//
//
//
//
//
//
module direct_interc_285 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_286__285 ( .A ( in[0] ) , 
    .X ( net_net_1939 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_1929 ( .A ( net_net_1930 ) , 
    .X ( out[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_1931 ( .A ( net_net_1933 ) , 
    .X ( net_net_1930 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_1934 ( .A ( net_net_1937 ) , 
    .X ( net_net_1933 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_1938 ( .A ( net_net_1939 ) , 
    .X ( net_net_1937 ) ) ;
endmodule


module direct_interc_284 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

wire aps_rename_14_ ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_285__284 ( .A ( in[0] ) , 
    .X ( aps_rename_14_ ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_1915 ( .A ( BUF_net_1917 ) , 
    .X ( out[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_1917 ( .A ( BUF_net_1920 ) , 
    .X ( BUF_net_1917 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_1920 ( .A ( BUF_net_1924 ) , 
    .X ( BUF_net_1920 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_1924 ( .A ( aps_rename_14_ ) , 
    .X ( BUF_net_1924 ) ) ;
endmodule


module direct_interc_283 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

wire aps_rename_13_ ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_284__283 ( .A ( in[0] ) , 
    .X ( aps_rename_13_ ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_1901 ( .A ( BUF_net_1903 ) , 
    .X ( out[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_1903 ( .A ( BUF_net_1906 ) , 
    .X ( BUF_net_1903 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_1906 ( .A ( BUF_net_1910 ) , 
    .X ( BUF_net_1906 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_1910 ( .A ( aps_rename_13_ ) , 
    .X ( BUF_net_1910 ) ) ;
endmodule


module direct_interc_282 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_283__282 ( .A ( in[0] ) , 
    .X ( net_net_1898 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_1889 ( .A ( net_net_1890 ) , 
    .X ( out[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_1891 ( .A ( net_net_1893 ) , 
    .X ( net_net_1890 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_1894 ( .A ( net_net_1897 ) , 
    .X ( net_net_1893 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_1898 ( .A ( net_net_1898 ) , 
    .X ( net_net_1897 ) ) ;
endmodule


module direct_interc_281 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_282__281 ( .A ( in[0] ) , 
    .X ( net_net_1886 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_1877 ( .A ( net_net_1881 ) , 
    .X ( out[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_1882 ( .A ( net_net_1885 ) , 
    .X ( net_net_1881 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_1886 ( .A ( net_net_1886 ) , 
    .X ( net_net_1885 ) ) ;
endmodule


module direct_interc_280 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_281__280 ( .A ( in[0] ) , 
    .X ( net_net_1874 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_1864 ( .A ( net_net_1865 ) , 
    .X ( out[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_1866 ( .A ( net_net_1868 ) , 
    .X ( net_net_1865 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_1869 ( .A ( net_net_1872 ) , 
    .X ( net_net_1868 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_1873 ( .A ( net_net_1874 ) , 
    .X ( net_net_1872 ) ) ;
endmodule


module direct_interc_279 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_280__279 ( .A ( in[0] ) , 
    .X ( net_net_1861 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_1852 ( .A ( net_net_1853 ) , 
    .X ( out[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_1854 ( .A ( net_net_1856 ) , 
    .X ( net_net_1853 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_1857 ( .A ( net_net_1857 ) , 
    .X ( net_net_1856 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_1858 ( .A ( net_net_1860 ) , 
    .X ( net_net_1857 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_1861 ( .A ( net_net_1861 ) , 
    .X ( net_net_1860 ) ) ;
endmodule


module direct_interc_278 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

wire aps_rename_12_ ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_279__278 ( .A ( in[0] ) , 
    .X ( aps_rename_12_ ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_1835 ( .A ( BUF_net_1837 ) , 
    .X ( out[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_1837 ( .A ( BUF_net_1840 ) , 
    .X ( BUF_net_1837 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_1840 ( .A ( BUF_net_1841 ) , 
    .X ( BUF_net_1840 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_1841 ( .A ( BUF_net_1844 ) , 
    .X ( BUF_net_1841 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_1844 ( .A ( BUF_net_1846 ) , 
    .X ( BUF_net_1844 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_1846 ( .A ( aps_rename_12_ ) , 
    .X ( BUF_net_1846 ) ) ;
endmodule


module direct_interc_277 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_278__277 ( .A ( in[0] ) , 
    .X ( net_net_1832 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_1822 ( .A ( net_net_1824 ) , 
    .X ( out[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_1825 ( .A ( net_net_1827 ) , 
    .X ( net_net_1824 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_1828 ( .A ( net_net_1831 ) , 
    .X ( net_net_1827 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_1832 ( .A ( net_net_1832 ) , 
    .X ( net_net_1831 ) ) ;
endmodule


module direct_interc_276 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_277__276 ( .A ( in[0] ) , 
    .X ( net_net_1820 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_1811 ( .A ( net_net_1812 ) , 
    .X ( out[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_1813 ( .A ( net_net_1815 ) , 
    .X ( net_net_1812 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_1816 ( .A ( net_net_1819 ) , 
    .X ( net_net_1815 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_1820 ( .A ( net_net_1820 ) , 
    .X ( net_net_1819 ) ) ;
endmodule


module direct_interc_275 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_276__275 ( .A ( in[0] ) , 
    .X ( net_net_1808 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_1799 ( .A ( net_net_1800 ) , 
    .X ( out[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_1801 ( .A ( net_net_1803 ) , 
    .X ( net_net_1800 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_1804 ( .A ( net_net_1807 ) , 
    .X ( net_net_1803 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_1808 ( .A ( net_net_1808 ) , 
    .X ( net_net_1807 ) ) ;
endmodule


module direct_interc_274 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_275__274 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_273 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_274__273 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_272 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_273__272 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_271 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_272__271 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_270 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_271__270 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_269 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_270__269 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_268 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_269__268 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_267 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_268__267 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_266 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_267__266 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_265 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_266__265 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_264 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_265__264 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_263 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_264__263 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_262 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_263__262 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_261 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_262__261 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_260 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_261__260 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_259 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_260__259 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_258 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_259__258 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_257 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_258__257 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_256 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_257__256 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_255 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_256__255 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_254 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_255__254 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_253 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_254__253 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_252 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_253__252 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_251 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_252__251 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_250 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_251__250 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_249 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_250__249 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_248 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_249__248 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_247 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_248__247 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_246 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_247__246 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_245 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_246__245 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_244 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_245__244 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_243 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_244__243 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_242 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_243__242 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_241 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_242__241 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_240 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_241__240 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_239 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_240__239 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_238 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_239__238 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_237 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_238__237 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_236 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_237__236 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_235 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_236__235 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_234 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_235__234 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_233 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_234__233 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_232 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_233__232 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_231 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_232__231 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_230 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_231__230 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_229 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_230__229 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_228 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_229__228 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_227 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_228__227 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_226 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_227__226 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_225 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_226__225 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_224 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_225__224 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_223 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_224__223 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_222 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_223__222 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_221 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_222__221 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_220 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_221__220 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_219 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_220__219 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_218 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_219__218 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_217 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_218__217 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_216 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_217__216 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_215 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_216__215 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_214 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_215__214 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_213 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_214__213 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_212 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_213__212 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_211 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_212__211 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_210 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_211__210 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_209 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_210__209 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_208 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_209__208 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_207 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_208__207 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_206 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_207__206 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_205 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_206__205 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_204 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_205__204 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_203 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_204__203 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_202 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_203__202 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_201 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_202__201 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_200 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_201__200 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_199 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_200__199 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_198 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_199__198 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_197 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_198__197 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_196 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_197__196 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_195 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_196__195 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_194 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_195__194 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_193 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_194__193 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_192 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_193__192 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_191 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_192__191 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_190 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_191__190 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_189 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_190__189 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_188 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_189__188 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_187 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_188__187 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_186 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_187__186 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_185 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_186__185 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_184 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_185__184 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_183 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_184__183 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_182 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_183__182 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_181 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_182__181 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_180 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_181__180 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_179 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_180__179 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_178 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_179__178 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_177 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_178__177 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_176 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_177__176 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_175 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_176__175 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_174 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_175__174 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_173 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_174__173 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_172 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_173__172 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_171 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_172__171 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_170 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_171__170 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_169 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_170__169 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_168 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_169__168 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_167 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_168__167 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_166 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_167__166 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_165 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_166__165 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_164 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_165__164 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_163 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_164__163 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_162 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_163__162 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_161 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_162__161 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_160 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_161__160 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_159 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_160__159 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_158 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_159__158 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_157 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_158__157 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_156 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_157__156 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_155 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_156__155 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_154 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_155__154 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_153 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_154__153 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_152 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_153__152 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_151 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_152__151 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_150 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_151__150 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_149 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_150__149 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_148 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_149__148 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_147 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_148__147 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_146 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_147__146 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_145 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_146__145 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_144 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_145__144 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_143 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_144__143 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_142 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

wire aps_rename_11_ ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_143__142 ( .A ( in[0] ) , 
    .X ( aps_rename_11_ ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_428 ( .A ( BUF_net_430 ) , 
    .X ( out[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_430 ( .A ( BUF_net_433 ) , 
    .X ( BUF_net_430 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_433 ( .A ( BUF_net_437 ) , 
    .X ( BUF_net_433 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_437 ( .A ( aps_rename_11_ ) , 
    .X ( BUF_net_437 ) ) ;
endmodule


module direct_interc_141 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

wire aps_rename_10_ ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_142__141 ( .A ( in[0] ) , 
    .X ( aps_rename_10_ ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_414 ( .A ( BUF_net_416 ) , 
    .X ( out[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_416 ( .A ( BUF_net_419 ) , 
    .X ( BUF_net_416 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_419 ( .A ( BUF_net_423 ) , 
    .X ( BUF_net_419 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_423 ( .A ( aps_rename_10_ ) , 
    .X ( BUF_net_423 ) ) ;
endmodule


module direct_interc_140 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

wire aps_rename_9_ ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_141__140 ( .A ( in[0] ) , 
    .X ( aps_rename_9_ ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_399 ( .A ( BUF_net_401 ) , 
    .X ( out[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_401 ( .A ( BUF_net_404 ) , 
    .X ( BUF_net_401 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_404 ( .A ( BUF_net_408 ) , 
    .X ( BUF_net_404 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_408 ( .A ( aps_rename_9_ ) , 
    .X ( BUF_net_408 ) ) ;
endmodule


module direct_interc_139 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

wire aps_rename_8_ ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_140__139 ( .A ( in[0] ) , 
    .X ( aps_rename_8_ ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_385 ( .A ( BUF_net_387 ) , 
    .X ( out[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_387 ( .A ( BUF_net_390 ) , 
    .X ( BUF_net_387 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_390 ( .A ( BUF_net_394 ) , 
    .X ( BUF_net_390 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_394 ( .A ( aps_rename_8_ ) , 
    .X ( BUF_net_394 ) ) ;
endmodule


module direct_interc_138 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

wire aps_rename_7_ ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_139__138 ( .A ( in[0] ) , 
    .X ( aps_rename_7_ ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_372 ( .A ( BUF_net_374 ) , 
    .X ( out[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_374 ( .A ( BUF_net_377 ) , 
    .X ( BUF_net_374 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_377 ( .A ( BUF_net_381 ) , 
    .X ( BUF_net_377 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_381 ( .A ( aps_rename_7_ ) , 
    .X ( BUF_net_381 ) ) ;
endmodule


module direct_interc_137 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

wire aps_rename_6_ ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_138__137 ( .A ( in[0] ) , 
    .X ( aps_rename_6_ ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_358 ( .A ( BUF_net_360 ) , 
    .X ( out[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_360 ( .A ( BUF_net_363 ) , 
    .X ( BUF_net_360 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_363 ( .A ( BUF_net_367 ) , 
    .X ( BUF_net_363 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_367 ( .A ( aps_rename_6_ ) , 
    .X ( BUF_net_367 ) ) ;
endmodule


module direct_interc_136 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

wire aps_rename_5_ ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_137__136 ( .A ( in[0] ) , 
    .X ( aps_rename_5_ ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_345 ( .A ( BUF_net_347 ) , 
    .X ( out[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_347 ( .A ( BUF_net_350 ) , 
    .X ( BUF_net_347 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_350 ( .A ( BUF_net_351 ) , 
    .X ( BUF_net_350 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_351 ( .A ( BUF_net_354 ) , 
    .X ( BUF_net_351 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_354 ( .A ( aps_rename_5_ ) , 
    .X ( BUF_net_354 ) ) ;
endmodule


module direct_interc_135 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

wire aps_rename_4_ ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_136__135 ( .A ( in[0] ) , 
    .X ( aps_rename_4_ ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_328 ( .A ( BUF_net_330 ) , 
    .X ( out[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_330 ( .A ( BUF_net_333 ) , 
    .X ( BUF_net_330 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_333 ( .A ( BUF_net_337 ) , 
    .X ( BUF_net_333 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_337 ( .A ( BUF_net_339 ) , 
    .X ( BUF_net_337 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_339 ( .A ( aps_rename_4_ ) , 
    .X ( BUF_net_339 ) ) ;
endmodule


module direct_interc_134 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

wire aps_rename_3_ ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_135__134 ( .A ( in[0] ) , 
    .X ( aps_rename_3_ ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_314 ( .A ( BUF_net_316 ) , 
    .X ( out[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_316 ( .A ( BUF_net_319 ) , 
    .X ( BUF_net_316 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_319 ( .A ( BUF_net_323 ) , 
    .X ( BUF_net_319 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_323 ( .A ( aps_rename_3_ ) , 
    .X ( BUF_net_323 ) ) ;
endmodule


module direct_interc_133 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

wire aps_rename_2_ ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_134__133 ( .A ( in[0] ) , 
    .X ( aps_rename_2_ ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_301 ( .A ( BUF_net_303 ) , 
    .X ( out[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_303 ( .A ( BUF_net_306 ) , 
    .X ( BUF_net_303 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_306 ( .A ( BUF_net_310 ) , 
    .X ( BUF_net_306 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_310 ( .A ( aps_rename_2_ ) , 
    .X ( BUF_net_310 ) ) ;
endmodule


module direct_interc_132 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

wire aps_rename_1_ ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_133__132 ( .A ( in[0] ) , 
    .X ( aps_rename_1_ ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_288 ( .A ( BUF_net_290 ) , 
    .X ( out[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_290 ( .A ( BUF_net_293 ) , 
    .X ( BUF_net_290 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_293 ( .A ( BUF_net_297 ) , 
    .X ( BUF_net_293 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_297 ( .A ( aps_rename_1_ ) , 
    .X ( BUF_net_297 ) ) ;
endmodule


module direct_interc_131 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_132__131 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_130 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_131__130 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_129 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_130__129 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_128 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_129__128 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_127 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_128__127 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_126 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_127__126 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_125 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_126__125 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_124 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_125__124 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_123 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_124__123 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_122 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_123__122 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_121 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_122__121 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_120 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_121__120 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_119 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_120__119 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_118 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_119__118 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_117 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_118__117 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_116 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_117__116 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_115 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_116__115 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_114 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_115__114 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_113 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_114__113 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_112 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_113__112 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_111 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_112__111 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_110 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_111__110 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_109 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_110__109 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_108 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_109__108 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_107 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_108__107 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_106 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_107__106 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_105 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_106__105 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_104 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_105__104 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_103 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_104__103 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_102 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_103__102 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_101 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_102__101 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_100 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_101__100 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_99 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_100__99 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_98 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_99__98 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_97 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_98__97 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_96 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_97__96 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_95 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_96__95 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_94 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_95__94 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_93 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_94__93 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_92 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_93__92 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_91 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_92__91 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_90 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_91__90 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_89 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_90__89 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_88 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_89__88 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_87 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_88__87 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_86 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_87__86 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_85 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_86__85 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_84 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_85__84 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_83 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_84__83 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_82 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_83__82 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_81 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_82__81 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_80 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_81__80 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_79 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_80__79 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_78 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_79__78 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_77 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_78__77 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_76 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_77__76 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_75 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_76__75 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_74 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_75__74 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_73 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_74__73 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_72 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_73__72 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_71 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_72__71 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_70 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_71__70 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_69 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_70__69 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_68 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_69__68 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_67 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_68__67 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_66 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_67__66 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_65 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_66__65 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_64 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_65__64 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_63 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_64__63 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_62 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_63__62 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_61 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_62__61 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_60 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_61__60 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_59 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_60__59 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_58 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_59__58 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_57 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_58__57 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_56 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_57__56 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_55 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_56__55 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_54 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_55__54 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_53 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_54__53 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_52 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_53__52 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_51 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_52__51 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_50 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_51__50 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_49 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_50__49 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_48 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_49__48 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_47 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_48__47 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_46 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_47__46 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_45 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_46__45 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_44 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_45__44 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_43 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_44__43 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_42 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_43__42 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_41 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_42__41 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_40 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_41__40 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_39 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_40__39 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_38 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_39__38 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_37 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_38__37 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_36 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_37__36 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_35 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_36__35 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_34 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_35__34 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_33 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_34__33 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_32 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_33__32 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_31 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_32__31 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_30 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_31__30 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_29 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_30__29 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_28 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_29__28 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_27 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_28__27 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_26 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_27__26 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_25 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_26__25 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_24 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_25__24 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_23 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_24__23 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_22 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_23__22 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_21 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_22__21 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_20 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_21__20 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_19 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_20__19 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_18 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_19__18 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_17 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_18__17 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_16 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_17__16 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_15 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_16__15 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_14 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_15__14 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_13 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_14__13 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_12 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_13__12 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_11 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_12__11 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_10 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_11__10 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_9 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_10__9 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_8 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_9__8 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_7 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_8__7 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_6 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_7__6 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_5 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_6__5 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_4 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_5__4 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_3 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_4__3 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_2 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_3__2 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_1 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_2__1 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_0 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_1__0 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module mux_tree_tapbuf_size8_mem_3_2 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd1_1 FTB_17__56 ( .A ( mem_out[3] ) , 
    .X ( net_net_85 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_RR_85 ( .A ( net_net_85 ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size8_mem_2_3 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_16__55 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size8_mem_1_4 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_15__54 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size8_mem_0_4 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_14__53 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size8_mem_9 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_13__52 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size8_mem_6_2 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_12__51 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size8_mem_5_2 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_11__50 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size8_mem_4_2 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_10__49 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_44 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size8_3_2 ( in , sram , sram_inv , out , p0 ) ;
input  [0:7] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;

const1_44 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( in[2] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[4] ) , .A1 ( in[3] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[6] ) , .A1 ( in[5] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
endmodule


module const1_15_10 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size8_2_3 ( in , sram , sram_inv , out , p0 ) ;
input  [0:7] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;

const1_15_10 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( in[2] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[4] ) , .A1 ( in[3] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[6] ) , .A1 ( in[5] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
endmodule


module const1_14_11 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size8_1_4 ( in , sram , sram_inv , out , p0 ) ;
input  [0:7] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;

const1_14_11 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( in[2] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[4] ) , .A1 ( in[3] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[6] ) , .A1 ( in[5] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
endmodule


module const1_13_11 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size8_0_4 ( in , sram , sram_inv , out , p0 ) ;
input  [0:7] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;

const1_13_11 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( in[2] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[4] ) , .A1 ( in[3] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[6] ) , .A1 ( in[5] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
endmodule


module const1_12_11 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size8_9 ( in , sram , sram_inv , out , p0 ) ;
input  [0:7] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;

const1_12_11 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( in[2] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[4] ) , .A1 ( in[3] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[6] ) , .A1 ( in[5] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
endmodule


module const1_11_11 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size8_6_2 ( in , sram , sram_inv , out , p0 ) ;
input  [0:7] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;

const1_11_11 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( in[2] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[4] ) , .A1 ( in[3] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[6] ) , .A1 ( in[5] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
endmodule


module const1_10_11 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size8_5_2 ( in , sram , sram_inv , out , p0 ) ;
input  [0:7] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;

const1_10_11 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( in[2] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[4] ) , .A1 ( in[3] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[6] ) , .A1 ( in[5] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
endmodule


module const1_9_11 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size8_4_2 ( in , sram , sram_inv , out , p0 ) ;
input  [0:7] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;

const1_9_11 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( in[2] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[4] ) , .A1 ( in[3] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[6] ) , .A1 ( in[5] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
endmodule


module mux_tree_tapbuf_size10_mem_4_3 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_9__48 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size10_mem_3_3 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_8__47 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size10_mem_16 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_7__46 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size10_mem_7_2 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_6__45 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size10_mem_6_3 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_5__44 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size10_mem_5_3 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_4__43 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size10_mem_2_3 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_3__42 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size10_mem_1_3 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_2__41 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size10_mem_0_5 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_1__40 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_8_11 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size10_4_3 ( in , sram , sram_inv , out , p0 ) ;
input  [0:9] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

const1_8_11 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[6] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[8] ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[9] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
endmodule


module const1_7_11 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size10_3_3 ( in , sram , sram_inv , out , p0 ) ;
input  [0:9] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

const1_7_11 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[6] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[8] ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[9] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
endmodule


module const1_6_12 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size10_16 ( in , sram , sram_inv , out , p0 ) ;
input  [0:9] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

const1_6_12 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[6] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[8] ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[9] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
endmodule


module const1_5_12 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size10_7_2 ( in , sram , sram_inv , out , p0 ) ;
input  [0:9] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

const1_5_12 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[6] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[8] ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[9] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
endmodule


module const1_4_12 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size10_6_3 ( in , sram , sram_inv , out , p0 ) ;
input  [0:9] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

const1_4_12 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[6] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[8] ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[9] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
endmodule


module const1_3_12 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size10_5_3 ( in , sram , sram_inv , out , p0 ) ;
input  [0:9] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

const1_3_12 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[6] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[8] ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[9] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
endmodule


module const1_2_12 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size10_2_3 ( in , sram , sram_inv , out , p0 ) ;
input  [0:9] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

const1_2_12 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[6] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[8] ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[9] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
endmodule


module const1_1_12 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size10_1_3 ( in , sram , sram_inv , out , p0 ) ;
input  [0:9] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

const1_1_12 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[6] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[8] ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[9] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
endmodule


module const1_0_13 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size10_0_5 ( in , sram , sram_inv , out , p0 ) ;
input  [0:9] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

const1_0_13 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[6] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[8] ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[9] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
endmodule


module cby_1__1_ ( prog_clk , chany_bottom_in , chany_top_in , ccff_head , 
    chany_bottom_out , chany_top_out , right_grid_pin_52_ , left_grid_pin_0_ , 
    left_grid_pin_1_ , left_grid_pin_2_ , left_grid_pin_3_ , 
    left_grid_pin_4_ , left_grid_pin_5_ , left_grid_pin_6_ , 
    left_grid_pin_7_ , left_grid_pin_8_ , left_grid_pin_9_ , 
    left_grid_pin_10_ , left_grid_pin_11_ , left_grid_pin_12_ , 
    left_grid_pin_13_ , left_grid_pin_14_ , left_grid_pin_15_ , ccff_tail ) ;
input  [0:0] prog_clk ;
input  [0:19] chany_bottom_in ;
input  [0:19] chany_top_in ;
input  [0:0] ccff_head ;
output [0:19] chany_bottom_out ;
output [0:19] chany_top_out ;
output [0:0] right_grid_pin_52_ ;
output [0:0] left_grid_pin_0_ ;
output [0:0] left_grid_pin_1_ ;
output [0:0] left_grid_pin_2_ ;
output [0:0] left_grid_pin_3_ ;
output [0:0] left_grid_pin_4_ ;
output [0:0] left_grid_pin_5_ ;
output [0:0] left_grid_pin_6_ ;
output [0:0] left_grid_pin_7_ ;
output [0:0] left_grid_pin_8_ ;
output [0:0] left_grid_pin_9_ ;
output [0:0] left_grid_pin_10_ ;
output [0:0] left_grid_pin_11_ ;
output [0:0] left_grid_pin_12_ ;
output [0:0] left_grid_pin_13_ ;
output [0:0] left_grid_pin_14_ ;
output [0:0] left_grid_pin_15_ ;
output [0:0] ccff_tail ;

wire [0:3] mux_tree_tapbuf_size10_0_sram ;
wire [0:3] mux_tree_tapbuf_size10_0_sram_inv ;
wire [0:3] mux_tree_tapbuf_size10_1_sram ;
wire [0:3] mux_tree_tapbuf_size10_1_sram_inv ;
wire [0:3] mux_tree_tapbuf_size10_2_sram ;
wire [0:3] mux_tree_tapbuf_size10_2_sram_inv ;
wire [0:3] mux_tree_tapbuf_size10_3_sram ;
wire [0:3] mux_tree_tapbuf_size10_3_sram_inv ;
wire [0:3] mux_tree_tapbuf_size10_4_sram ;
wire [0:3] mux_tree_tapbuf_size10_4_sram_inv ;
wire [0:3] mux_tree_tapbuf_size10_5_sram ;
wire [0:3] mux_tree_tapbuf_size10_5_sram_inv ;
wire [0:3] mux_tree_tapbuf_size10_6_sram ;
wire [0:3] mux_tree_tapbuf_size10_6_sram_inv ;
wire [0:3] mux_tree_tapbuf_size10_7_sram ;
wire [0:3] mux_tree_tapbuf_size10_7_sram_inv ;
wire [0:3] mux_tree_tapbuf_size10_8_sram ;
wire [0:3] mux_tree_tapbuf_size10_8_sram_inv ;
wire [0:0] mux_tree_tapbuf_size10_mem_0_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size10_mem_1_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size10_mem_2_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size10_mem_3_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size10_mem_4_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size10_mem_5_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size10_mem_6_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size10_mem_7_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size10_mem_8_ccff_tail ;
wire [0:3] mux_tree_tapbuf_size8_0_sram ;
wire [0:3] mux_tree_tapbuf_size8_0_sram_inv ;
wire [0:3] mux_tree_tapbuf_size8_1_sram ;
wire [0:3] mux_tree_tapbuf_size8_1_sram_inv ;
wire [0:3] mux_tree_tapbuf_size8_2_sram ;
wire [0:3] mux_tree_tapbuf_size8_2_sram_inv ;
wire [0:3] mux_tree_tapbuf_size8_3_sram ;
wire [0:3] mux_tree_tapbuf_size8_3_sram_inv ;
wire [0:3] mux_tree_tapbuf_size8_4_sram ;
wire [0:3] mux_tree_tapbuf_size8_4_sram_inv ;
wire [0:3] mux_tree_tapbuf_size8_5_sram ;
wire [0:3] mux_tree_tapbuf_size8_5_sram_inv ;
wire [0:3] mux_tree_tapbuf_size8_6_sram ;
wire [0:3] mux_tree_tapbuf_size8_6_sram_inv ;
wire [0:3] mux_tree_tapbuf_size8_7_sram ;
wire [0:3] mux_tree_tapbuf_size8_7_sram_inv ;
wire [0:0] mux_tree_tapbuf_size8_mem_0_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size8_mem_1_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size8_mem_2_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size8_mem_3_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size8_mem_4_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size8_mem_5_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size8_mem_6_ccff_tail ;

mux_tree_tapbuf_size10_0_5 mux_left_ipin_0 (
    .in ( { chany_bottom_in[0] , chany_top_in[0] , chany_bottom_in[2] , 
        chany_top_in[2] , chany_bottom_in[4] , chany_top_in[4] , 
        chany_bottom_in[10] , chany_top_in[10] , chany_bottom_in[16] , 
        chany_top_in[16] } ) ,
    .sram ( mux_tree_tapbuf_size10_0_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size10_0_sram_inv ) , 
    .out ( right_grid_pin_52_ ) , .p0 ( optlc_net_96 ) ) ;
mux_tree_tapbuf_size10_1_3 mux_right_ipin_0 (
    .in ( { chany_bottom_in[1] , chany_top_in[1] , chany_bottom_in[3] , 
        chany_top_in[3] , chany_bottom_in[5] , chany_top_in[5] , 
        chany_bottom_in[11] , chany_top_in[11] , chany_bottom_in[17] , 
        chany_top_in[17] } ) ,
    .sram ( mux_tree_tapbuf_size10_1_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size10_1_sram_inv ) , 
    .out ( left_grid_pin_0_ ) , .p0 ( optlc_net_96 ) ) ;
mux_tree_tapbuf_size10_2_3 mux_right_ipin_1 (
    .in ( { chany_bottom_in[0] , chany_top_in[0] , chany_bottom_in[2] , 
        chany_top_in[2] , chany_bottom_in[6] , chany_top_in[6] , 
        chany_bottom_in[12] , chany_top_in[12] , chany_bottom_in[18] , 
        chany_top_in[18] } ) ,
    .sram ( mux_tree_tapbuf_size10_2_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size10_2_sram_inv ) , 
    .out ( left_grid_pin_1_ ) , .p0 ( optlc_net_97 ) ) ;
mux_tree_tapbuf_size10_5_3 mux_right_ipin_4 (
    .in ( { chany_bottom_in[1] , chany_top_in[1] , chany_bottom_in[3] , 
        chany_top_in[3] , chany_bottom_in[5] , chany_top_in[5] , 
        chany_bottom_in[9] , chany_top_in[9] , chany_bottom_in[15] , 
        chany_top_in[15] } ) ,
    .sram ( mux_tree_tapbuf_size10_3_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size10_3_sram_inv ) , 
    .out ( left_grid_pin_4_ ) , .p0 ( optlc_net_97 ) ) ;
mux_tree_tapbuf_size10_6_3 mux_right_ipin_5 (
    .in ( { chany_bottom_in[0] , chany_top_in[0] , chany_bottom_in[2] , 
        chany_top_in[2] , chany_bottom_in[6] , chany_top_in[6] , 
        chany_bottom_in[10] , chany_top_in[10] , chany_bottom_in[16] , 
        chany_top_in[16] } ) ,
    .sram ( mux_tree_tapbuf_size10_4_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size10_4_sram_inv ) , 
    .out ( left_grid_pin_5_ ) , .p0 ( optlc_net_96 ) ) ;
mux_tree_tapbuf_size10_7_2 mux_right_ipin_8 (
    .in ( { chany_bottom_in[1] , chany_top_in[1] , chany_bottom_in[3] , 
        chany_top_in[3] , chany_bottom_in[9] , chany_top_in[9] , 
        chany_bottom_in[13] , chany_top_in[13] , chany_bottom_in[19] , 
        chany_top_in[19] } ) ,
    .sram ( mux_tree_tapbuf_size10_5_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size10_5_sram_inv ) , 
    .out ( left_grid_pin_8_ ) , .p0 ( optlc_net_95 ) ) ;
mux_tree_tapbuf_size10_16 mux_right_ipin_9 (
    .in ( { chany_bottom_in[0] , chany_top_in[0] , chany_bottom_in[2] , 
        chany_top_in[2] , chany_bottom_in[4] , chany_top_in[4] , 
        chany_bottom_in[10] , chany_top_in[10] , chany_bottom_in[14] , 
        chany_top_in[14] } ) ,
    .sram ( mux_tree_tapbuf_size10_6_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size10_6_sram_inv ) , 
    .out ( left_grid_pin_9_ ) , .p0 ( optlc_net_95 ) ) ;
mux_tree_tapbuf_size10_3_3 mux_right_ipin_12 (
    .in ( { chany_bottom_in[1] , chany_top_in[1] , chany_bottom_in[3] , 
        chany_top_in[3] , chany_bottom_in[7] , chany_top_in[7] , 
        chany_bottom_in[13] , chany_top_in[13] , chany_bottom_in[17] , 
        chany_top_in[17] } ) ,
    .sram ( mux_tree_tapbuf_size10_7_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size10_7_sram_inv ) , 
    .out ( left_grid_pin_12_ ) , .p0 ( optlc_net_96 ) ) ;
mux_tree_tapbuf_size10_4_3 mux_right_ipin_13 (
    .in ( { chany_bottom_in[0] , chany_top_in[0] , chany_bottom_in[2] , 
        chany_top_in[2] , chany_bottom_in[8] , chany_top_in[8] , 
        chany_bottom_in[14] , chany_top_in[14] , chany_bottom_in[18] , 
        chany_top_in[18] } ) ,
    .sram ( mux_tree_tapbuf_size10_8_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size10_8_sram_inv ) , 
    .out ( left_grid_pin_13_ ) , .p0 ( optlc_net_96 ) ) ;
mux_tree_tapbuf_size10_mem_0_5 mem_left_ipin_0 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( ccff_head ) , 
    .ccff_tail ( mux_tree_tapbuf_size10_mem_0_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size10_0_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size10_0_sram_inv ) ) ;
mux_tree_tapbuf_size10_mem_1_3 mem_right_ipin_0 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size10_mem_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size10_mem_1_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size10_1_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size10_1_sram_inv ) ) ;
mux_tree_tapbuf_size10_mem_2_3 mem_right_ipin_1 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size10_mem_1_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size10_mem_2_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size10_2_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size10_2_sram_inv ) ) ;
mux_tree_tapbuf_size10_mem_5_3 mem_right_ipin_4 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size8_mem_1_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size10_mem_3_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size10_3_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size10_3_sram_inv ) ) ;
mux_tree_tapbuf_size10_mem_6_3 mem_right_ipin_5 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size10_mem_3_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size10_mem_4_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size10_4_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size10_4_sram_inv ) ) ;
mux_tree_tapbuf_size10_mem_7_2 mem_right_ipin_8 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size8_mem_3_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size10_mem_5_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size10_5_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size10_5_sram_inv ) ) ;
mux_tree_tapbuf_size10_mem_16 mem_right_ipin_9 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size10_mem_5_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size10_mem_6_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size10_6_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size10_6_sram_inv ) ) ;
mux_tree_tapbuf_size10_mem_3_3 mem_right_ipin_12 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size8_mem_5_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size10_mem_7_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size10_7_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size10_7_sram_inv ) ) ;
mux_tree_tapbuf_size10_mem_4_3 mem_right_ipin_13 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size10_mem_7_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size10_mem_8_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size10_8_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size10_8_sram_inv ) ) ;
mux_tree_tapbuf_size8_4_2 mux_right_ipin_2 (
    .in ( { chany_bottom_in[1] , chany_top_in[1] , chany_bottom_in[3] , 
        chany_top_in[3] , chany_bottom_in[7] , chany_top_in[7] , 
        chany_bottom_in[15] , chany_top_in[15] } ) ,
    .sram ( mux_tree_tapbuf_size8_0_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size8_0_sram_inv ) , 
    .out ( left_grid_pin_2_ ) , .p0 ( optlc_net_97 ) ) ;
mux_tree_tapbuf_size8_5_2 mux_right_ipin_3 (
    .in ( { chany_bottom_in[0] , chany_top_in[0] , chany_bottom_in[2] , 
        chany_top_in[2] , chany_bottom_in[8] , chany_top_in[8] , 
        chany_bottom_in[16] , chany_top_in[16] } ) ,
    .sram ( mux_tree_tapbuf_size8_1_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size8_1_sram_inv ) , 
    .out ( left_grid_pin_3_ ) , .p0 ( optlc_net_96 ) ) ;
mux_tree_tapbuf_size8_6_2 mux_right_ipin_6 (
    .in ( { chany_bottom_in[1] , chany_top_in[1] , chany_bottom_in[3] , 
        chany_top_in[3] , chany_bottom_in[11] , chany_top_in[11] , 
        chany_bottom_in[19] , chany_top_in[19] } ) ,
    .sram ( mux_tree_tapbuf_size8_2_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size8_2_sram_inv ) , 
    .out ( left_grid_pin_6_ ) , .p0 ( optlc_net_97 ) ) ;
mux_tree_tapbuf_size8_9 mux_right_ipin_7 (
    .in ( { chany_bottom_in[0] , chany_top_in[0] , chany_bottom_in[2] , 
        chany_top_in[2] , chany_bottom_in[4] , chany_top_in[4] , 
        chany_bottom_in[12] , chany_top_in[12] } ) ,
    .sram ( mux_tree_tapbuf_size8_3_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size8_3_sram_inv ) , 
    .out ( left_grid_pin_7_ ) , .p0 ( optlc_net_96 ) ) ;
mux_tree_tapbuf_size8_0_4 mux_right_ipin_10 (
    .in ( { chany_bottom_in[1] , chany_top_in[1] , chany_bottom_in[3] , 
        chany_top_in[3] , chany_bottom_in[7] , chany_top_in[7] , 
        chany_bottom_in[15] , chany_top_in[15] } ) ,
    .sram ( mux_tree_tapbuf_size8_4_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size8_4_sram_inv ) , 
    .out ( left_grid_pin_10_ ) , .p0 ( optlc_net_95 ) ) ;
mux_tree_tapbuf_size8_1_4 mux_right_ipin_11 (
    .in ( { chany_bottom_in[0] , chany_top_in[0] , chany_bottom_in[2] , 
        chany_top_in[2] , chany_bottom_in[8] , chany_top_in[8] , 
        chany_bottom_in[16] , chany_top_in[16] } ) ,
    .sram ( mux_tree_tapbuf_size8_5_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size8_5_sram_inv ) , 
    .out ( left_grid_pin_11_ ) , .p0 ( optlc_net_96 ) ) ;
mux_tree_tapbuf_size8_2_3 mux_right_ipin_14 (
    .in ( { chany_bottom_in[1] , chany_top_in[1] , chany_bottom_in[3] , 
        chany_top_in[3] , chany_bottom_in[11] , chany_top_in[11] , 
        chany_bottom_in[19] , chany_top_in[19] } ) ,
    .sram ( mux_tree_tapbuf_size8_6_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size8_6_sram_inv ) , 
    .out ( left_grid_pin_14_ ) , .p0 ( optlc_net_97 ) ) ;
mux_tree_tapbuf_size8_3_2 mux_right_ipin_15 (
    .in ( { chany_bottom_in[0] , chany_top_in[0] , chany_bottom_in[2] , 
        chany_top_in[2] , chany_bottom_in[4] , chany_top_in[4] , 
        chany_bottom_in[12] , chany_top_in[12] } ) ,
    .sram ( mux_tree_tapbuf_size8_7_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size8_7_sram_inv ) , 
    .out ( left_grid_pin_15_ ) , .p0 ( optlc_net_96 ) ) ;
mux_tree_tapbuf_size8_mem_4_2 mem_right_ipin_2 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size10_mem_2_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size8_mem_0_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size8_0_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size8_0_sram_inv ) ) ;
mux_tree_tapbuf_size8_mem_5_2 mem_right_ipin_3 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size8_mem_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size8_mem_1_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size8_1_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size8_1_sram_inv ) ) ;
mux_tree_tapbuf_size8_mem_6_2 mem_right_ipin_6 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size10_mem_4_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size8_mem_2_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size8_2_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size8_2_sram_inv ) ) ;
mux_tree_tapbuf_size8_mem_9 mem_right_ipin_7 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size8_mem_2_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size8_mem_3_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size8_3_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size8_3_sram_inv ) ) ;
mux_tree_tapbuf_size8_mem_0_4 mem_right_ipin_10 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size10_mem_6_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size8_mem_4_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size8_4_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size8_4_sram_inv ) ) ;
mux_tree_tapbuf_size8_mem_1_4 mem_right_ipin_11 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size8_mem_4_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size8_mem_5_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size8_5_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size8_5_sram_inv ) ) ;
mux_tree_tapbuf_size8_mem_2_3 mem_right_ipin_14 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size10_mem_8_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size8_mem_6_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size8_6_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size8_6_sram_inv ) ) ;
mux_tree_tapbuf_size8_mem_3_2 mem_right_ipin_15 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size8_mem_6_ccff_tail ) , 
    .ccff_tail ( ccff_tail ) , .mem_out ( mux_tree_tapbuf_size8_7_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size8_7_sram_inv ) ) ;
sky130_fd_sc_hd__dlygate4sd1_1 FTB_1__0 ( .A ( chany_bottom_in[0] ) , 
    .X ( chany_top_out[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd1_1 FTB_2__1 ( .A ( chany_bottom_in[1] ) , 
    .X ( chany_top_out[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd1_1 FTB_3__2 ( .A ( chany_bottom_in[2] ) , 
    .X ( chany_top_out[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd1_1 FTB_4__3 ( .A ( chany_bottom_in[3] ) , 
    .X ( chany_top_out[3] ) ) ;
sky130_fd_sc_hd__conb_1 optlc_94 ( .LO ( SYNOPSYS_UNCONNECTED_1 ) , 
    .HI ( optlc_net_95 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_96 ( .LO ( SYNOPSYS_UNCONNECTED_2 ) , 
    .HI ( optlc_net_96 ) ) ;
sky130_fd_sc_hd__dlygate4sd1_1 FTB_7__6 ( .A ( chany_bottom_in[6] ) , 
    .X ( chany_top_out[6] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_9__8 ( .A ( chany_bottom_in[8] ) , 
    .X ( aps_rename_3_ ) ) ;
sky130_fd_sc_hd__dlygate4sd1_1 FTB_10__9 ( .A ( chany_bottom_in[9] ) , 
    .X ( chany_top_out[9] ) ) ;
sky130_fd_sc_hd__conb_1 optlc_98 ( .LO ( SYNOPSYS_UNCONNECTED_3 ) , 
    .HI ( optlc_net_97 ) ) ;
sky130_fd_sc_hd__dlygate4sd1_1 FTB_12__11 ( .A ( chany_bottom_in[11] ) , 
    .X ( chany_top_out[11] ) ) ;
sky130_fd_sc_hd__dlygate4sd1_1 FTB_13__12 ( .A ( chany_bottom_in[12] ) , 
    .X ( chany_top_out[12] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_15__14 ( .A ( chany_bottom_in[14] ) , 
    .X ( aps_rename_4_ ) ) ;
sky130_fd_sc_hd__dlygate4sd1_1 FTB_16__15 ( .A ( chany_bottom_in[15] ) , 
    .X ( chany_top_out[15] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_17__16 ( .A ( chany_bottom_in[16] ) , 
    .X ( aps_rename_5_ ) ) ;
sky130_fd_sc_hd__dlygate4sd1_1 FTB_19__18 ( .A ( chany_bottom_in[18] ) , 
    .X ( chany_top_out[18] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_20__19 ( .A ( chany_bottom_in[19] ) , 
    .X ( aps_rename_6_ ) ) ;
sky130_fd_sc_hd__dlygate4sd1_1 FTB_21__20 ( .A ( chany_top_in[0] ) , 
    .X ( chany_bottom_out[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd1_1 FTB_22__21 ( .A ( chany_top_in[1] ) , 
    .X ( chany_bottom_out[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd1_1 FTB_23__22 ( .A ( chany_top_in[2] ) , 
    .X ( chany_bottom_out[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd1_1 FTB_24__23 ( .A ( chany_top_in[3] ) , 
    .X ( chany_bottom_out[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd1_1 FTB_25__24 ( .A ( chany_top_in[4] ) , 
    .X ( chany_bottom_out[4] ) ) ;
sky130_fd_sc_hd__dlygate4sd1_1 FTB_27__26 ( .A ( chany_top_in[6] ) , 
    .X ( chany_bottom_out[6] ) ) ;
sky130_fd_sc_hd__dlygate4sd1_1 FTB_28__27 ( .A ( chany_top_in[7] ) , 
    .X ( chany_bottom_out[7] ) ) ;
sky130_fd_sc_hd__dlygate4sd1_1 FTB_29__28 ( .A ( chany_top_in[8] ) , 
    .X ( chany_bottom_out[8] ) ) ;
sky130_fd_sc_hd__dlygate4sd1_1 FTB_30__29 ( .A ( chany_top_in[9] ) , 
    .X ( chany_bottom_out[9] ) ) ;
sky130_fd_sc_hd__dlygate4sd1_1 FTB_31__30 ( .A ( chany_top_in[10] ) , 
    .X ( chany_bottom_out[10] ) ) ;
sky130_fd_sc_hd__dlygate4sd1_1 FTB_32__31 ( .A ( chany_top_in[11] ) , 
    .X ( chany_bottom_out[11] ) ) ;
sky130_fd_sc_hd__dlygate4sd1_1 FTB_33__32 ( .A ( chany_top_in[12] ) , 
    .X ( chany_bottom_out[12] ) ) ;
sky130_fd_sc_hd__dlygate4sd1_1 FTB_34__33 ( .A ( chany_top_in[13] ) , 
    .X ( chany_bottom_out[13] ) ) ;
sky130_fd_sc_hd__dlygate4sd1_1 FTB_35__34 ( .A ( chany_top_in[14] ) , 
    .X ( chany_bottom_out[14] ) ) ;
sky130_fd_sc_hd__dlygate4sd1_1 FTB_36__35 ( .A ( chany_top_in[15] ) , 
    .X ( chany_bottom_out[15] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_40__39 ( .A ( chany_top_in[19] ) , 
    .X ( aps_rename_2_ ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_57 ( .A ( chany_bottom_in[4] ) , 
    .X ( BUF_net_57 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_60 ( .A ( chany_bottom_in[10] ) , 
    .X ( BUF_net_60 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_RR_61 ( .A ( chany_bottom_in[13] ) , 
    .X ( chany_top_out[13] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_66 ( .A ( chany_top_in[5] ) , 
    .X ( BUF_net_66 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_68 ( .A ( chany_top_in[18] ) , 
    .X ( BUF_net_68 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 BUFT_RR_70 ( .A ( BUF_net_57 ) , 
    .X ( chany_top_out[4] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_RR_71 ( .A ( chany_bottom_in[7] ) , 
    .X ( chany_top_out[7] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 BUFT_RR_72 ( .A ( aps_rename_3_ ) , 
    .X ( chany_top_out[8] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 BUFT_RR_73 ( .A ( BUF_net_60 ) , 
    .X ( chany_top_out[10] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 BUFT_RR_74 ( .A ( aps_rename_4_ ) , 
    .X ( chany_top_out[14] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_RR_75 ( .A ( chany_bottom_in[17] ) , 
    .X ( chany_top_out[17] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 BUFT_RR_76 ( .A ( aps_rename_6_ ) , 
    .X ( chany_top_out[19] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 BUFT_RR_77 ( .A ( BUF_net_66 ) , 
    .X ( chany_bottom_out[5] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 BUFT_RR_79 ( .A ( aps_rename_2_ ) , 
    .X ( chany_bottom_out[19] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_P_83 ( .A ( chany_bottom_in[5] ) , 
    .X ( chany_top_out[5] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_P_84 ( .A ( chany_top_in[17] ) , 
    .X ( chany_bottom_out[17] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 BUFT_P_87 ( .A ( aps_rename_5_ ) , 
    .X ( chany_top_out[16] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_P_88 ( .A ( chany_top_in[16] ) , 
    .X ( chany_bottom_out[16] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 BUFT_P_91 ( .A ( BUF_net_68 ) , 
    .X ( chany_bottom_out[18] ) ) ;
endmodule


module mux_tree_tapbuf_size10_mem_15 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd1_1 FTB_2__41 ( .A ( mem_out[3] ) , 
    .X ( net_net_73 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_RR_110 ( .A ( net_net_73 ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size10_mem_0_4 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_1__40 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_43 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size10_15 ( in , sram , sram_inv , out , p0 ) ;
input  [0:9] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

const1_43 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[6] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[8] ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[9] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
endmodule


module const1_0_12 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size10_0_4 ( in , sram , sram_inv , out , p0 ) ;
input  [0:9] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

const1_0_12 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[6] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[8] ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[9] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
endmodule


module cby_0__1_ ( prog_clk , chany_bottom_in , chany_top_in , ccff_head , 
    chany_bottom_out , chany_top_out , right_grid_pin_52_ , left_grid_pin_0_ , 
    ccff_tail ) ;
input  [0:0] prog_clk ;
input  [0:19] chany_bottom_in ;
input  [0:19] chany_top_in ;
input  [0:0] ccff_head ;
output [0:19] chany_bottom_out ;
output [0:19] chany_top_out ;
output [0:0] right_grid_pin_52_ ;
output [0:0] left_grid_pin_0_ ;
output [0:0] ccff_tail ;

wire [0:3] mux_tree_tapbuf_size10_0_sram ;
wire [0:3] mux_tree_tapbuf_size10_0_sram_inv ;
wire [0:3] mux_tree_tapbuf_size10_1_sram ;
wire [0:3] mux_tree_tapbuf_size10_1_sram_inv ;
wire [0:0] mux_tree_tapbuf_size10_mem_0_ccff_tail ;

mux_tree_tapbuf_size10_0_4 mux_left_ipin_0 (
    .in ( { chany_bottom_in[0] , chany_top_in[0] , chany_bottom_in[2] , 
        chany_top_in[2] , chany_bottom_in[4] , chany_top_in[4] , 
        chany_bottom_in[10] , chany_top_in[10] , chany_bottom_in[16] , 
        chany_top_in[16] } ) ,
    .sram ( mux_tree_tapbuf_size10_0_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size10_0_sram_inv ) , 
    .out ( right_grid_pin_52_ ) , .p0 ( optlc_net_135 ) ) ;
mux_tree_tapbuf_size10_15 mux_right_ipin_0 (
    .in ( { chany_bottom_in[1] , chany_top_in[1] , chany_bottom_in[3] , 
        chany_top_in[3] , chany_bottom_in[5] , chany_top_in[5] , 
        chany_bottom_in[11] , chany_top_in[11] , chany_bottom_in[17] , 
        chany_top_in[17] } ) ,
    .sram ( mux_tree_tapbuf_size10_1_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size10_1_sram_inv ) , 
    .out ( left_grid_pin_0_ ) , .p0 ( optlc_net_135 ) ) ;
mux_tree_tapbuf_size10_mem_0_4 mem_left_ipin_0 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( ccff_head ) , 
    .ccff_tail ( mux_tree_tapbuf_size10_mem_0_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size10_0_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size10_0_sram_inv ) ) ;
mux_tree_tapbuf_size10_mem_15 mem_right_ipin_0 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size10_mem_0_ccff_tail ) ,
    .ccff_tail ( { ropt_net_161 } ) ,
    .mem_out ( mux_tree_tapbuf_size10_1_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size10_1_sram_inv ) ) ;
sky130_fd_sc_hd__conb_1 optlc_136 ( .LO ( SYNOPSYS_UNCONNECTED_1 ) , 
    .HI ( optlc_net_135 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_715 ( .A ( chany_bottom_in[8] ) , 
    .X ( ropt_net_181 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_3__2 ( .A ( chany_bottom_in[2] ) , 
    .X ( ropt_net_156 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_716 ( .A ( chany_bottom_in[1] ) , 
    .X ( ropt_net_200 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_717 ( .A ( ropt_net_138 ) , 
    .X ( ropt_net_182 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_718 ( .A ( chany_top_in[13] ) , 
    .X ( chany_bottom_out[13] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_753 ( .A ( ropt_net_174 ) , 
    .X ( chany_bottom_out[12] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_719 ( .A ( chany_top_in[9] ) , 
    .X ( chany_bottom_out[9] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_720 ( 
    .A ( chany_bottom_in[17] ) , .X ( ropt_net_203 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_721 ( 
    .A ( chany_bottom_in[16] ) , .X ( ropt_net_202 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_722 ( .A ( chany_bottom_in[6] ) , 
    .X ( ropt_net_199 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_723 ( .A ( chany_top_in[1] ) , 
    .X ( ropt_net_201 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_724 ( 
    .A ( chany_bottom_in[15] ) , .X ( ropt_net_177 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_725 ( .A ( chany_top_in[10] ) , 
    .X ( chany_bottom_out[10] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_726 ( .A ( ropt_net_147 ) , 
    .X ( ropt_net_180 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_727 ( .A ( ropt_net_148 ) , 
    .X ( ropt_net_185 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_754 ( .A ( ropt_net_175 ) , 
    .X ( chany_bottom_out[2] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_728 ( .A ( ropt_net_149 ) , 
    .X ( ropt_net_189 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_729 ( .A ( ropt_net_150 ) , 
    .X ( ropt_net_184 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_730 ( .A ( ropt_net_151 ) , 
    .X ( ropt_net_197 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_21__20 ( .A ( chany_top_in[0] ) , 
    .X ( ropt_net_168 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_731 ( .A ( ropt_net_152 ) , 
    .X ( ropt_net_195 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_732 ( .A ( ropt_net_153 ) , 
    .X ( ropt_net_174 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_733 ( .A ( ropt_net_154 ) , 
    .X ( ropt_net_194 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_734 ( .A ( ropt_net_155 ) , 
    .X ( ropt_net_176 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_26__25 ( .A ( chany_top_in[5] ) , 
    .X ( ropt_net_169 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_27__26 ( .A ( chany_top_in[6] ) , 
    .X ( aps_rename_1_ ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_735 ( .A ( ropt_net_156 ) , 
    .X ( ropt_net_178 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_736 ( .A ( ropt_net_157 ) , 
    .X ( ropt_net_179 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_737 ( .A ( ropt_net_158 ) , 
    .X ( ropt_net_192 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_738 ( .A ( ropt_net_159 ) , 
    .X ( ropt_net_188 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_32__31 ( .A ( chany_top_in[11] ) , 
    .X ( ropt_net_172 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_739 ( .A ( ropt_net_160 ) , 
    .X ( ropt_net_187 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_755 ( .A ( ropt_net_176 ) , 
    .X ( chany_bottom_out[15] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_740 ( .A ( ropt_net_161 ) , 
    .X ( ccff_tail[0] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_741 ( .A ( ropt_net_162 ) , 
    .X ( ropt_net_198 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_37__36 ( .A ( chany_top_in[16] ) , 
    .X ( chany_bottom_out[16] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_742 ( .A ( ropt_net_163 ) , 
    .X ( ropt_net_191 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_743 ( .A ( ropt_net_164 ) , 
    .X ( chany_bottom_out[17] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_744 ( .A ( ropt_net_165 ) , 
    .X ( ropt_net_183 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_745 ( .A ( ropt_net_166 ) , 
    .X ( chany_bottom_out[7] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_746 ( .A ( ropt_net_167 ) , 
    .X ( ropt_net_190 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_747 ( .A ( ropt_net_168 ) , 
    .X ( chany_bottom_out[0] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_748 ( .A ( ropt_net_169 ) , 
    .X ( ropt_net_186 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_749 ( .A ( ropt_net_170 ) , 
    .X ( ropt_net_193 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_756 ( .A ( ropt_net_177 ) , 
    .X ( chany_top_out[15] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_750 ( .A ( ropt_net_171 ) , 
    .X ( chany_bottom_out[19] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_757 ( .A ( ropt_net_178 ) , 
    .X ( chany_top_out[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_50 ( .A ( chany_bottom_in[9] ) , 
    .X ( ropt_net_151 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_51 ( .A ( chany_bottom_in[10] ) , 
    .X ( ropt_net_157 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_751 ( .A ( ropt_net_172 ) , 
    .X ( ropt_net_196 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_752 ( .A ( ropt_net_173 ) , 
    .X ( ropt_net_175 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_54 ( .A ( chany_bottom_in[13] ) , 
    .X ( ropt_net_147 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_758 ( .A ( ropt_net_179 ) , 
    .X ( chany_top_out[10] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_759 ( .A ( ropt_net_180 ) , 
    .X ( chany_top_out[13] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_760 ( .A ( ropt_net_181 ) , 
    .X ( chany_top_out[8] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_761 ( .A ( ropt_net_182 ) , 
    .X ( chany_bottom_out[18] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_59 ( .A ( chany_bottom_in[18] ) , 
    .X ( ropt_net_159 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_60 ( .A ( chany_bottom_in[19] ) , 
    .X ( ropt_net_167 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_762 ( .A ( ropt_net_183 ) , 
    .X ( chany_top_out[0] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_763 ( .A ( ropt_net_184 ) , 
    .X ( chany_bottom_out[3] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_765 ( .A ( ropt_net_185 ) , 
    .X ( chany_top_out[5] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_766 ( .A ( ropt_net_186 ) , 
    .X ( chany_bottom_out[5] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_767 ( .A ( ropt_net_187 ) , 
    .X ( chany_top_out[12] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_768 ( .A ( ropt_net_188 ) , 
    .X ( chany_top_out[18] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_769 ( .A ( ropt_net_189 ) , 
    .X ( chany_bottom_out[8] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_770 ( .A ( ropt_net_190 ) , 
    .X ( chany_top_out[19] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_771 ( .A ( ropt_net_191 ) , 
    .X ( chany_top_out[11] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_772 ( .A ( ropt_net_192 ) , 
    .X ( chany_top_out[3] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_773 ( .A ( ropt_net_193 ) , 
    .X ( chany_top_out[14] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_774 ( .A ( ropt_net_194 ) , 
    .X ( chany_bottom_out[14] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_775 ( .A ( ropt_net_195 ) , 
    .X ( chany_top_out[7] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_776 ( .A ( ropt_net_196 ) , 
    .X ( chany_bottom_out[11] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_777 ( .A ( ropt_net_197 ) , 
    .X ( chany_top_out[9] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_779 ( .A ( ropt_net_198 ) , 
    .X ( chany_bottom_out[4] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_78 ( .A ( chany_bottom_in[5] ) , 
    .X ( ropt_net_148 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_783 ( .A ( ropt_net_199 ) , 
    .X ( chany_top_out[6] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_784 ( .A ( ropt_net_200 ) , 
    .X ( chany_top_out[1] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_786 ( .A ( ropt_net_201 ) , 
    .X ( chany_bottom_out[1] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_787 ( .A ( ropt_net_202 ) , 
    .X ( chany_top_out[16] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_790 ( .A ( ropt_net_203 ) , 
    .X ( chany_top_out[17] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 BUFT_RR_92 ( .A ( aps_rename_1_ ) , 
    .X ( chany_bottom_out[6] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_P_101 ( .A ( chany_top_in[2] ) , 
    .X ( ropt_net_173 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_P_102 ( .A ( chany_top_in[4] ) , 
    .X ( ropt_net_162 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_P_103 ( .A ( chany_top_in[8] ) , 
    .X ( ropt_net_149 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_P_105 ( .A ( chany_top_in[17] ) , 
    .X ( ropt_net_164 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_P_108 ( .A ( chany_top_in[3] ) , 
    .X ( ropt_net_150 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_P_111 ( .A ( chany_bottom_in[0] ) , 
    .X ( ropt_net_165 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_P_113 ( .A ( chany_bottom_in[3] ) , 
    .X ( ropt_net_158 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_P_114 ( .A ( chany_bottom_in[4] ) , 
    .X ( chany_top_out[4] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_P_115 ( .A ( chany_bottom_in[7] ) , 
    .X ( ropt_net_152 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_P_118 ( .A ( chany_bottom_in[11] ) , 
    .X ( ropt_net_163 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_P_119 ( .A ( chany_bottom_in[12] ) , 
    .X ( ropt_net_160 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_P_121 ( .A ( chany_bottom_in[14] ) , 
    .X ( ropt_net_170 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_P_127 ( .A ( chany_top_in[7] ) , 
    .X ( ropt_net_166 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_P_129 ( .A ( chany_top_in[12] ) , 
    .X ( ropt_net_153 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_P_130 ( .A ( chany_top_in[14] ) , 
    .X ( ropt_net_154 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_P_131 ( .A ( chany_top_in[15] ) , 
    .X ( ropt_net_155 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_P_132 ( .A ( chany_top_in[18] ) , 
    .X ( ropt_net_138 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_P_133 ( .A ( chany_top_in[19] ) , 
    .X ( ropt_net_171 ) ) ;
endmodule


module mux_tree_tapbuf_size10_mem_14 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_1__40 ( .A ( mem_out[3] ) , 
    .X ( net_net_80 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_122 ( .A ( net_net_80 ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_42 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size10_14 ( in , sram , sram_inv , out , p0 ) ;
input  [0:9] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;

const1_42 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[6] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[8] ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[9] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_8 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .S ( sram[3] ) , .X ( out[0] ) ) ;
endmodule


module cbx_1__2_ ( prog_clk , chanx_left_in , chanx_right_in , ccff_head , 
    chanx_left_out , chanx_right_out , top_grid_pin_0_ , ccff_tail ) ;
input  [0:0] prog_clk ;
input  [0:19] chanx_left_in ;
input  [0:19] chanx_right_in ;
input  [0:0] ccff_head ;
output [0:19] chanx_left_out ;
output [0:19] chanx_right_out ;
output [0:0] top_grid_pin_0_ ;
output [0:0] ccff_tail ;

wire [0:3] mux_tree_tapbuf_size10_0_sram ;
wire [0:3] mux_tree_tapbuf_size10_0_sram_inv ;

mux_tree_tapbuf_size10_14 mux_bottom_ipin_0 (
    .in ( { chanx_left_in[0] , chanx_right_in[0] , chanx_left_in[2] , 
        chanx_right_in[2] , chanx_left_in[4] , chanx_right_in[4] , 
        chanx_left_in[10] , chanx_right_in[10] , chanx_left_in[16] , 
        chanx_right_in[16] } ) ,
    .sram ( mux_tree_tapbuf_size10_0_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size10_0_sram_inv ) , 
    .out ( top_grid_pin_0_ ) , .p0 ( optlc_net_159 ) ) ;
mux_tree_tapbuf_size10_mem_14 mem_bottom_ipin_0 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( ccff_head ) ,
    .ccff_tail ( { ropt_net_165 } ) ,
    .mem_out ( mux_tree_tapbuf_size10_0_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size10_0_sram_inv ) ) ;
sky130_fd_sc_hd__conb_1 optlc_160 ( .LO ( SYNOPSYS_UNCONNECTED_1 ) , 
    .HI ( optlc_net_159 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_739 ( .A ( chanx_right_in[14] ) , 
    .X ( ropt_net_219 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_740 ( .A ( chanx_right_in[11] ) , 
    .X ( ropt_net_214 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_741 ( .A ( chanx_right_in[5] ) , 
    .X ( chanx_left_out[5] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_742 ( .A ( chanx_right_in[18] ) , 
    .X ( ropt_net_220 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_743 ( .A ( ropt_net_165 ) , 
    .X ( ropt_net_215 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_744 ( .A ( chanx_right_in[9] ) , 
    .X ( ropt_net_222 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_745 ( .A ( chanx_left_in[14] ) , 
    .X ( ropt_net_212 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_746 ( .A ( chanx_left_in[15] ) , 
    .X ( ropt_net_210 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_747 ( .A ( chanx_right_in[17] ) , 
    .X ( ropt_net_223 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_748 ( .A ( chanx_right_in[12] ) , 
    .X ( ropt_net_218 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_749 ( .A ( chanx_right_in[1] ) , 
    .X ( ropt_net_213 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_750 ( .A ( chanx_right_in[2] ) , 
    .X ( chanx_left_out[2] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_751 ( .A ( chanx_left_in[11] ) , 
    .X ( ropt_net_221 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_752 ( .A ( chanx_right_in[6] ) , 
    .X ( ropt_net_217 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_753 ( .A ( chanx_left_in[12] ) , 
    .X ( ropt_net_225 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_754 ( .A ( chanx_left_in[13] ) , 
    .X ( ropt_net_224 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_755 ( .A ( chanx_right_in[13] ) , 
    .X ( ropt_net_216 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_756 ( .A ( chanx_left_in[7] ) , 
    .X ( chanx_right_out[7] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_757 ( .A ( chanx_left_in[19] ) , 
    .X ( chanx_right_out[19] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_758 ( .A ( ropt_net_180 ) , 
    .X ( ropt_net_205 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_759 ( .A ( chanx_right_in[19] ) , 
    .X ( ropt_net_211 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_760 ( .A ( ropt_net_182 ) , 
    .X ( ropt_net_209 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_761 ( .A ( ropt_net_183 ) , 
    .X ( chanx_right_out[5] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_762 ( .A ( ropt_net_184 ) , 
    .X ( ropt_net_201 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_763 ( .A ( ropt_net_185 ) , 
    .X ( chanx_right_out[3] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_764 ( .A ( ropt_net_186 ) , 
    .X ( ropt_net_198 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_765 ( .A ( ropt_net_187 ) , 
    .X ( ropt_net_206 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_766 ( .A ( ropt_net_188 ) , 
    .X ( ropt_net_208 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_767 ( .A ( ropt_net_189 ) , 
    .X ( chanx_right_out[9] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_768 ( .A ( ropt_net_190 ) , 
    .X ( chanx_right_out[6] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_769 ( .A ( ropt_net_191 ) , 
    .X ( ropt_net_199 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_770 ( .A ( ropt_net_192 ) , 
    .X ( ropt_net_202 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_771 ( .A ( ropt_net_193 ) , 
    .X ( ropt_net_200 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_772 ( .A ( ropt_net_194 ) , 
    .X ( ropt_net_207 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_773 ( .A ( ropt_net_195 ) , 
    .X ( chanx_left_out[0] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_774 ( .A ( ropt_net_196 ) , 
    .X ( chanx_right_out[2] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_776 ( .A ( ropt_net_198 ) , 
    .X ( chanx_left_out[10] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_775 ( .A ( ropt_net_197 ) , 
    .X ( ropt_net_204 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_777 ( .A ( ropt_net_199 ) , 
    .X ( chanx_left_out[16] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_778 ( .A ( ropt_net_200 ) , 
    .X ( chanx_left_out[4] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_779 ( .A ( ropt_net_201 ) , 
    .X ( chanx_left_out[8] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_780 ( .A ( ropt_net_202 ) , 
    .X ( chanx_left_out[7] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_781 ( .A ( ropt_net_203 ) , 
    .X ( chanx_right_out[17] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_46 ( .A ( chanx_left_in[4] ) , 
    .X ( BUF_net_46 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_782 ( .A ( ropt_net_204 ) , 
    .X ( chanx_left_out[3] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_784 ( .A ( ropt_net_205 ) , 
    .X ( chanx_right_out[18] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_785 ( .A ( ropt_net_206 ) , 
    .X ( chanx_right_out[0] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_786 ( .A ( ropt_net_207 ) , 
    .X ( chanx_right_out[8] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_787 ( .A ( ropt_net_208 ) , 
    .X ( chanx_right_out[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_52 ( .A ( chanx_left_in[10] ) , 
    .X ( BUF_net_52 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_788 ( .A ( ropt_net_209 ) , 
    .X ( chanx_right_out[16] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_791 ( .A ( ropt_net_210 ) , 
    .X ( chanx_right_out[15] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_792 ( .A ( ropt_net_211 ) , 
    .X ( chanx_left_out[19] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_794 ( .A ( ropt_net_212 ) , 
    .X ( chanx_right_out[14] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_795 ( .A ( ropt_net_213 ) , 
    .X ( chanx_left_out[1] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_796 ( .A ( ropt_net_214 ) , 
    .X ( chanx_left_out[11] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_59 ( .A ( chanx_left_in[17] ) , 
    .X ( BUF_net_59 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_797 ( .A ( ropt_net_215 ) , 
    .X ( ccff_tail[0] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_799 ( .A ( ropt_net_216 ) , 
    .X ( chanx_left_out[13] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_RR_62 ( .A ( chanx_right_in[0] ) , 
    .X ( ropt_net_195 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_800 ( .A ( ropt_net_217 ) , 
    .X ( chanx_left_out[6] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_801 ( .A ( ropt_net_218 ) , 
    .X ( chanx_left_out[12] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_802 ( .A ( ropt_net_219 ) , 
    .X ( chanx_left_out[14] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_804 ( .A ( ropt_net_220 ) , 
    .X ( chanx_left_out[18] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_805 ( .A ( ropt_net_221 ) , 
    .X ( chanx_right_out[11] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_68 ( .A ( chanx_right_in[7] ) , 
    .X ( ropt_net_192 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_806 ( .A ( ropt_net_222 ) , 
    .X ( chanx_left_out[9] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_808 ( .A ( ropt_net_223 ) , 
    .X ( chanx_left_out[17] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_71 ( .A ( chanx_right_in[10] ) , 
    .X ( ropt_net_186 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_810 ( .A ( ropt_net_224 ) , 
    .X ( chanx_right_out[13] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_811 ( .A ( ropt_net_225 ) , 
    .X ( chanx_right_out[12] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_76 ( .A ( chanx_right_in[15] ) , 
    .X ( BUF_net_76 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_P_117 ( .A ( chanx_right_in[3] ) , 
    .X ( ropt_net_197 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_P_118 ( .A ( chanx_right_in[16] ) , 
    .X ( ropt_net_191 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_P_124 ( .A ( chanx_left_in[0] ) , 
    .X ( ropt_net_187 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_P_125 ( .A ( chanx_left_in[1] ) , 
    .X ( ropt_net_188 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_P_126 ( .A ( chanx_left_in[2] ) , 
    .X ( ropt_net_196 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_P_127 ( .A ( chanx_left_in[3] ) , 
    .X ( ropt_net_185 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 BUFT_P_128 ( .A ( BUF_net_46 ) , 
    .X ( chanx_right_out[4] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_P_129 ( .A ( chanx_left_in[5] ) , 
    .X ( ropt_net_183 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_P_130 ( .A ( chanx_left_in[6] ) , 
    .X ( ropt_net_190 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_P_132 ( .A ( chanx_left_in[8] ) , 
    .X ( ropt_net_194 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_P_133 ( .A ( chanx_left_in[9] ) , 
    .X ( ropt_net_189 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 BUFT_P_134 ( .A ( BUF_net_52 ) , 
    .X ( chanx_right_out[10] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_P_140 ( .A ( chanx_left_in[16] ) , 
    .X ( ropt_net_182 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 BUFT_P_141 ( .A ( BUF_net_59 ) , 
    .X ( ropt_net_203 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_P_142 ( .A ( chanx_left_in[18] ) , 
    .X ( ropt_net_180 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_P_146 ( .A ( chanx_right_in[4] ) , 
    .X ( ropt_net_193 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_P_149 ( .A ( chanx_right_in[8] ) , 
    .X ( ropt_net_184 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 BUFT_P_156 ( .A ( BUF_net_76 ) , 
    .X ( chanx_left_out[15] ) ) ;
endmodule


module mux_tree_tapbuf_size8_mem_3_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_16__55 ( .A ( mem_out[3] ) , 
    .X ( net_net_74 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_RR_73 ( .A ( net_net_73 ) , 
    .X ( ccff_tail[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd1_1 BUFT_RR_74 ( .A ( net_net_74 ) , 
    .X ( net_net_73 ) ) ;
endmodule


module mux_tree_tapbuf_size8_mem_2_2 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_15__54 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size8_mem_1_3 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_14__53 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size8_mem_0_3 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_13__52 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size8_mem_8 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_12__51 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size8_mem_6_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_11__50 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size8_mem_5_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_10__49 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size8_mem_4_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_9__48 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_41 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size8_3_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:7] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;

const1_41 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( in[2] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[4] ) , .A1 ( in[3] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[6] ) , .A1 ( in[5] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_4 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[3] ) , .X ( out[0] ) ) ;
endmodule


module const1_14_10 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size8_2_2 ( in , sram , sram_inv , out , p0 ) ;
input  [0:7] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;

const1_14_10 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( in[2] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[4] ) , .A1 ( in[3] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[6] ) , .A1 ( in[5] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
endmodule


module const1_13_10 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size8_1_3 ( in , sram , sram_inv , out , p0 ) ;
input  [0:7] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;

const1_13_10 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( in[2] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[4] ) , .A1 ( in[3] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[6] ) , .A1 ( in[5] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
endmodule


module const1_12_10 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size8_0_3 ( in , sram , sram_inv , out , p0 ) ;
input  [0:7] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;

const1_12_10 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( in[2] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[4] ) , .A1 ( in[3] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[6] ) , .A1 ( in[5] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
endmodule


module const1_11_10 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size8_8 ( in , sram , sram_inv , out , p0 ) ;
input  [0:7] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;

const1_11_10 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( in[2] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[4] ) , .A1 ( in[3] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[6] ) , .A1 ( in[5] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_4 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[3] ) , .X ( out[0] ) ) ;
endmodule


module const1_10_10 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size8_6_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:7] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;

const1_10_10 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( in[2] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[4] ) , .A1 ( in[3] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[6] ) , .A1 ( in[5] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
endmodule


module const1_9_10 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size8_5_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:7] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;

const1_9_10 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( in[2] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[4] ) , .A1 ( in[3] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[6] ) , .A1 ( in[5] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
endmodule


module const1_8_10 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size8_4_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:7] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;

const1_8_10 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( in[2] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[4] ) , .A1 ( in[3] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[6] ) , .A1 ( in[5] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
endmodule


module mux_tree_tapbuf_size10_mem_3_2 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_8__47 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size10_mem_2_2 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_7__46 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size10_mem_13 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_6__45 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size10_mem_6_2 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_5__44 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size10_mem_5_2 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_4__43 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size10_mem_4_2 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_3__42 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size10_mem_1_2 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_2__41 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size10_mem_0_3 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_1__40 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_7_10 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size10_3_2 ( in , sram , sram_inv , out , p0 ) ;
input  [0:9] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

const1_7_10 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[6] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[8] ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[9] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
endmodule


module const1_6_11 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size10_2_2 ( in , sram , sram_inv , out , p0 ) ;
input  [0:9] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

const1_6_11 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[6] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[8] ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[9] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
endmodule


module const1_5_11 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size10_13 ( in , sram , sram_inv , out , p0 ) ;
input  [0:9] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

const1_5_11 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[6] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[8] ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[9] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
endmodule


module const1_4_11 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size10_6_2 ( in , sram , sram_inv , out , p0 ) ;
input  [0:9] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

const1_4_11 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[6] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[8] ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[9] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
endmodule


module const1_3_11 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size10_5_2 ( in , sram , sram_inv , out , p0 ) ;
input  [0:9] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

const1_3_11 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[6] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[8] ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[9] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
endmodule


module const1_2_11 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size10_4_2 ( in , sram , sram_inv , out , p0 ) ;
input  [0:9] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

const1_2_11 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[6] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[8] ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[9] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
endmodule


module const1_1_11 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size10_1_2 ( in , sram , sram_inv , out , p0 ) ;
input  [0:9] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

const1_1_11 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[6] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[8] ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[9] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
endmodule


module const1_0_11 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size10_0_3 ( in , sram , sram_inv , out , p0 ) ;
input  [0:9] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

const1_0_11 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[6] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[8] ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[9] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
endmodule


module cbx_1__1_ ( prog_clk , chanx_left_in , chanx_right_in , ccff_head , 
    chanx_left_out , chanx_right_out , top_grid_pin_16_ , top_grid_pin_17_ , 
    top_grid_pin_18_ , top_grid_pin_19_ , top_grid_pin_20_ , 
    top_grid_pin_21_ , top_grid_pin_22_ , top_grid_pin_23_ , 
    top_grid_pin_24_ , top_grid_pin_25_ , top_grid_pin_26_ , 
    top_grid_pin_27_ , top_grid_pin_28_ , top_grid_pin_29_ , 
    top_grid_pin_30_ , top_grid_pin_31_ , ccff_tail ) ;
input  [0:0] prog_clk ;
input  [0:19] chanx_left_in ;
input  [0:19] chanx_right_in ;
input  [0:0] ccff_head ;
output [0:19] chanx_left_out ;
output [0:19] chanx_right_out ;
output [0:0] top_grid_pin_16_ ;
output [0:0] top_grid_pin_17_ ;
output [0:0] top_grid_pin_18_ ;
output [0:0] top_grid_pin_19_ ;
output [0:0] top_grid_pin_20_ ;
output [0:0] top_grid_pin_21_ ;
output [0:0] top_grid_pin_22_ ;
output [0:0] top_grid_pin_23_ ;
output [0:0] top_grid_pin_24_ ;
output [0:0] top_grid_pin_25_ ;
output [0:0] top_grid_pin_26_ ;
output [0:0] top_grid_pin_27_ ;
output [0:0] top_grid_pin_28_ ;
output [0:0] top_grid_pin_29_ ;
output [0:0] top_grid_pin_30_ ;
output [0:0] top_grid_pin_31_ ;
output [0:0] ccff_tail ;

wire [0:3] mux_tree_tapbuf_size10_0_sram ;
wire [0:3] mux_tree_tapbuf_size10_0_sram_inv ;
wire [0:3] mux_tree_tapbuf_size10_1_sram ;
wire [0:3] mux_tree_tapbuf_size10_1_sram_inv ;
wire [0:3] mux_tree_tapbuf_size10_2_sram ;
wire [0:3] mux_tree_tapbuf_size10_2_sram_inv ;
wire [0:3] mux_tree_tapbuf_size10_3_sram ;
wire [0:3] mux_tree_tapbuf_size10_3_sram_inv ;
wire [0:3] mux_tree_tapbuf_size10_4_sram ;
wire [0:3] mux_tree_tapbuf_size10_4_sram_inv ;
wire [0:3] mux_tree_tapbuf_size10_5_sram ;
wire [0:3] mux_tree_tapbuf_size10_5_sram_inv ;
wire [0:3] mux_tree_tapbuf_size10_6_sram ;
wire [0:3] mux_tree_tapbuf_size10_6_sram_inv ;
wire [0:3] mux_tree_tapbuf_size10_7_sram ;
wire [0:3] mux_tree_tapbuf_size10_7_sram_inv ;
wire [0:0] mux_tree_tapbuf_size10_mem_0_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size10_mem_1_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size10_mem_2_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size10_mem_3_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size10_mem_4_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size10_mem_5_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size10_mem_6_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size10_mem_7_ccff_tail ;
wire [0:3] mux_tree_tapbuf_size8_0_sram ;
wire [0:3] mux_tree_tapbuf_size8_0_sram_inv ;
wire [0:3] mux_tree_tapbuf_size8_1_sram ;
wire [0:3] mux_tree_tapbuf_size8_1_sram_inv ;
wire [0:3] mux_tree_tapbuf_size8_2_sram ;
wire [0:3] mux_tree_tapbuf_size8_2_sram_inv ;
wire [0:3] mux_tree_tapbuf_size8_3_sram ;
wire [0:3] mux_tree_tapbuf_size8_3_sram_inv ;
wire [0:3] mux_tree_tapbuf_size8_4_sram ;
wire [0:3] mux_tree_tapbuf_size8_4_sram_inv ;
wire [0:3] mux_tree_tapbuf_size8_5_sram ;
wire [0:3] mux_tree_tapbuf_size8_5_sram_inv ;
wire [0:3] mux_tree_tapbuf_size8_6_sram ;
wire [0:3] mux_tree_tapbuf_size8_6_sram_inv ;
wire [0:3] mux_tree_tapbuf_size8_7_sram ;
wire [0:3] mux_tree_tapbuf_size8_7_sram_inv ;
wire [0:0] mux_tree_tapbuf_size8_mem_0_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size8_mem_1_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size8_mem_2_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size8_mem_3_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size8_mem_4_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size8_mem_5_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size8_mem_6_ccff_tail ;

mux_tree_tapbuf_size10_0_3 mux_bottom_ipin_0 (
    .in ( { chanx_left_in[0] , chanx_right_in[0] , chanx_left_in[2] , 
        chanx_right_in[2] , chanx_left_in[4] , chanx_right_in[4] , 
        chanx_left_in[10] , chanx_right_in[10] , chanx_left_in[16] , 
        chanx_right_in[16] } ) ,
    .sram ( mux_tree_tapbuf_size10_0_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size10_0_sram_inv ) , 
    .out ( top_grid_pin_16_ ) , .p0 ( optlc_net_108 ) ) ;
mux_tree_tapbuf_size10_1_2 mux_bottom_ipin_1 (
    .in ( { chanx_left_in[1] , chanx_right_in[1] , chanx_left_in[3] , 
        chanx_right_in[3] , chanx_left_in[5] , chanx_right_in[5] , 
        chanx_left_in[11] , chanx_right_in[11] , chanx_left_in[17] , 
        chanx_right_in[17] } ) ,
    .sram ( mux_tree_tapbuf_size10_1_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size10_1_sram_inv ) , 
    .out ( top_grid_pin_17_ ) , .p0 ( optlc_net_109 ) ) ;
mux_tree_tapbuf_size10_4_2 mux_bottom_ipin_4 (
    .in ( { chanx_left_in[0] , chanx_right_in[0] , chanx_left_in[2] , 
        chanx_right_in[2] , chanx_left_in[4] , chanx_right_in[4] , 
        chanx_left_in[8] , chanx_right_in[8] , chanx_left_in[14] , 
        chanx_right_in[14] } ) ,
    .sram ( mux_tree_tapbuf_size10_2_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size10_2_sram_inv ) , 
    .out ( top_grid_pin_20_ ) , .p0 ( optlc_net_108 ) ) ;
mux_tree_tapbuf_size10_5_2 mux_bottom_ipin_5 (
    .in ( { chanx_left_in[1] , chanx_right_in[1] , chanx_left_in[3] , 
        chanx_right_in[3] , chanx_left_in[5] , chanx_right_in[5] , 
        chanx_left_in[9] , chanx_right_in[9] , chanx_left_in[15] , 
        chanx_right_in[15] } ) ,
    .sram ( mux_tree_tapbuf_size10_3_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size10_3_sram_inv ) , 
    .out ( top_grid_pin_21_ ) , .p0 ( optlc_net_109 ) ) ;
mux_tree_tapbuf_size10_6_2 mux_bottom_ipin_8 (
    .in ( { chanx_left_in[0] , chanx_right_in[0] , chanx_left_in[2] , 
        chanx_right_in[2] , chanx_left_in[8] , chanx_right_in[8] , 
        chanx_left_in[12] , chanx_right_in[12] , chanx_left_in[18] , 
        chanx_right_in[18] } ) ,
    .sram ( mux_tree_tapbuf_size10_4_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size10_4_sram_inv ) , 
    .out ( top_grid_pin_24_ ) , .p0 ( optlc_net_109 ) ) ;
mux_tree_tapbuf_size10_13 mux_bottom_ipin_9 (
    .in ( { chanx_left_in[1] , chanx_right_in[1] , chanx_left_in[3] , 
        chanx_right_in[3] , chanx_left_in[9] , chanx_right_in[9] , 
        chanx_left_in[13] , chanx_right_in[13] , chanx_left_in[19] , 
        chanx_right_in[19] } ) ,
    .sram ( mux_tree_tapbuf_size10_5_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size10_5_sram_inv ) , 
    .out ( top_grid_pin_25_ ) , .p0 ( optlc_net_108 ) ) ;
mux_tree_tapbuf_size10_2_2 mux_bottom_ipin_12 (
    .in ( { chanx_left_in[0] , chanx_right_in[0] , chanx_left_in[2] , 
        chanx_right_in[2] , chanx_left_in[6] , chanx_right_in[6] , 
        chanx_left_in[12] , chanx_right_in[12] , chanx_left_in[16] , 
        chanx_right_in[16] } ) ,
    .sram ( mux_tree_tapbuf_size10_6_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size10_6_sram_inv ) , 
    .out ( top_grid_pin_28_ ) , .p0 ( optlc_net_109 ) ) ;
mux_tree_tapbuf_size10_3_2 mux_bottom_ipin_13 (
    .in ( { chanx_left_in[1] , chanx_right_in[1] , chanx_left_in[3] , 
        chanx_right_in[3] , chanx_left_in[7] , chanx_right_in[7] , 
        chanx_left_in[13] , chanx_right_in[13] , chanx_left_in[17] , 
        chanx_right_in[17] } ) ,
    .sram ( mux_tree_tapbuf_size10_7_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size10_7_sram_inv ) , 
    .out ( top_grid_pin_29_ ) , .p0 ( optlc_net_109 ) ) ;
mux_tree_tapbuf_size10_mem_0_3 mem_bottom_ipin_0 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( ccff_head ) , 
    .ccff_tail ( mux_tree_tapbuf_size10_mem_0_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size10_0_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size10_0_sram_inv ) ) ;
mux_tree_tapbuf_size10_mem_1_2 mem_bottom_ipin_1 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size10_mem_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size10_mem_1_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size10_1_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size10_1_sram_inv ) ) ;
mux_tree_tapbuf_size10_mem_4_2 mem_bottom_ipin_4 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size8_mem_1_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size10_mem_2_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size10_2_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size10_2_sram_inv ) ) ;
mux_tree_tapbuf_size10_mem_5_2 mem_bottom_ipin_5 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size10_mem_2_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size10_mem_3_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size10_3_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size10_3_sram_inv ) ) ;
mux_tree_tapbuf_size10_mem_6_2 mem_bottom_ipin_8 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size8_mem_3_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size10_mem_4_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size10_4_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size10_4_sram_inv ) ) ;
mux_tree_tapbuf_size10_mem_13 mem_bottom_ipin_9 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size10_mem_4_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size10_mem_5_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size10_5_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size10_5_sram_inv ) ) ;
mux_tree_tapbuf_size10_mem_2_2 mem_bottom_ipin_12 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size8_mem_5_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size10_mem_6_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size10_6_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size10_6_sram_inv ) ) ;
mux_tree_tapbuf_size10_mem_3_2 mem_bottom_ipin_13 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size10_mem_6_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size10_mem_7_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size10_7_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size10_7_sram_inv ) ) ;
mux_tree_tapbuf_size8_4_1 mux_bottom_ipin_2 (
    .in ( { chanx_left_in[0] , chanx_right_in[0] , chanx_left_in[2] , 
        chanx_right_in[2] , chanx_left_in[6] , chanx_right_in[6] , 
        chanx_left_in[14] , chanx_right_in[14] } ) ,
    .sram ( mux_tree_tapbuf_size8_0_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size8_0_sram_inv ) , 
    .out ( top_grid_pin_18_ ) , .p0 ( optlc_net_109 ) ) ;
mux_tree_tapbuf_size8_5_1 mux_bottom_ipin_3 (
    .in ( { chanx_left_in[1] , chanx_right_in[1] , chanx_left_in[3] , 
        chanx_right_in[3] , chanx_left_in[7] , chanx_right_in[7] , 
        chanx_left_in[15] , chanx_right_in[15] } ) ,
    .sram ( mux_tree_tapbuf_size8_1_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size8_1_sram_inv ) , 
    .out ( top_grid_pin_19_ ) , .p0 ( optlc_net_109 ) ) ;
mux_tree_tapbuf_size8_6_1 mux_bottom_ipin_6 (
    .in ( { chanx_left_in[0] , chanx_right_in[0] , chanx_left_in[2] , 
        chanx_right_in[2] , chanx_left_in[10] , chanx_right_in[10] , 
        chanx_left_in[18] , chanx_right_in[18] } ) ,
    .sram ( mux_tree_tapbuf_size8_2_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size8_2_sram_inv ) , 
    .out ( top_grid_pin_22_ ) , .p0 ( optlc_net_108 ) ) ;
mux_tree_tapbuf_size8_8 mux_bottom_ipin_7 (
    .in ( { chanx_left_in[1] , chanx_right_in[1] , chanx_left_in[3] , 
        chanx_right_in[3] , chanx_left_in[11] , chanx_right_in[11] , 
        chanx_left_in[19] , chanx_right_in[19] } ) ,
    .sram ( mux_tree_tapbuf_size8_3_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size8_3_sram_inv ) , 
    .out ( top_grid_pin_23_ ) , .p0 ( optlc_net_109 ) ) ;
mux_tree_tapbuf_size8_0_3 mux_bottom_ipin_10 (
    .in ( { chanx_left_in[0] , chanx_right_in[0] , chanx_left_in[2] , 
        chanx_right_in[2] , chanx_left_in[6] , chanx_right_in[6] , 
        chanx_left_in[14] , chanx_right_in[14] } ) ,
    .sram ( mux_tree_tapbuf_size8_4_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size8_4_sram_inv ) , 
    .out ( top_grid_pin_26_ ) , .p0 ( optlc_net_108 ) ) ;
mux_tree_tapbuf_size8_1_3 mux_bottom_ipin_11 (
    .in ( { chanx_left_in[1] , chanx_right_in[1] , chanx_left_in[3] , 
        chanx_right_in[3] , chanx_left_in[7] , chanx_right_in[7] , 
        chanx_left_in[15] , chanx_right_in[15] } ) ,
    .sram ( mux_tree_tapbuf_size8_5_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size8_5_sram_inv ) , 
    .out ( top_grid_pin_27_ ) , .p0 ( optlc_net_108 ) ) ;
mux_tree_tapbuf_size8_2_2 mux_bottom_ipin_14 (
    .in ( { chanx_left_in[0] , chanx_right_in[0] , chanx_left_in[2] , 
        chanx_right_in[2] , chanx_left_in[10] , chanx_right_in[10] , 
        chanx_left_in[18] , chanx_right_in[18] } ) ,
    .sram ( mux_tree_tapbuf_size8_6_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size8_6_sram_inv ) , 
    .out ( top_grid_pin_30_ ) , .p0 ( optlc_net_109 ) ) ;
mux_tree_tapbuf_size8_3_1 mux_bottom_ipin_15 (
    .in ( { chanx_left_in[1] , chanx_right_in[1] , chanx_left_in[3] , 
        chanx_right_in[3] , chanx_left_in[11] , chanx_right_in[11] , 
        chanx_left_in[19] , chanx_right_in[19] } ) ,
    .sram ( mux_tree_tapbuf_size8_7_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size8_7_sram_inv ) , 
    .out ( top_grid_pin_31_ ) , .p0 ( optlc_net_109 ) ) ;
mux_tree_tapbuf_size8_mem_4_1 mem_bottom_ipin_2 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size10_mem_1_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size8_mem_0_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size8_0_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size8_0_sram_inv ) ) ;
mux_tree_tapbuf_size8_mem_5_1 mem_bottom_ipin_3 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size8_mem_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size8_mem_1_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size8_1_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size8_1_sram_inv ) ) ;
mux_tree_tapbuf_size8_mem_6_1 mem_bottom_ipin_6 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size10_mem_3_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size8_mem_2_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size8_2_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size8_2_sram_inv ) ) ;
mux_tree_tapbuf_size8_mem_8 mem_bottom_ipin_7 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size8_mem_2_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size8_mem_3_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size8_3_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size8_3_sram_inv ) ) ;
mux_tree_tapbuf_size8_mem_0_3 mem_bottom_ipin_10 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size10_mem_5_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size8_mem_4_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size8_4_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size8_4_sram_inv ) ) ;
mux_tree_tapbuf_size8_mem_1_3 mem_bottom_ipin_11 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size8_mem_4_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size8_mem_5_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size8_5_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size8_5_sram_inv ) ) ;
mux_tree_tapbuf_size8_mem_2_2 mem_bottom_ipin_14 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size10_mem_7_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size8_mem_6_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size8_6_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size8_6_sram_inv ) ) ;
mux_tree_tapbuf_size8_mem_3_1 mem_bottom_ipin_15 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size8_mem_6_ccff_tail ) , 
    .ccff_tail ( ccff_tail ) , .mem_out ( mux_tree_tapbuf_size8_7_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size8_7_sram_inv ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_1__0 ( .A ( chanx_left_in[0] ) , 
    .X ( chanx_right_out[0] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_2__1 ( .A ( chanx_left_in[1] ) , 
    .X ( chanx_right_out[1] ) ) ;
sky130_fd_sc_hd__conb_1 optlc_102 ( .LO ( SYNOPSYS_UNCONNECTED_1 ) , 
    .HI ( optlc_net_108 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_104 ( .LO ( SYNOPSYS_UNCONNECTED_2 ) , 
    .HI ( optlc_net_109 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_684 ( .A ( chanx_right_in[12] ) , 
    .X ( chanx_left_out[12] ) ) ;
sky130_fd_sc_hd__dlygate4sd1_1 FTB_6__5 ( .A ( chanx_left_in[5] ) , 
    .X ( chanx_right_out[5] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_703 ( .A ( ropt_net_117 ) , 
    .X ( chanx_right_out[4] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_687 ( .A ( chanx_left_in[10] ) , 
    .X ( chanx_right_out[10] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_689 ( .A ( ropt_net_112 ) , 
    .X ( ropt_net_117 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_10__9 ( .A ( chanx_left_in[9] ) , 
    .X ( chanx_right_out[9] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_690 ( .A ( chanx_left_in[6] ) , 
    .X ( chanx_right_out[6] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_692 ( .A ( ropt_net_114 ) , 
    .X ( ropt_net_118 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_13__12 ( .A ( chanx_left_in[12] ) , 
    .X ( ropt_net_115 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_14__13 ( .A ( chanx_left_in[13] ) , 
    .X ( chanx_right_out[13] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_15__14 ( .A ( chanx_left_in[14] ) , 
    .X ( ropt_net_116 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_16__15 ( .A ( chanx_left_in[15] ) , 
    .X ( chanx_right_out[15] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_694 ( .A ( ropt_net_115 ) , 
    .X ( ropt_net_119 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_699 ( .A ( ropt_net_116 ) , 
    .X ( ropt_net_120 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_704 ( .A ( ropt_net_118 ) , 
    .X ( chanx_left_out[2] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_20__19 ( .A ( chanx_left_in[19] ) , 
    .X ( chanx_right_out[19] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_21__20 ( .A ( chanx_right_in[0] ) , 
    .X ( aps_rename_1_ ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_705 ( .A ( ropt_net_119 ) , 
    .X ( chanx_right_out[12] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_706 ( .A ( ropt_net_120 ) , 
    .X ( chanx_right_out[14] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_24__23 ( .A ( chanx_right_in[3] ) , 
    .X ( chanx_left_out[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_25__24 ( .A ( chanx_right_in[4] ) , 
    .X ( aps_rename_2_ ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_26__25 ( .A ( chanx_right_in[5] ) , 
    .X ( aps_rename_3_ ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_709 ( .A ( ropt_net_121 ) , 
    .X ( chanx_right_out[17] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_28__27 ( .A ( chanx_right_in[7] ) , 
    .X ( chanx_left_out[7] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_31__30 ( .A ( chanx_right_in[10] ) , 
    .X ( chanx_left_out[10] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_32__31 ( .A ( chanx_right_in[11] ) , 
    .X ( chanx_left_out[11] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_34__33 ( .A ( chanx_right_in[13] ) , 
    .X ( chanx_left_out[13] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_36__35 ( .A ( chanx_right_in[15] ) , 
    .X ( chanx_left_out[15] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_38__37 ( .A ( chanx_right_in[17] ) , 
    .X ( chanx_left_out[17] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_40__39 ( .A ( chanx_right_in[19] ) , 
    .X ( chanx_left_out[19] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_RR_61 ( .A ( chanx_left_in[7] ) , 
    .X ( chanx_right_out[7] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_RR_63 ( .A ( chanx_left_in[11] ) , 
    .X ( chanx_right_out[11] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_67 ( .A ( chanx_right_in[2] ) , 
    .X ( ropt_net_114 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_71 ( .A ( chanx_right_in[16] ) , 
    .X ( BUF_net_71 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_76 ( .A ( chanx_left_in[4] ) , 
    .X ( ropt_net_112 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_RR_77 ( .A ( chanx_left_in[8] ) , 
    .X ( chanx_right_out[8] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_RR_78 ( .A ( chanx_left_in[17] ) , 
    .X ( ropt_net_121 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_RR_79 ( .A ( chanx_right_in[8] ) , 
    .X ( chanx_left_out[8] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_RR_83 ( .A ( chanx_left_in[16] ) , 
    .X ( chanx_right_out[16] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_RR_84 ( .A ( chanx_left_in[18] ) , 
    .X ( chanx_right_out[18] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 BUFT_RR_85 ( .A ( aps_rename_1_ ) , 
    .X ( chanx_left_out[0] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 BUFT_RR_86 ( .A ( aps_rename_2_ ) , 
    .X ( chanx_left_out[4] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 BUFT_RR_87 ( .A ( aps_rename_3_ ) , 
    .X ( chanx_left_out[5] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_P_90 ( .A ( chanx_left_in[2] ) , 
    .X ( chanx_right_out[2] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_P_91 ( .A ( chanx_left_in[3] ) , 
    .X ( chanx_right_out[3] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_P_92 ( .A ( chanx_right_in[1] ) , 
    .X ( chanx_left_out[1] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_P_93 ( .A ( chanx_right_in[6] ) , 
    .X ( chanx_left_out[6] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_P_94 ( .A ( chanx_right_in[9] ) , 
    .X ( chanx_left_out[9] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_P_95 ( .A ( chanx_right_in[14] ) , 
    .X ( chanx_left_out[14] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 BUFT_P_97 ( .A ( BUF_net_71 ) , 
    .X ( chanx_left_out[16] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_P_98 ( .A ( chanx_right_in[18] ) , 
    .X ( chanx_left_out[18] ) ) ;
endmodule


module mux_tree_tapbuf_size8_mem_3 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_17__56 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size8_mem_2_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_16__55 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size8_mem_1_2 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_15__54 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size8_mem_0_2 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_14__53 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size8_mem_7 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_13__52 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size8_mem_6 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_12__51 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size8_mem_5 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_11__50 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size8_mem_4 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_10__49 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_40 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size8_3 ( in , sram , sram_inv , out , p0 ) ;
input  [0:7] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;

const1_40 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( in[2] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[4] ) , .A1 ( in[3] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[6] ) , .A1 ( in[5] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
endmodule


module const1_15_9 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size8_2_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:7] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;

const1_15_9 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( in[2] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[4] ) , .A1 ( in[3] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[6] ) , .A1 ( in[5] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
endmodule


module const1_14_9 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size8_1_2 ( in , sram , sram_inv , out , p0 ) ;
input  [0:7] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;

const1_14_9 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( in[2] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[4] ) , .A1 ( in[3] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[6] ) , .A1 ( in[5] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
endmodule


module const1_13_9 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size8_0_2 ( in , sram , sram_inv , out , p0 ) ;
input  [0:7] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;

const1_13_9 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( in[2] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[4] ) , .A1 ( in[3] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[6] ) , .A1 ( in[5] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
endmodule


module const1_12_9 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size8_7 ( in , sram , sram_inv , out , p0 ) ;
input  [0:7] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;

const1_12_9 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( in[2] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[4] ) , .A1 ( in[3] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[6] ) , .A1 ( in[5] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
endmodule


module const1_11_9 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size8_6 ( in , sram , sram_inv , out , p0 ) ;
input  [0:7] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;

const1_11_9 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( in[2] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[4] ) , .A1 ( in[3] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[6] ) , .A1 ( in[5] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
endmodule


module const1_10_9 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size8_5 ( in , sram , sram_inv , out , p0 ) ;
input  [0:7] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;

const1_10_9 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( in[2] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[4] ) , .A1 ( in[3] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[6] ) , .A1 ( in[5] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_2 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[3] ) , .X ( out[0] ) ) ;
endmodule


module const1_9_9 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size8_4 ( in , sram , sram_inv , out , p0 ) ;
input  [0:7] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;

const1_9_9 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( in[2] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[4] ) , .A1 ( in[3] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[6] ) , .A1 ( in[5] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
endmodule


module mux_tree_tapbuf_size10_mem_12 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd1_1 FTB_9__48 ( .A ( mem_out[3] ) , 
    .X ( net_net_69 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 BUFT_RR_69 ( .A ( net_net_69 ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size10_mem_3_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_8__47 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size10_mem_2_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_7__46 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size10_mem_7_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_6__45 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size10_mem_6_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_5__44 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size10_mem_5_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_4__43 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size10_mem_4_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_3__42 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size10_mem_1_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_2__41 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size10_mem_0_2 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_1__40 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_8_9 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size10_12 ( in , sram , sram_inv , out , p0 ) ;
input  [0:9] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

const1_8_9 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[6] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[8] ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[9] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
endmodule


module const1_7_9 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size10_3_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:9] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

const1_7_9 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[6] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[8] ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[9] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
endmodule


module const1_6_10 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size10_2_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:9] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

const1_6_10 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[6] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[8] ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[9] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
endmodule


module const1_5_10 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size10_7_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:9] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

const1_5_10 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[6] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[8] ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[9] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
endmodule


module const1_4_10 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size10_6_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:9] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

const1_4_10 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[6] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[8] ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[9] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
endmodule


module const1_3_10 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size10_5_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:9] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

const1_3_10 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[6] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[8] ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[9] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
endmodule


module const1_2_10 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size10_4_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:9] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

const1_2_10 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[6] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[8] ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[9] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
endmodule


module const1_1_10 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size10_1_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:9] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

const1_1_10 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[6] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[8] ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[9] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
endmodule


module const1_0_10 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size10_0_2 ( in , sram , sram_inv , out , p0 ) ;
input  [0:9] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

const1_0_10 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[6] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[8] ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[9] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
endmodule


module cbx_1__0_ ( prog_clk , chanx_left_in , chanx_right_in , ccff_head , 
    chanx_left_out , chanx_right_out , top_grid_pin_16_ , top_grid_pin_17_ , 
    top_grid_pin_18_ , top_grid_pin_19_ , top_grid_pin_20_ , 
    top_grid_pin_21_ , top_grid_pin_22_ , top_grid_pin_23_ , 
    top_grid_pin_24_ , top_grid_pin_25_ , top_grid_pin_26_ , 
    top_grid_pin_27_ , top_grid_pin_28_ , top_grid_pin_29_ , 
    top_grid_pin_30_ , top_grid_pin_31_ , bottom_grid_pin_0_ , ccff_tail ) ;
input  [0:0] prog_clk ;
input  [0:19] chanx_left_in ;
input  [0:19] chanx_right_in ;
input  [0:0] ccff_head ;
output [0:19] chanx_left_out ;
output [0:19] chanx_right_out ;
output [0:0] top_grid_pin_16_ ;
output [0:0] top_grid_pin_17_ ;
output [0:0] top_grid_pin_18_ ;
output [0:0] top_grid_pin_19_ ;
output [0:0] top_grid_pin_20_ ;
output [0:0] top_grid_pin_21_ ;
output [0:0] top_grid_pin_22_ ;
output [0:0] top_grid_pin_23_ ;
output [0:0] top_grid_pin_24_ ;
output [0:0] top_grid_pin_25_ ;
output [0:0] top_grid_pin_26_ ;
output [0:0] top_grid_pin_27_ ;
output [0:0] top_grid_pin_28_ ;
output [0:0] top_grid_pin_29_ ;
output [0:0] top_grid_pin_30_ ;
output [0:0] top_grid_pin_31_ ;
output [0:0] bottom_grid_pin_0_ ;
output [0:0] ccff_tail ;

wire [0:3] mux_tree_tapbuf_size10_0_sram ;
wire [0:3] mux_tree_tapbuf_size10_0_sram_inv ;
wire [0:3] mux_tree_tapbuf_size10_1_sram ;
wire [0:3] mux_tree_tapbuf_size10_1_sram_inv ;
wire [0:3] mux_tree_tapbuf_size10_2_sram ;
wire [0:3] mux_tree_tapbuf_size10_2_sram_inv ;
wire [0:3] mux_tree_tapbuf_size10_3_sram ;
wire [0:3] mux_tree_tapbuf_size10_3_sram_inv ;
wire [0:3] mux_tree_tapbuf_size10_4_sram ;
wire [0:3] mux_tree_tapbuf_size10_4_sram_inv ;
wire [0:3] mux_tree_tapbuf_size10_5_sram ;
wire [0:3] mux_tree_tapbuf_size10_5_sram_inv ;
wire [0:3] mux_tree_tapbuf_size10_6_sram ;
wire [0:3] mux_tree_tapbuf_size10_6_sram_inv ;
wire [0:3] mux_tree_tapbuf_size10_7_sram ;
wire [0:3] mux_tree_tapbuf_size10_7_sram_inv ;
wire [0:3] mux_tree_tapbuf_size10_8_sram ;
wire [0:3] mux_tree_tapbuf_size10_8_sram_inv ;
wire [0:0] mux_tree_tapbuf_size10_mem_0_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size10_mem_1_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size10_mem_2_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size10_mem_3_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size10_mem_4_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size10_mem_5_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size10_mem_6_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size10_mem_7_ccff_tail ;
wire [0:3] mux_tree_tapbuf_size8_0_sram ;
wire [0:3] mux_tree_tapbuf_size8_0_sram_inv ;
wire [0:3] mux_tree_tapbuf_size8_1_sram ;
wire [0:3] mux_tree_tapbuf_size8_1_sram_inv ;
wire [0:3] mux_tree_tapbuf_size8_2_sram ;
wire [0:3] mux_tree_tapbuf_size8_2_sram_inv ;
wire [0:3] mux_tree_tapbuf_size8_3_sram ;
wire [0:3] mux_tree_tapbuf_size8_3_sram_inv ;
wire [0:3] mux_tree_tapbuf_size8_4_sram ;
wire [0:3] mux_tree_tapbuf_size8_4_sram_inv ;
wire [0:3] mux_tree_tapbuf_size8_5_sram ;
wire [0:3] mux_tree_tapbuf_size8_5_sram_inv ;
wire [0:3] mux_tree_tapbuf_size8_6_sram ;
wire [0:3] mux_tree_tapbuf_size8_6_sram_inv ;
wire [0:3] mux_tree_tapbuf_size8_7_sram ;
wire [0:3] mux_tree_tapbuf_size8_7_sram_inv ;
wire [0:0] mux_tree_tapbuf_size8_mem_0_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size8_mem_1_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size8_mem_2_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size8_mem_3_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size8_mem_4_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size8_mem_5_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size8_mem_6_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size8_mem_7_ccff_tail ;

mux_tree_tapbuf_size10_0_2 mux_bottom_ipin_0 (
    .in ( { chanx_left_in[0] , chanx_right_in[0] , chanx_left_in[2] , 
        chanx_right_in[2] , chanx_left_in[4] , chanx_right_in[4] , 
        chanx_left_in[10] , chanx_right_in[10] , chanx_left_in[16] , 
        chanx_right_in[16] } ) ,
    .sram ( mux_tree_tapbuf_size10_0_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size10_0_sram_inv ) , 
    .out ( top_grid_pin_16_ ) , .p0 ( optlc_net_94 ) ) ;
mux_tree_tapbuf_size10_1_1 mux_bottom_ipin_1 (
    .in ( { chanx_left_in[1] , chanx_right_in[1] , chanx_left_in[3] , 
        chanx_right_in[3] , chanx_left_in[5] , chanx_right_in[5] , 
        chanx_left_in[11] , chanx_right_in[11] , chanx_left_in[17] , 
        chanx_right_in[17] } ) ,
    .sram ( mux_tree_tapbuf_size10_1_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size10_1_sram_inv ) , 
    .out ( top_grid_pin_17_ ) , .p0 ( optlc_net_94 ) ) ;
mux_tree_tapbuf_size10_4_1 mux_bottom_ipin_4 (
    .in ( { chanx_left_in[0] , chanx_right_in[0] , chanx_left_in[2] , 
        chanx_right_in[2] , chanx_left_in[4] , chanx_right_in[4] , 
        chanx_left_in[8] , chanx_right_in[8] , chanx_left_in[14] , 
        chanx_right_in[14] } ) ,
    .sram ( mux_tree_tapbuf_size10_2_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size10_2_sram_inv ) , 
    .out ( top_grid_pin_20_ ) , .p0 ( optlc_net_95 ) ) ;
mux_tree_tapbuf_size10_5_1 mux_bottom_ipin_5 (
    .in ( { chanx_left_in[1] , chanx_right_in[1] , chanx_left_in[3] , 
        chanx_right_in[3] , chanx_left_in[5] , chanx_right_in[5] , 
        chanx_left_in[9] , chanx_right_in[9] , chanx_left_in[15] , 
        chanx_right_in[15] } ) ,
    .sram ( mux_tree_tapbuf_size10_3_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size10_3_sram_inv ) , 
    .out ( top_grid_pin_21_ ) , .p0 ( optlc_net_95 ) ) ;
mux_tree_tapbuf_size10_6_1 mux_bottom_ipin_8 (
    .in ( { chanx_left_in[0] , chanx_right_in[0] , chanx_left_in[2] , 
        chanx_right_in[2] , chanx_left_in[8] , chanx_right_in[8] , 
        chanx_left_in[12] , chanx_right_in[12] , chanx_left_in[18] , 
        chanx_right_in[18] } ) ,
    .sram ( mux_tree_tapbuf_size10_4_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size10_4_sram_inv ) , 
    .out ( top_grid_pin_24_ ) , .p0 ( optlc_net_95 ) ) ;
mux_tree_tapbuf_size10_7_1 mux_bottom_ipin_9 (
    .in ( { chanx_left_in[1] , chanx_right_in[1] , chanx_left_in[3] , 
        chanx_right_in[3] , chanx_left_in[9] , chanx_right_in[9] , 
        chanx_left_in[13] , chanx_right_in[13] , chanx_left_in[19] , 
        chanx_right_in[19] } ) ,
    .sram ( mux_tree_tapbuf_size10_5_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size10_5_sram_inv ) , 
    .out ( top_grid_pin_25_ ) , .p0 ( optlc_net_95 ) ) ;
mux_tree_tapbuf_size10_2_1 mux_bottom_ipin_12 (
    .in ( { chanx_left_in[0] , chanx_right_in[0] , chanx_left_in[2] , 
        chanx_right_in[2] , chanx_left_in[6] , chanx_right_in[6] , 
        chanx_left_in[12] , chanx_right_in[12] , chanx_left_in[16] , 
        chanx_right_in[16] } ) ,
    .sram ( mux_tree_tapbuf_size10_6_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size10_6_sram_inv ) , 
    .out ( top_grid_pin_28_ ) , .p0 ( optlc_net_94 ) ) ;
mux_tree_tapbuf_size10_3_1 mux_bottom_ipin_13 (
    .in ( { chanx_left_in[1] , chanx_right_in[1] , chanx_left_in[3] , 
        chanx_right_in[3] , chanx_left_in[7] , chanx_right_in[7] , 
        chanx_left_in[13] , chanx_right_in[13] , chanx_left_in[17] , 
        chanx_right_in[17] } ) ,
    .sram ( mux_tree_tapbuf_size10_7_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size10_7_sram_inv ) , 
    .out ( top_grid_pin_29_ ) , .p0 ( optlc_net_94 ) ) ;
mux_tree_tapbuf_size10_12 mux_top_ipin_0 (
    .in ( { chanx_left_in[0] , chanx_right_in[0] , chanx_left_in[2] , 
        chanx_right_in[2] , chanx_left_in[4] , chanx_right_in[4] , 
        chanx_left_in[10] , chanx_right_in[10] , chanx_left_in[16] , 
        chanx_right_in[16] } ) ,
    .sram ( mux_tree_tapbuf_size10_8_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size10_8_sram_inv ) , 
    .out ( bottom_grid_pin_0_ ) , .p0 ( optlc_net_95 ) ) ;
mux_tree_tapbuf_size10_mem_0_2 mem_bottom_ipin_0 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( ccff_head ) , 
    .ccff_tail ( mux_tree_tapbuf_size10_mem_0_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size10_0_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size10_0_sram_inv ) ) ;
mux_tree_tapbuf_size10_mem_1_1 mem_bottom_ipin_1 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size10_mem_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size10_mem_1_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size10_1_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size10_1_sram_inv ) ) ;
mux_tree_tapbuf_size10_mem_4_1 mem_bottom_ipin_4 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size8_mem_1_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size10_mem_2_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size10_2_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size10_2_sram_inv ) ) ;
mux_tree_tapbuf_size10_mem_5_1 mem_bottom_ipin_5 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size10_mem_2_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size10_mem_3_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size10_3_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size10_3_sram_inv ) ) ;
mux_tree_tapbuf_size10_mem_6_1 mem_bottom_ipin_8 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size8_mem_3_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size10_mem_4_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size10_4_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size10_4_sram_inv ) ) ;
mux_tree_tapbuf_size10_mem_7_1 mem_bottom_ipin_9 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size10_mem_4_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size10_mem_5_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size10_5_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size10_5_sram_inv ) ) ;
mux_tree_tapbuf_size10_mem_2_1 mem_bottom_ipin_12 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size8_mem_5_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size10_mem_6_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size10_6_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size10_6_sram_inv ) ) ;
mux_tree_tapbuf_size10_mem_3_1 mem_bottom_ipin_13 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size10_mem_6_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size10_mem_7_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size10_7_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size10_7_sram_inv ) ) ;
mux_tree_tapbuf_size10_mem_12 mem_top_ipin_0 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size8_mem_7_ccff_tail ) ,
    .ccff_tail ( { ropt_net_98 } ) ,
    .mem_out ( mux_tree_tapbuf_size10_8_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size10_8_sram_inv ) ) ;
mux_tree_tapbuf_size8_4 mux_bottom_ipin_2 (
    .in ( { chanx_left_in[0] , chanx_right_in[0] , chanx_left_in[2] , 
        chanx_right_in[2] , chanx_left_in[6] , chanx_right_in[6] , 
        chanx_left_in[14] , chanx_right_in[14] } ) ,
    .sram ( mux_tree_tapbuf_size8_0_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size8_0_sram_inv ) , 
    .out ( top_grid_pin_18_ ) , .p0 ( optlc_net_94 ) ) ;
mux_tree_tapbuf_size8_5 mux_bottom_ipin_3 (
    .in ( { chanx_left_in[1] , chanx_right_in[1] , chanx_left_in[3] , 
        chanx_right_in[3] , chanx_left_in[7] , chanx_right_in[7] , 
        chanx_left_in[15] , chanx_right_in[15] } ) ,
    .sram ( mux_tree_tapbuf_size8_1_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size8_1_sram_inv ) , 
    .out ( top_grid_pin_19_ ) , .p0 ( optlc_net_94 ) ) ;
mux_tree_tapbuf_size8_6 mux_bottom_ipin_6 (
    .in ( { chanx_left_in[0] , chanx_right_in[0] , chanx_left_in[2] , 
        chanx_right_in[2] , chanx_left_in[10] , chanx_right_in[10] , 
        chanx_left_in[18] , chanx_right_in[18] } ) ,
    .sram ( mux_tree_tapbuf_size8_2_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size8_2_sram_inv ) , 
    .out ( top_grid_pin_22_ ) , .p0 ( optlc_net_95 ) ) ;
mux_tree_tapbuf_size8_7 mux_bottom_ipin_7 (
    .in ( { chanx_left_in[1] , chanx_right_in[1] , chanx_left_in[3] , 
        chanx_right_in[3] , chanx_left_in[11] , chanx_right_in[11] , 
        chanx_left_in[19] , chanx_right_in[19] } ) ,
    .sram ( mux_tree_tapbuf_size8_3_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size8_3_sram_inv ) , 
    .out ( top_grid_pin_23_ ) , .p0 ( optlc_net_95 ) ) ;
mux_tree_tapbuf_size8_0_2 mux_bottom_ipin_10 (
    .in ( { chanx_left_in[0] , chanx_right_in[0] , chanx_left_in[2] , 
        chanx_right_in[2] , chanx_left_in[6] , chanx_right_in[6] , 
        chanx_left_in[14] , chanx_right_in[14] } ) ,
    .sram ( mux_tree_tapbuf_size8_4_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size8_4_sram_inv ) , 
    .out ( top_grid_pin_26_ ) , .p0 ( optlc_net_95 ) ) ;
mux_tree_tapbuf_size8_1_2 mux_bottom_ipin_11 (
    .in ( { chanx_left_in[1] , chanx_right_in[1] , chanx_left_in[3] , 
        chanx_right_in[3] , chanx_left_in[7] , chanx_right_in[7] , 
        chanx_left_in[15] , chanx_right_in[15] } ) ,
    .sram ( mux_tree_tapbuf_size8_5_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size8_5_sram_inv ) , 
    .out ( top_grid_pin_27_ ) , .p0 ( optlc_net_94 ) ) ;
mux_tree_tapbuf_size8_2_1 mux_bottom_ipin_14 (
    .in ( { chanx_left_in[0] , chanx_right_in[0] , chanx_left_in[2] , 
        chanx_right_in[2] , chanx_left_in[10] , chanx_right_in[10] , 
        chanx_left_in[18] , chanx_right_in[18] } ) ,
    .sram ( mux_tree_tapbuf_size8_6_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size8_6_sram_inv ) , 
    .out ( top_grid_pin_30_ ) , .p0 ( optlc_net_95 ) ) ;
mux_tree_tapbuf_size8_3 mux_bottom_ipin_15 (
    .in ( { chanx_left_in[1] , chanx_right_in[1] , chanx_left_in[3] , 
        chanx_right_in[3] , chanx_left_in[11] , chanx_right_in[11] , 
        chanx_left_in[19] , chanx_right_in[19] } ) ,
    .sram ( mux_tree_tapbuf_size8_7_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size8_7_sram_inv ) , 
    .out ( top_grid_pin_31_ ) , .p0 ( optlc_net_94 ) ) ;
mux_tree_tapbuf_size8_mem_4 mem_bottom_ipin_2 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size10_mem_1_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size8_mem_0_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size8_0_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size8_0_sram_inv ) ) ;
mux_tree_tapbuf_size8_mem_5 mem_bottom_ipin_3 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size8_mem_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size8_mem_1_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size8_1_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size8_1_sram_inv ) ) ;
mux_tree_tapbuf_size8_mem_6 mem_bottom_ipin_6 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size10_mem_3_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size8_mem_2_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size8_2_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size8_2_sram_inv ) ) ;
mux_tree_tapbuf_size8_mem_7 mem_bottom_ipin_7 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size8_mem_2_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size8_mem_3_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size8_3_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size8_3_sram_inv ) ) ;
mux_tree_tapbuf_size8_mem_0_2 mem_bottom_ipin_10 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size10_mem_5_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size8_mem_4_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size8_4_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size8_4_sram_inv ) ) ;
mux_tree_tapbuf_size8_mem_1_2 mem_bottom_ipin_11 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size8_mem_4_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size8_mem_5_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size8_5_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size8_5_sram_inv ) ) ;
mux_tree_tapbuf_size8_mem_2_1 mem_bottom_ipin_14 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size10_mem_7_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size8_mem_6_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size8_6_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size8_6_sram_inv ) ) ;
mux_tree_tapbuf_size8_mem_3 mem_bottom_ipin_15 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size8_mem_6_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size8_mem_7_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size8_7_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size8_7_sram_inv ) ) ;
sky130_fd_sc_hd__conb_1 optlc_89 ( .LO ( SYNOPSYS_UNCONNECTED_1 ) , 
    .HI ( optlc_net_94 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_2__1 ( .A ( chanx_left_in[1] ) , 
    .X ( chanx_right_out[1] ) ) ;
sky130_fd_sc_hd__conb_1 optlc_91 ( .LO ( SYNOPSYS_UNCONNECTED_2 ) , 
    .HI ( optlc_net_95 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_670 ( .A ( chanx_right_in[7] ) , 
    .X ( chanx_left_out[7] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_5__4 ( .A ( chanx_left_in[4] ) , 
    .X ( chanx_right_out[4] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_671 ( .A ( ropt_net_98 ) , 
    .X ( ccff_tail[0] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_7__6 ( .A ( chanx_left_in[6] ) , 
    .X ( chanx_right_out[6] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_673 ( .A ( ropt_net_99 ) , 
    .X ( chanx_left_out[10] ) ) ;
sky130_fd_sc_hd__dlygate4sd1_1 FTB_9__8 ( .A ( chanx_left_in[8] ) , 
    .X ( chanx_right_out[8] ) ) ;
sky130_fd_sc_hd__dlygate4sd1_1 FTB_11__10 ( .A ( chanx_left_in[10] ) , 
    .X ( chanx_right_out[10] ) ) ;
sky130_fd_sc_hd__dlygate4sd1_1 FTB_14__13 ( .A ( chanx_left_in[13] ) , 
    .X ( chanx_right_out[13] ) ) ;
sky130_fd_sc_hd__dlygate4sd1_1 FTB_15__14 ( .A ( chanx_left_in[14] ) , 
    .X ( chanx_right_out[14] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_16__15 ( .A ( chanx_left_in[15] ) , 
    .X ( chanx_right_out[15] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_17__16 ( .A ( chanx_left_in[16] ) , 
    .X ( chanx_right_out[16] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_18__17 ( .A ( chanx_left_in[17] ) , 
    .X ( chanx_right_out[17] ) ) ;
sky130_fd_sc_hd__dlygate4sd1_1 FTB_20__19 ( .A ( chanx_left_in[19] ) , 
    .X ( chanx_right_out[19] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_21__20 ( .A ( chanx_right_in[0] ) , 
    .X ( chanx_left_out[0] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_22__21 ( .A ( chanx_right_in[1] ) , 
    .X ( chanx_left_out[1] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_23__22 ( .A ( chanx_right_in[2] ) , 
    .X ( chanx_left_out[2] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_24__23 ( .A ( chanx_right_in[3] ) , 
    .X ( chanx_left_out[3] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_25__24 ( .A ( chanx_right_in[4] ) , 
    .X ( chanx_left_out[4] ) ) ;
sky130_fd_sc_hd__dlygate4sd1_1 FTB_26__25 ( .A ( chanx_right_in[5] ) , 
    .X ( chanx_left_out[5] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_27__26 ( .A ( chanx_right_in[6] ) , 
    .X ( chanx_left_out[6] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_29__28 ( .A ( chanx_right_in[8] ) , 
    .X ( chanx_left_out[8] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_30__29 ( .A ( chanx_right_in[9] ) , 
    .X ( chanx_left_out[9] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_31__30 ( .A ( chanx_right_in[10] ) , 
    .X ( aps_rename_1_ ) ) ;
sky130_fd_sc_hd__dlygate4sd1_1 FTB_32__31 ( .A ( chanx_right_in[11] ) , 
    .X ( chanx_left_out[11] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_33__32 ( .A ( chanx_right_in[12] ) , 
    .X ( chanx_left_out[12] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_34__33 ( .A ( chanx_right_in[13] ) , 
    .X ( chanx_left_out[13] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_35__34 ( .A ( chanx_right_in[14] ) , 
    .X ( chanx_left_out[14] ) ) ;
sky130_fd_sc_hd__dlygate4sd1_1 FTB_36__35 ( .A ( chanx_right_in[15] ) , 
    .X ( chanx_left_out[15] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_40__39 ( .A ( chanx_right_in[19] ) , 
    .X ( chanx_left_out[19] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_RR_60 ( .A ( chanx_left_in[0] ) , 
    .X ( chanx_right_out[0] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_RR_61 ( .A ( chanx_left_in[5] ) , 
    .X ( chanx_right_out[5] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_RR_62 ( .A ( chanx_left_in[7] ) , 
    .X ( chanx_right_out[7] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_RR_63 ( .A ( chanx_left_in[9] ) , 
    .X ( chanx_right_out[9] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_RR_64 ( .A ( chanx_left_in[11] ) , 
    .X ( chanx_right_out[11] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 BUFT_RR_65 ( .A ( aps_rename_1_ ) , 
    .X ( ropt_net_99 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_RR_67 ( .A ( chanx_right_in[18] ) , 
    .X ( chanx_left_out[18] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_RR_72 ( .A ( chanx_left_in[18] ) , 
    .X ( chanx_right_out[18] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_P_79 ( .A ( chanx_left_in[2] ) , 
    .X ( chanx_right_out[2] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_P_80 ( .A ( chanx_left_in[3] ) , 
    .X ( chanx_right_out[3] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_P_81 ( .A ( chanx_left_in[12] ) , 
    .X ( chanx_right_out[12] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_P_82 ( .A ( chanx_right_in[16] ) , 
    .X ( chanx_left_out[16] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_P_86 ( .A ( chanx_right_in[17] ) , 
    .X ( chanx_left_out[17] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_15_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd1_1 FTB_24__39 ( .A ( mem_out[1] ) , 
    .X ( net_net_75 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_75 ( .A ( net_net_75 ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_22 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_23__38 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_16_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_22__37 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_14_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_21__36 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_13_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_20__35 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_12_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_19__34 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_11_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_18__33 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_10_2 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_17__32 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_9_2 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_16__31 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_8_2 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_15__30 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_7_2 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_14__29 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_6_3 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_13__28 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_5_4 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_12__27 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_4_4 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_11__26 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_3_5 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_10__25 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_2_5 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_9__24 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_1_5 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_8__23 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_0_5 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_7__22 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_39 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_15_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_39 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
endmodule


module const1_22_7 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_22 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_22_7 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
endmodule


module const1_21_7 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_16_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_21_7 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
endmodule


module const1_20_7 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_14_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_20_7 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
endmodule


module const1_19_7 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_13_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_19_7 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
endmodule


module const1_18_7 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_12_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_18_7 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
endmodule


module const1_17_7 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_11_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_17_7 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
endmodule


module const1_16_8 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_10_2 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_16_8 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
endmodule


module const1_15_8 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_9_2 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_15_8 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
endmodule


module const1_14_8 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_8_2 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_14_8 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
endmodule


module const1_13_8 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_7_2 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;

const1_13_8 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_8 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , .X ( out[0] ) ) ;
endmodule


module const1_12_8 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_6_3 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_12_8 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
endmodule


module const1_11_8 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_5_4 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_11_8 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
endmodule


module const1_10_8 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_4_4 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_10_8 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
endmodule


module const1_9_8 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_3_5 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_9_8 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
endmodule


module const1_8_8 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_2_5 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_8_8 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
endmodule


module const1_7_8 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_1_5 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_7_8 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
endmodule


module const1_6_9 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_0_5 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_6_9 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
endmodule


module mux_tree_tapbuf_size3_mem_0_6 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_6__21 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size3_mem_11 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_5__20 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_5_9 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size3_0_6 ( in , sram , sram_inv , out , p0 ) ;
input  [0:2] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;

const1_5_9 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( p0 ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
endmodule


module const1_4_9 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size3_11 ( in , sram , sram_inv , out , p0 ) ;
input  [0:2] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;

const1_4_9 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( p0 ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
endmodule


module mux_tree_tapbuf_size5_mem_8 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_4__19 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size5_mem_0_4 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_3__18 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_3_9 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size5_8 ( in , sram , sram_inv , out , p0 ) ;
input  [0:4] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;

const1_3_9 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , .A1 ( in[4] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
endmodule


module const1_2_9 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size5_0_4 ( in , sram , sram_inv , out , p0 ) ;
input  [0:4] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;

const1_2_9 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , .A1 ( in[4] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
endmodule


module mux_tree_tapbuf_size6_mem_10 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_2__17 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size6_mem_0_6 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_1__16 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_1_9 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size6_10 ( in , sram , sram_inv , out , p0 ) ;
input  [0:5] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;

const1_1_9 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
endmodule


module const1_0_9 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size6_0_6 ( in , sram , sram_inv , out , p0 ) ;
input  [0:5] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;

const1_0_9 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
endmodule


module sb_2__2_ ( prog_clk , chany_bottom_in , bottom_right_grid_pin_1_ , 
    bottom_left_grid_pin_34_ , bottom_left_grid_pin_35_ , 
    bottom_left_grid_pin_36_ , bottom_left_grid_pin_37_ , 
    bottom_left_grid_pin_38_ , bottom_left_grid_pin_39_ , 
    bottom_left_grid_pin_40_ , bottom_left_grid_pin_41_ , chanx_left_in , 
    left_top_grid_pin_1_ , ccff_head , chany_bottom_out , chanx_left_out , 
    ccff_tail ) ;
input  [0:0] prog_clk ;
input  [0:19] chany_bottom_in ;
input  [0:0] bottom_right_grid_pin_1_ ;
input  [0:0] bottom_left_grid_pin_34_ ;
input  [0:0] bottom_left_grid_pin_35_ ;
input  [0:0] bottom_left_grid_pin_36_ ;
input  [0:0] bottom_left_grid_pin_37_ ;
input  [0:0] bottom_left_grid_pin_38_ ;
input  [0:0] bottom_left_grid_pin_39_ ;
input  [0:0] bottom_left_grid_pin_40_ ;
input  [0:0] bottom_left_grid_pin_41_ ;
input  [0:19] chanx_left_in ;
input  [0:0] left_top_grid_pin_1_ ;
input  [0:0] ccff_head ;
output [0:19] chany_bottom_out ;
output [0:19] chanx_left_out ;
output [0:0] ccff_tail ;

wire [0:1] mux_tree_tapbuf_size2_0_sram ;
wire [0:1] mux_tree_tapbuf_size2_0_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_10_sram ;
wire [0:1] mux_tree_tapbuf_size2_10_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_11_sram ;
wire [0:1] mux_tree_tapbuf_size2_11_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_12_sram ;
wire [0:1] mux_tree_tapbuf_size2_12_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_13_sram ;
wire [0:1] mux_tree_tapbuf_size2_13_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_14_sram ;
wire [0:1] mux_tree_tapbuf_size2_14_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_15_sram ;
wire [0:1] mux_tree_tapbuf_size2_15_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_16_sram ;
wire [0:1] mux_tree_tapbuf_size2_16_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_17_sram ;
wire [0:1] mux_tree_tapbuf_size2_17_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_1_sram ;
wire [0:1] mux_tree_tapbuf_size2_1_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_2_sram ;
wire [0:1] mux_tree_tapbuf_size2_2_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_3_sram ;
wire [0:1] mux_tree_tapbuf_size2_3_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_4_sram ;
wire [0:1] mux_tree_tapbuf_size2_4_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_5_sram ;
wire [0:1] mux_tree_tapbuf_size2_5_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_6_sram ;
wire [0:1] mux_tree_tapbuf_size2_6_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_7_sram ;
wire [0:1] mux_tree_tapbuf_size2_7_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_8_sram ;
wire [0:1] mux_tree_tapbuf_size2_8_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_9_sram ;
wire [0:1] mux_tree_tapbuf_size2_9_sram_inv ;
wire [0:0] mux_tree_tapbuf_size2_mem_0_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_10_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_11_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_12_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_13_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_14_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_15_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_16_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_1_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_2_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_3_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_4_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_5_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_6_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_7_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_8_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_9_ccff_tail ;
wire [0:1] mux_tree_tapbuf_size3_0_sram ;
wire [0:1] mux_tree_tapbuf_size3_0_sram_inv ;
wire [0:1] mux_tree_tapbuf_size3_1_sram ;
wire [0:1] mux_tree_tapbuf_size3_1_sram_inv ;
wire [0:0] mux_tree_tapbuf_size3_mem_0_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size3_mem_1_ccff_tail ;
wire [0:2] mux_tree_tapbuf_size5_0_sram ;
wire [0:2] mux_tree_tapbuf_size5_0_sram_inv ;
wire [0:2] mux_tree_tapbuf_size5_1_sram ;
wire [0:2] mux_tree_tapbuf_size5_1_sram_inv ;
wire [0:0] mux_tree_tapbuf_size5_mem_0_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size5_mem_1_ccff_tail ;
wire [0:2] mux_tree_tapbuf_size6_0_sram ;
wire [0:2] mux_tree_tapbuf_size6_0_sram_inv ;
wire [0:2] mux_tree_tapbuf_size6_1_sram ;
wire [0:2] mux_tree_tapbuf_size6_1_sram_inv ;
wire [0:0] mux_tree_tapbuf_size6_mem_0_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size6_mem_1_ccff_tail ;

mux_tree_tapbuf_size6_0_6 mux_bottom_track_1 (
    .in ( { bottom_right_grid_pin_1_[0] , bottom_left_grid_pin_35_[0] , 
        bottom_left_grid_pin_37_[0] , bottom_left_grid_pin_39_[0] , 
        bottom_left_grid_pin_41_[0] , chanx_left_in[1] } ) ,
    .sram ( mux_tree_tapbuf_size6_0_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size6_0_sram_inv ) , 
    .out ( chany_bottom_out[0] ) , .p0 ( optlc_net_96 ) ) ;
mux_tree_tapbuf_size6_10 mux_bottom_track_5 (
    .in ( { bottom_right_grid_pin_1_[0] , bottom_left_grid_pin_35_[0] , 
        bottom_left_grid_pin_37_[0] , bottom_left_grid_pin_39_[0] , 
        bottom_left_grid_pin_41_[0] , chanx_left_in[3] } ) ,
    .sram ( mux_tree_tapbuf_size6_1_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size6_1_sram_inv ) , 
    .out ( chany_bottom_out[2] ) , .p0 ( optlc_net_96 ) ) ;
mux_tree_tapbuf_size6_mem_0_6 mem_bottom_track_1 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( ccff_head ) , 
    .ccff_tail ( mux_tree_tapbuf_size6_mem_0_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size6_0_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size6_0_sram_inv ) ) ;
mux_tree_tapbuf_size6_mem_10 mem_bottom_track_5 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size5_mem_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size6_mem_1_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size6_1_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size6_1_sram_inv ) ) ;
mux_tree_tapbuf_size5_0_4 mux_bottom_track_3 (
    .in ( { bottom_left_grid_pin_34_[0] , bottom_left_grid_pin_36_[0] , 
        bottom_left_grid_pin_38_[0] , bottom_left_grid_pin_40_[0] , 
        chanx_left_in[2] } ) ,
    .sram ( mux_tree_tapbuf_size5_0_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size5_0_sram_inv ) , 
    .out ( chany_bottom_out[1] ) , .p0 ( optlc_net_95 ) ) ;
mux_tree_tapbuf_size5_8 mux_bottom_track_7 (
    .in ( { bottom_left_grid_pin_34_[0] , bottom_left_grid_pin_36_[0] , 
        bottom_left_grid_pin_38_[0] , bottom_left_grid_pin_40_[0] , 
        chanx_left_in[4] } ) ,
    .sram ( mux_tree_tapbuf_size5_1_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size5_1_sram_inv ) , 
    .out ( chany_bottom_out[3] ) , .p0 ( optlc_net_96 ) ) ;
mux_tree_tapbuf_size5_mem_0_4 mem_bottom_track_3 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size6_mem_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size5_mem_0_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size5_0_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size5_0_sram_inv ) ) ;
mux_tree_tapbuf_size5_mem_8 mem_bottom_track_7 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size6_mem_1_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size5_mem_1_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size5_1_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size5_1_sram_inv ) ) ;
mux_tree_tapbuf_size3_11 mux_bottom_track_9 (
    .in ( { bottom_right_grid_pin_1_[0] , bottom_left_grid_pin_41_[0] , 
        chanx_left_in[5] } ) ,
    .sram ( mux_tree_tapbuf_size3_0_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size3_0_sram_inv ) , 
    .out ( chany_bottom_out[4] ) , .p0 ( optlc_net_96 ) ) ;
mux_tree_tapbuf_size3_0_6 mux_bottom_track_25 (
    .in ( { bottom_right_grid_pin_1_[0] , bottom_left_grid_pin_41_[0] , 
        chanx_left_in[13] } ) ,
    .sram ( mux_tree_tapbuf_size3_1_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size3_1_sram_inv ) , 
    .out ( chany_bottom_out[12] ) , .p0 ( optlc_net_97 ) ) ;
mux_tree_tapbuf_size3_mem_11 mem_bottom_track_9 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size5_mem_1_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size3_mem_0_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size3_0_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size3_0_sram_inv ) ) ;
mux_tree_tapbuf_size3_mem_0_6 mem_bottom_track_25 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_6_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size3_mem_1_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size3_1_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size3_1_sram_inv ) ) ;
mux_tree_tapbuf_size2_0_5 mux_bottom_track_11 (
    .in ( { bottom_left_grid_pin_34_[0] , chanx_left_in[6] } ) ,
    .sram ( mux_tree_tapbuf_size2_0_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_0_sram_inv ) , 
    .out ( chany_bottom_out[5] ) , .p0 ( optlc_net_97 ) ) ;
mux_tree_tapbuf_size2_1_5 mux_bottom_track_13 (
    .in ( { bottom_left_grid_pin_35_[0] , chanx_left_in[7] } ) ,
    .sram ( mux_tree_tapbuf_size2_1_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_1_sram_inv ) , 
    .out ( chany_bottom_out[6] ) , .p0 ( optlc_net_97 ) ) ;
mux_tree_tapbuf_size2_2_5 mux_bottom_track_15 (
    .in ( { bottom_left_grid_pin_36_[0] , chanx_left_in[8] } ) ,
    .sram ( mux_tree_tapbuf_size2_2_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_2_sram_inv ) , 
    .out ( chany_bottom_out[7] ) , .p0 ( optlc_net_95 ) ) ;
mux_tree_tapbuf_size2_3_5 mux_bottom_track_17 (
    .in ( { bottom_left_grid_pin_37_[0] , chanx_left_in[9] } ) ,
    .sram ( mux_tree_tapbuf_size2_3_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_3_sram_inv ) , 
    .out ( chany_bottom_out[8] ) , .p0 ( optlc_net_95 ) ) ;
mux_tree_tapbuf_size2_4_4 mux_bottom_track_19 (
    .in ( { bottom_left_grid_pin_38_[0] , chanx_left_in[10] } ) ,
    .sram ( mux_tree_tapbuf_size2_4_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_4_sram_inv ) , 
    .out ( chany_bottom_out[9] ) , .p0 ( optlc_net_95 ) ) ;
mux_tree_tapbuf_size2_5_4 mux_bottom_track_21 (
    .in ( { bottom_left_grid_pin_39_[0] , chanx_left_in[11] } ) ,
    .sram ( mux_tree_tapbuf_size2_5_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_5_sram_inv ) , 
    .out ( chany_bottom_out[10] ) , .p0 ( optlc_net_97 ) ) ;
mux_tree_tapbuf_size2_6_3 mux_bottom_track_23 (
    .in ( { bottom_left_grid_pin_40_[0] , chanx_left_in[12] } ) ,
    .sram ( mux_tree_tapbuf_size2_6_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_6_sram_inv ) , 
    .out ( chany_bottom_out[11] ) , .p0 ( optlc_net_96 ) ) ;
mux_tree_tapbuf_size2_7_2 mux_bottom_track_27 (
    .in ( { bottom_left_grid_pin_34_[0] , chanx_left_in[14] } ) ,
    .sram ( mux_tree_tapbuf_size2_7_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_7_sram_inv ) , 
    .out ( chany_bottom_out[13] ) , .p0 ( optlc_net_97 ) ) ;
mux_tree_tapbuf_size2_8_2 mux_bottom_track_29 (
    .in ( { bottom_left_grid_pin_35_[0] , chanx_left_in[15] } ) ,
    .sram ( mux_tree_tapbuf_size2_8_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_8_sram_inv ) , 
    .out ( chany_bottom_out[14] ) , .p0 ( optlc_net_97 ) ) ;
mux_tree_tapbuf_size2_9_2 mux_bottom_track_31 (
    .in ( { bottom_left_grid_pin_36_[0] , chanx_left_in[16] } ) ,
    .sram ( mux_tree_tapbuf_size2_9_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_9_sram_inv ) , 
    .out ( chany_bottom_out[15] ) , .p0 ( optlc_net_95 ) ) ;
mux_tree_tapbuf_size2_10_2 mux_bottom_track_33 (
    .in ( { bottom_left_grid_pin_37_[0] , chanx_left_in[17] } ) ,
    .sram ( mux_tree_tapbuf_size2_10_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_10_sram_inv ) , 
    .out ( chany_bottom_out[16] ) , .p0 ( optlc_net_95 ) ) ;
mux_tree_tapbuf_size2_11_1 mux_bottom_track_35 (
    .in ( { bottom_left_grid_pin_38_[0] , chanx_left_in[18] } ) ,
    .sram ( mux_tree_tapbuf_size2_11_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_11_sram_inv ) , 
    .out ( chany_bottom_out[17] ) , .p0 ( optlc_net_95 ) ) ;
mux_tree_tapbuf_size2_12_1 mux_bottom_track_37 (
    .in ( { bottom_left_grid_pin_39_[0] , chanx_left_in[19] } ) ,
    .sram ( mux_tree_tapbuf_size2_12_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_12_sram_inv ) , 
    .out ( chany_bottom_out[18] ) , .p0 ( optlc_net_97 ) ) ;
mux_tree_tapbuf_size2_13_1 mux_bottom_track_39 (
    .in ( { bottom_left_grid_pin_40_[0] , chanx_left_in[0] } ) ,
    .sram ( mux_tree_tapbuf_size2_13_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_13_sram_inv ) , 
    .out ( chany_bottom_out[19] ) , .p0 ( optlc_net_96 ) ) ;
mux_tree_tapbuf_size2_14_1 mux_left_track_1 (
    .in ( { chany_bottom_in[19] , left_top_grid_pin_1_[0] } ) ,
    .sram ( mux_tree_tapbuf_size2_14_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_14_sram_inv ) , 
    .out ( chanx_left_out[0] ) , .p0 ( optlc_net_95 ) ) ;
mux_tree_tapbuf_size2_16_1 mux_left_track_5 (
    .in ( { chany_bottom_in[1] , left_top_grid_pin_1_[0] } ) ,
    .sram ( mux_tree_tapbuf_size2_15_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_15_sram_inv ) , 
    .out ( chanx_left_out[2] ) , .p0 ( optlc_net_95 ) ) ;
mux_tree_tapbuf_size2_22 mux_left_track_9 (
    .in ( { chany_bottom_in[3] , left_top_grid_pin_1_[0] } ) ,
    .sram ( mux_tree_tapbuf_size2_16_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_16_sram_inv ) , 
    .out ( chanx_left_out[4] ) , .p0 ( optlc_net_95 ) ) ;
mux_tree_tapbuf_size2_15_1 mux_left_track_25 (
    .in ( { chany_bottom_in[11] , left_top_grid_pin_1_[0] } ) ,
    .sram ( mux_tree_tapbuf_size2_17_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_17_sram_inv ) , 
    .out ( chanx_left_out[12] ) , .p0 ( optlc_net_95 ) ) ;
mux_tree_tapbuf_size2_mem_0_5 mem_bottom_track_11 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size3_mem_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_0_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_0_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_0_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem_1_5 mem_bottom_track_13 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_1_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_1_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_1_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem_2_5 mem_bottom_track_15 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_1_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_2_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_2_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_2_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem_3_5 mem_bottom_track_17 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_2_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_3_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_3_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_3_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem_4_4 mem_bottom_track_19 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_3_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_4_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_4_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_4_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem_5_4 mem_bottom_track_21 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_4_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_5_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_5_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_5_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem_6_3 mem_bottom_track_23 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_5_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_6_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_6_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_6_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem_7_2 mem_bottom_track_27 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size3_mem_1_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_7_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_7_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_7_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem_8_2 mem_bottom_track_29 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_7_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_8_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_8_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_8_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem_9_2 mem_bottom_track_31 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_8_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_9_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_9_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_9_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem_10_2 mem_bottom_track_33 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_9_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_10_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_10_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_10_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem_11_1 mem_bottom_track_35 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_10_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_11_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_11_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_11_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem_12_1 mem_bottom_track_37 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_11_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_12_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_12_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_12_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem_13_1 mem_bottom_track_39 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_12_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_13_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_13_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_13_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem_14_1 mem_left_track_1 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_13_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_14_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_14_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_14_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem_16_1 mem_left_track_5 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_14_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_15_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_15_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_15_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem_22 mem_left_track_9 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_15_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_16_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_16_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_16_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem_15_1 mem_left_track_25 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_16_ccff_tail ) ,
    .ccff_tail ( { ropt_net_102 } ) ,
    .mem_out ( mux_tree_tapbuf_size2_17_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_17_sram_inv ) ) ;
sky130_fd_sc_hd__conb_1 optlc_88 ( .LO ( SYNOPSYS_UNCONNECTED_1 ) , 
    .HI ( optlc_net_95 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_90 ( .LO ( SYNOPSYS_UNCONNECTED_2 ) , 
    .HI ( optlc_net_96 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_92 ( .LO ( SYNOPSYS_UNCONNECTED_3 ) , 
    .HI ( optlc_net_97 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_696 ( .A ( ropt_net_112 ) , 
    .X ( chanx_left_out[3] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_682 ( .A ( chany_bottom_in[2] ) , 
    .X ( ropt_net_112 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_683 ( .A ( ropt_net_99 ) , 
    .X ( ropt_net_117 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_697 ( .A ( ropt_net_113 ) , 
    .X ( chanx_left_out[7] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_698 ( .A ( ropt_net_114 ) , 
    .X ( chanx_left_out[8] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_699 ( .A ( ropt_net_115 ) , 
    .X ( chanx_left_out[9] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_700 ( .A ( ropt_net_116 ) , 
    .X ( chanx_left_out[5] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_701 ( .A ( ropt_net_117 ) , 
    .X ( chanx_left_out[1] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_684 ( .A ( ropt_net_100 ) , 
    .X ( ropt_net_113 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_702 ( .A ( ropt_net_118 ) , 
    .X ( ccff_tail[0] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_685 ( 
    .A ( chany_bottom_in[16] ) , .X ( ropt_net_122 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_703 ( .A ( ropt_net_119 ) , 
    .X ( chanx_left_out[15] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_686 ( .A ( ropt_net_102 ) , 
    .X ( ropt_net_118 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_704 ( .A ( ropt_net_120 ) , 
    .X ( chanx_left_out[19] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_42 ( .A ( chany_bottom_in[4] ) , 
    .X ( ropt_net_110 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_705 ( .A ( ropt_net_121 ) , 
    .X ( chanx_left_out[6] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_706 ( .A ( ropt_net_122 ) , 
    .X ( chanx_left_out[17] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_45 ( .A ( chany_bottom_in[7] ) , 
    .X ( ropt_net_111 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_707 ( .A ( ropt_net_123 ) , 
    .X ( chanx_left_out[13] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_47 ( .A ( chany_bottom_in[9] ) , 
    .X ( BUF_net_47 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_48 ( .A ( chany_bottom_in[10] ) , 
    .X ( BUF_net_48 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_50 ( .A ( chany_bottom_in[13] ) , 
    .X ( BUF_net_50 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_687 ( .A ( ropt_net_103 ) , 
    .X ( ropt_net_115 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_688 ( 
    .A ( chany_bottom_in[12] ) , .X ( ropt_net_123 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_689 ( 
    .A ( chany_bottom_in[15] ) , .X ( chanx_left_out[16] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 BUFT_RR_60 ( .A ( BUF_net_47 ) , 
    .X ( chanx_left_out[10] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 BUFT_RR_61 ( .A ( BUF_net_48 ) , 
    .X ( chanx_left_out[11] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_690 ( 
    .A ( chany_bottom_in[17] ) , .X ( chanx_left_out[18] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_691 ( .A ( chany_bottom_in[5] ) , 
    .X ( ropt_net_121 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_692 ( 
    .A ( chany_bottom_in[18] ) , .X ( ropt_net_120 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_P_76 ( .A ( chany_bottom_in[8] ) , 
    .X ( ropt_net_103 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 BUFT_P_78 ( .A ( BUF_net_50 ) , 
    .X ( chanx_left_out[14] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_P_81 ( .A ( chany_bottom_in[0] ) , 
    .X ( ropt_net_99 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_P_82 ( .A ( chany_bottom_in[6] ) , 
    .X ( ropt_net_100 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_693 ( 
    .A ( chany_bottom_in[14] ) , .X ( ropt_net_119 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_694 ( .A ( ropt_net_110 ) , 
    .X ( ropt_net_116 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_695 ( .A ( ropt_net_111 ) , 
    .X ( ropt_net_114 ) ) ;
endmodule


module mux_tree_tapbuf_size3_mem_10 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_27__59 ( .A ( mem_out[1] ) , 
    .X ( net_net_75 ) ) ;
sky130_fd_sc_hd__dlygate4sd1_1 BUFT_RR_75 ( .A ( net_net_75 ) , 
    .X ( net_net_74 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_90 ( .A ( net_net_74 ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size3_mem_3_3 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_26__58 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size3_mem_2_4 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_25__57 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size3_mem_1_4 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_24__56 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size3_mem_0_5 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_23__55 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_38 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size3_10 ( in , sram , sram_inv , out , p0 ) ;
input  [0:2] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;

const1_38 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( p0 ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
endmodule


module const1_25_6 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size3_3_3 ( in , sram , sram_inv , out , p0 ) ;
input  [0:2] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;

const1_25_6 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( p0 ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
endmodule


module const1_24_6 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size3_2_4 ( in , sram , sram_inv , out , p0 ) ;
input  [0:2] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;

const1_24_6 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( p0 ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
endmodule


module const1_23_6 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size3_1_4 ( in , sram , sram_inv , out , p0 ) ;
input  [0:2] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;

const1_23_6 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( p0 ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
endmodule


module const1_22_6 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size3_0_5 ( in , sram , sram_inv , out , p0 ) ;
input  [0:2] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;

const1_22_6 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( p0 ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
endmodule


module mux_tree_tapbuf_size4_mem_2_2 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_22__54 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size4_mem_1_2 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_21__53 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size4_mem_0_3 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_20__52 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size4_mem_8 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_19__51 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_21_6 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size4_2_2 ( in , sram , sram_inv , out , p0 ) ;
input  [0:3] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;

const1_21_6 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( in[2] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , .A1 ( in[3] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
endmodule


module const1_20_6 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size4_1_2 ( in , sram , sram_inv , out , p0 ) ;
input  [0:3] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;

const1_20_6 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( in[2] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , .A1 ( in[3] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
endmodule


module const1_19_6 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size4_0_3 ( in , sram , sram_inv , out , p0 ) ;
input  [0:3] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;

const1_19_6 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( in[2] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , .A1 ( in[3] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
endmodule


module const1_18_6 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size4_8 ( in , sram , sram_inv , out , p0 ) ;
input  [0:3] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;

const1_18_6 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( in[2] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , .A1 ( in[3] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
endmodule


module mux_tree_tapbuf_size9_mem_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_18__50 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_17_6 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size9_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:8] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;

const1_17_6 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[7] ) , .A1 ( in[6] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[8] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
endmodule


module mux_tree_tapbuf_size6_mem_1_3 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_17__49 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size6_mem_0_5 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_16__48 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size6_mem_9 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_15__47 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_16_7 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size6_1_3 ( in , sram , sram_inv , out , p0 ) ;
input  [0:5] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;

const1_16_7 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
endmodule


module const1_15_7 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size6_0_5 ( in , sram , sram_inv , out , p0 ) ;
input  [0:5] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;

const1_15_7 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
endmodule


module const1_14_7 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size6_9 ( in , sram , sram_inv , out , p0 ) ;
input  [0:5] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;

const1_14_7 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
endmodule


module mux_tree_tapbuf_size7_mem_4_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_14__46 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size7_mem_3_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_13__45 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size7_mem_2_3 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_12__44 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size7_mem_1_4 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_11__43 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size7_mem_0_4 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_10__42 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size7_mem_8 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_9__41 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size7_mem_5_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_8__40 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_13_7 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size7_4_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:6] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;

const1_13_7 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_3_ ( .A0 ( p0 ) , .A1 ( in[6] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
endmodule


module const1_12_7 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size7_3_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:6] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;

const1_12_7 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_3_ ( .A0 ( p0 ) , .A1 ( in[6] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
endmodule


module const1_11_7 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size7_2_3 ( in , sram , sram_inv , out , p0 ) ;
input  [0:6] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;

const1_11_7 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_3_ ( .A0 ( p0 ) , .A1 ( in[6] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_61 ( 
    .A ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , .X ( out[0] ) ) ;
endmodule


module const1_10_7 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size7_1_4 ( in , sram , sram_inv , out , p0 ) ;
input  [0:6] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;

const1_10_7 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_3_ ( .A0 ( p0 ) , .A1 ( in[6] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
endmodule


module const1_9_7 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size7_0_4 ( in , sram , sram_inv , out , p0 ) ;
input  [0:6] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;

const1_9_7 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_3_ ( .A0 ( p0 ) , .A1 ( in[6] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
endmodule


module const1_8_7 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size7_8 ( in , sram , sram_inv , out , p0 ) ;
input  [0:6] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;

const1_8_7 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_3_ ( .A0 ( p0 ) , .A1 ( in[6] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
endmodule


module const1_7_7 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size7_5_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:6] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;

const1_7_7 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_3_ ( .A0 ( p0 ) , .A1 ( in[6] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
endmodule


module mux_tree_tapbuf_size14_mem_0_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_7__39 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size14_mem_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_6__38 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_6_8 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size14_0_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:13] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_10_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_11_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_12_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_13_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

const1_6_8 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_13_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_3_ ( .A0 ( in[7] ) , .A1 ( in[6] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_4_ ( .A0 ( in[9] ) , .A1 ( in[8] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_5_ ( .A0 ( in[11] ) , .A1 ( in[10] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_6_ ( .A0 ( in[13] ) , .A1 ( in[12] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_10_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_11_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_10_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_12_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_12_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_11_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_13_X[0] ) ) ;
endmodule


module const1_5_8 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size14_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:13] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_10_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_11_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_12_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_13_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

const1_5_8 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_13_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_3_ ( .A0 ( in[7] ) , .A1 ( in[6] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_4_ ( .A0 ( in[9] ) , .A1 ( in[8] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_5_ ( .A0 ( in[11] ) , .A1 ( in[10] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_6_ ( .A0 ( in[13] ) , .A1 ( in[12] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_10_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_11_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_10_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_12_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_12_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_11_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_13_X[0] ) ) ;
endmodule


module mux_tree_tapbuf_size8_mem_0_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_5__37 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size8_mem_3 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_4__36 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size8_mem_1_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_3__35 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_4_8 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size8_0_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:7] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;

const1_4_8 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( in[2] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[4] ) , .A1 ( in[3] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[6] ) , .A1 ( in[5] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
endmodule


module const1_3_8 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size8_3 ( in , sram , sram_inv , out , p0 ) ;
input  [0:7] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;

const1_3_8 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( in[2] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[4] ) , .A1 ( in[3] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[6] ) , .A1 ( in[5] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
endmodule


module const1_2_8 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size8_1_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:7] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;

const1_2_8 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( in[2] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[4] ) , .A1 ( in[3] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[6] ) , .A1 ( in[5] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
endmodule


module mux_tree_tapbuf_size10_mem_0_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_2__34 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size10_mem_11 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_1__33 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_1_8 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size10_0_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:9] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

const1_1_8 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[6] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[8] ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[9] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
endmodule


module const1_0_8 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size10_11 ( in , sram , sram_inv , out , p0 ) ;
input  [0:9] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

const1_0_8 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[6] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[8] ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[9] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
endmodule


module sb_2__1_ ( prog_clk , chany_top_in , top_left_grid_pin_34_ , 
    top_left_grid_pin_35_ , top_left_grid_pin_36_ , top_left_grid_pin_37_ , 
    top_left_grid_pin_38_ , top_left_grid_pin_39_ , top_left_grid_pin_40_ , 
    top_left_grid_pin_41_ , top_right_grid_pin_1_ , chany_bottom_in , 
    bottom_right_grid_pin_1_ , bottom_left_grid_pin_34_ , 
    bottom_left_grid_pin_35_ , bottom_left_grid_pin_36_ , 
    bottom_left_grid_pin_37_ , bottom_left_grid_pin_38_ , 
    bottom_left_grid_pin_39_ , bottom_left_grid_pin_40_ , 
    bottom_left_grid_pin_41_ , chanx_left_in , left_top_grid_pin_42_ , 
    left_top_grid_pin_43_ , left_top_grid_pin_44_ , left_top_grid_pin_45_ , 
    left_top_grid_pin_46_ , left_top_grid_pin_47_ , left_top_grid_pin_48_ , 
    left_top_grid_pin_49_ , ccff_head , chany_top_out , chany_bottom_out , 
    chanx_left_out , ccff_tail ) ;
input  [0:0] prog_clk ;
input  [0:19] chany_top_in ;
input  [0:0] top_left_grid_pin_34_ ;
input  [0:0] top_left_grid_pin_35_ ;
input  [0:0] top_left_grid_pin_36_ ;
input  [0:0] top_left_grid_pin_37_ ;
input  [0:0] top_left_grid_pin_38_ ;
input  [0:0] top_left_grid_pin_39_ ;
input  [0:0] top_left_grid_pin_40_ ;
input  [0:0] top_left_grid_pin_41_ ;
input  [0:0] top_right_grid_pin_1_ ;
input  [0:19] chany_bottom_in ;
input  [0:0] bottom_right_grid_pin_1_ ;
input  [0:0] bottom_left_grid_pin_34_ ;
input  [0:0] bottom_left_grid_pin_35_ ;
input  [0:0] bottom_left_grid_pin_36_ ;
input  [0:0] bottom_left_grid_pin_37_ ;
input  [0:0] bottom_left_grid_pin_38_ ;
input  [0:0] bottom_left_grid_pin_39_ ;
input  [0:0] bottom_left_grid_pin_40_ ;
input  [0:0] bottom_left_grid_pin_41_ ;
input  [0:19] chanx_left_in ;
input  [0:0] left_top_grid_pin_42_ ;
input  [0:0] left_top_grid_pin_43_ ;
input  [0:0] left_top_grid_pin_44_ ;
input  [0:0] left_top_grid_pin_45_ ;
input  [0:0] left_top_grid_pin_46_ ;
input  [0:0] left_top_grid_pin_47_ ;
input  [0:0] left_top_grid_pin_48_ ;
input  [0:0] left_top_grid_pin_49_ ;
input  [0:0] ccff_head ;
output [0:19] chany_top_out ;
output [0:19] chany_bottom_out ;
output [0:19] chanx_left_out ;
output [0:0] ccff_tail ;

wire [0:3] mux_tree_tapbuf_size10_0_sram ;
wire [0:3] mux_tree_tapbuf_size10_0_sram_inv ;
wire [0:3] mux_tree_tapbuf_size10_1_sram ;
wire [0:3] mux_tree_tapbuf_size10_1_sram_inv ;
wire [0:0] mux_tree_tapbuf_size10_mem_0_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size10_mem_1_ccff_tail ;
wire [0:3] mux_tree_tapbuf_size14_0_sram ;
wire [0:3] mux_tree_tapbuf_size14_0_sram_inv ;
wire [0:3] mux_tree_tapbuf_size14_1_sram ;
wire [0:3] mux_tree_tapbuf_size14_1_sram_inv ;
wire [0:0] mux_tree_tapbuf_size14_mem_0_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size14_mem_1_ccff_tail ;
wire [0:1] mux_tree_tapbuf_size3_0_sram ;
wire [0:1] mux_tree_tapbuf_size3_0_sram_inv ;
wire [0:1] mux_tree_tapbuf_size3_1_sram ;
wire [0:1] mux_tree_tapbuf_size3_1_sram_inv ;
wire [0:1] mux_tree_tapbuf_size3_2_sram ;
wire [0:1] mux_tree_tapbuf_size3_2_sram_inv ;
wire [0:1] mux_tree_tapbuf_size3_3_sram ;
wire [0:1] mux_tree_tapbuf_size3_3_sram_inv ;
wire [0:1] mux_tree_tapbuf_size3_4_sram ;
wire [0:1] mux_tree_tapbuf_size3_4_sram_inv ;
wire [0:0] mux_tree_tapbuf_size3_mem_0_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size3_mem_1_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size3_mem_2_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size3_mem_3_ccff_tail ;
wire [0:2] mux_tree_tapbuf_size4_0_sram ;
wire [0:2] mux_tree_tapbuf_size4_0_sram_inv ;
wire [0:2] mux_tree_tapbuf_size4_1_sram ;
wire [0:2] mux_tree_tapbuf_size4_1_sram_inv ;
wire [0:2] mux_tree_tapbuf_size4_2_sram ;
wire [0:2] mux_tree_tapbuf_size4_2_sram_inv ;
wire [0:2] mux_tree_tapbuf_size4_3_sram ;
wire [0:2] mux_tree_tapbuf_size4_3_sram_inv ;
wire [0:0] mux_tree_tapbuf_size4_mem_0_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size4_mem_1_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size4_mem_2_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size4_mem_3_ccff_tail ;
wire [0:2] mux_tree_tapbuf_size6_0_sram ;
wire [0:2] mux_tree_tapbuf_size6_0_sram_inv ;
wire [0:2] mux_tree_tapbuf_size6_1_sram ;
wire [0:2] mux_tree_tapbuf_size6_1_sram_inv ;
wire [0:2] mux_tree_tapbuf_size6_2_sram ;
wire [0:2] mux_tree_tapbuf_size6_2_sram_inv ;
wire [0:0] mux_tree_tapbuf_size6_mem_0_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size6_mem_1_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size6_mem_2_ccff_tail ;
wire [0:2] mux_tree_tapbuf_size7_0_sram ;
wire [0:2] mux_tree_tapbuf_size7_0_sram_inv ;
wire [0:2] mux_tree_tapbuf_size7_1_sram ;
wire [0:2] mux_tree_tapbuf_size7_1_sram_inv ;
wire [0:2] mux_tree_tapbuf_size7_2_sram ;
wire [0:2] mux_tree_tapbuf_size7_2_sram_inv ;
wire [0:2] mux_tree_tapbuf_size7_3_sram ;
wire [0:2] mux_tree_tapbuf_size7_3_sram_inv ;
wire [0:2] mux_tree_tapbuf_size7_4_sram ;
wire [0:2] mux_tree_tapbuf_size7_4_sram_inv ;
wire [0:2] mux_tree_tapbuf_size7_5_sram ;
wire [0:2] mux_tree_tapbuf_size7_5_sram_inv ;
wire [0:2] mux_tree_tapbuf_size7_6_sram ;
wire [0:2] mux_tree_tapbuf_size7_6_sram_inv ;
wire [0:0] mux_tree_tapbuf_size7_mem_0_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size7_mem_1_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size7_mem_2_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size7_mem_3_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size7_mem_4_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size7_mem_5_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size7_mem_6_ccff_tail ;
wire [0:3] mux_tree_tapbuf_size8_0_sram ;
wire [0:3] mux_tree_tapbuf_size8_0_sram_inv ;
wire [0:3] mux_tree_tapbuf_size8_1_sram ;
wire [0:3] mux_tree_tapbuf_size8_1_sram_inv ;
wire [0:3] mux_tree_tapbuf_size8_2_sram ;
wire [0:3] mux_tree_tapbuf_size8_2_sram_inv ;
wire [0:0] mux_tree_tapbuf_size8_mem_0_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size8_mem_1_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size8_mem_2_ccff_tail ;
wire [0:3] mux_tree_tapbuf_size9_0_sram ;
wire [0:3] mux_tree_tapbuf_size9_0_sram_inv ;
wire [0:0] mux_tree_tapbuf_size9_mem_0_ccff_tail ;

mux_tree_tapbuf_size10_11 mux_top_track_0 (
    .in ( { top_left_grid_pin_34_[0] , top_left_grid_pin_36_[0] , 
        top_left_grid_pin_38_[0] , top_left_grid_pin_40_[0] , 
        top_right_grid_pin_1_[0] , chany_bottom_in[2] , chany_bottom_in[12] , 
        chanx_left_in[0] , chanx_left_in[7] , chanx_left_in[14] } ) ,
    .sram ( mux_tree_tapbuf_size10_0_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size10_0_sram_inv ) , 
    .out ( chany_top_out[0] ) , .p0 ( optlc_net_104 ) ) ;
mux_tree_tapbuf_size10_0_1 mux_bottom_track_1 (
    .in ( { chany_top_in[2] , chany_top_in[12] , bottom_right_grid_pin_1_[0] , 
        bottom_left_grid_pin_35_[0] , bottom_left_grid_pin_37_[0] , 
        bottom_left_grid_pin_39_[0] , bottom_left_grid_pin_41_[0] , 
        chanx_left_in[1] , chanx_left_in[8] , chanx_left_in[15] } ) ,
    .sram ( mux_tree_tapbuf_size10_1_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size10_1_sram_inv ) , 
    .out ( chany_bottom_out[0] ) , .p0 ( optlc_net_105 ) ) ;
mux_tree_tapbuf_size10_mem_11 mem_top_track_0 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( ccff_head ) , 
    .ccff_tail ( mux_tree_tapbuf_size10_mem_0_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size10_0_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size10_0_sram_inv ) ) ;
mux_tree_tapbuf_size10_mem_0_1 mem_bottom_track_1 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size6_mem_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size10_mem_1_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size10_1_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size10_1_sram_inv ) ) ;
mux_tree_tapbuf_size8_1_1 mux_top_track_2 (
    .in ( { top_left_grid_pin_35_[0] , top_left_grid_pin_37_[0] , 
        top_left_grid_pin_39_[0] , top_left_grid_pin_41_[0] , 
        chany_bottom_in[4] , chany_bottom_in[13] , chanx_left_in[6] , 
        chanx_left_in[13] } ) ,
    .sram ( mux_tree_tapbuf_size8_0_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size8_0_sram_inv ) , 
    .out ( chany_top_out[1] ) , .p0 ( optlc_net_104 ) ) ;
mux_tree_tapbuf_size8_3 mux_top_track_8 (
    .in ( { top_left_grid_pin_34_[0] , top_left_grid_pin_38_[0] , 
        top_right_grid_pin_1_[0] , chany_bottom_in[6] , chany_bottom_in[16] , 
        chanx_left_in[4] , chanx_left_in[11] , chanx_left_in[18] } ) ,
    .sram ( mux_tree_tapbuf_size8_1_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size8_1_sram_inv ) , 
    .out ( chany_top_out[4] ) , .p0 ( optlc_net_106 ) ) ;
mux_tree_tapbuf_size8_0_1 mux_bottom_track_9 (
    .in ( { chany_top_in[6] , chany_top_in[16] , bottom_right_grid_pin_1_[0] , 
        bottom_left_grid_pin_37_[0] , bottom_left_grid_pin_41_[0] , 
        chanx_left_in[4] , chanx_left_in[11] , chanx_left_in[18] } ) ,
    .sram ( mux_tree_tapbuf_size8_2_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size8_2_sram_inv ) , 
    .out ( chany_bottom_out[4] ) , .p0 ( optlc_net_103 ) ) ;
mux_tree_tapbuf_size8_mem_1_1 mem_top_track_2 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size10_mem_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size8_mem_0_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size8_0_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size8_0_sram_inv ) ) ;
mux_tree_tapbuf_size8_mem_3 mem_top_track_8 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size14_mem_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size8_mem_1_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size8_1_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size8_1_sram_inv ) ) ;
mux_tree_tapbuf_size8_mem_0_1 mem_bottom_track_9 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size14_mem_1_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size8_mem_2_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size8_2_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size8_2_sram_inv ) ) ;
mux_tree_tapbuf_size14_1 mux_top_track_4 (
    .in ( { top_left_grid_pin_34_[0] , top_left_grid_pin_35_[0] , 
        top_left_grid_pin_36_[0] , top_left_grid_pin_37_[0] , 
        top_left_grid_pin_38_[0] , top_left_grid_pin_39_[0] , 
        top_left_grid_pin_40_[0] , top_left_grid_pin_41_[0] , 
        top_right_grid_pin_1_[0] , chany_bottom_in[5] , chany_bottom_in[14] , 
        chanx_left_in[5] , chanx_left_in[12] , chanx_left_in[19] } ) ,
    .sram ( mux_tree_tapbuf_size14_0_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size14_0_sram_inv ) , 
    .out ( chany_top_out[2] ) , .p0 ( optlc_net_104 ) ) ;
mux_tree_tapbuf_size14_0_1 mux_bottom_track_5 (
    .in ( { chany_top_in[5] , chany_top_in[14] , bottom_right_grid_pin_1_[0] , 
        bottom_left_grid_pin_34_[0] , bottom_left_grid_pin_35_[0] , 
        bottom_left_grid_pin_36_[0] , bottom_left_grid_pin_37_[0] , 
        bottom_left_grid_pin_38_[0] , bottom_left_grid_pin_39_[0] , 
        bottom_left_grid_pin_40_[0] , bottom_left_grid_pin_41_[0] , 
        chanx_left_in[3] , chanx_left_in[10] , chanx_left_in[17] } ) ,
    .sram ( mux_tree_tapbuf_size14_1_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size14_1_sram_inv ) , 
    .out ( chany_bottom_out[2] ) , .p0 ( optlc_net_103 ) ) ;
mux_tree_tapbuf_size14_mem_1 mem_top_track_4 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size8_mem_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size14_mem_0_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size14_0_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size14_0_sram_inv ) ) ;
mux_tree_tapbuf_size14_mem_0_1 mem_bottom_track_5 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size9_mem_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size14_mem_1_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size14_1_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size14_1_sram_inv ) ) ;
mux_tree_tapbuf_size7_5_1 mux_top_track_16 (
    .in ( { top_left_grid_pin_35_[0] , top_left_grid_pin_39_[0] , 
        chany_bottom_in[8] , chany_bottom_in[17] , chanx_left_in[3] , 
        chanx_left_in[10] , chanx_left_in[17] } ) ,
    .sram ( mux_tree_tapbuf_size7_0_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size7_0_sram_inv ) , 
    .out ( chany_top_out[8] ) , .p0 ( optlc_net_104 ) ) ;
mux_tree_tapbuf_size7_8 mux_top_track_24 (
    .in ( { top_left_grid_pin_36_[0] , top_left_grid_pin_40_[0] , 
        chany_bottom_in[9] , chany_bottom_in[18] , chanx_left_in[2] , 
        chanx_left_in[9] , chanx_left_in[16] } ) ,
    .sram ( mux_tree_tapbuf_size7_1_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size7_1_sram_inv ) , 
    .out ( chany_top_out[12] ) , .p0 ( optlc_net_105 ) ) ;
mux_tree_tapbuf_size7_0_4 mux_bottom_track_17 (
    .in ( { chany_top_in[8] , chany_top_in[17] , bottom_left_grid_pin_34_[0] , 
        bottom_left_grid_pin_38_[0] , chanx_left_in[5] , chanx_left_in[12] , 
        chanx_left_in[19] } ) ,
    .sram ( mux_tree_tapbuf_size7_2_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size7_2_sram_inv ) , 
    .out ( chany_bottom_out[8] ) , .p0 ( optlc_net_103 ) ) ;
mux_tree_tapbuf_size7_1_4 mux_left_track_1 (
    .in ( { chany_top_in[0] , chany_top_in[2] , chany_bottom_in[2] , 
        left_top_grid_pin_42_[0] , left_top_grid_pin_44_[0] , 
        left_top_grid_pin_46_[0] , left_top_grid_pin_48_[0] } ) ,
    .sram ( mux_tree_tapbuf_size7_3_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size7_3_sram_inv ) , 
    .out ( chanx_left_out[0] ) , .p0 ( optlc_net_104 ) ) ;
mux_tree_tapbuf_size7_2_3 mux_left_track_3 (
    .in ( { chany_top_in[4] , chany_bottom_in[0] , chany_bottom_in[4] , 
        left_top_grid_pin_43_[0] , left_top_grid_pin_45_[0] , 
        left_top_grid_pin_47_[0] , left_top_grid_pin_49_[0] } ) ,
    .sram ( mux_tree_tapbuf_size7_4_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size7_4_sram_inv ) ,
    .out ( { ropt_net_108 } ) ,
    .p0 ( optlc_net_104 ) ) ;
mux_tree_tapbuf_size7_3_1 mux_left_track_5 (
    .in ( { chany_top_in[5] , chany_bottom_in[1] , chany_bottom_in[5] , 
        left_top_grid_pin_42_[0] , left_top_grid_pin_44_[0] , 
        left_top_grid_pin_46_[0] , left_top_grid_pin_48_[0] } ) ,
    .sram ( mux_tree_tapbuf_size7_5_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size7_5_sram_inv ) , 
    .out ( chanx_left_out[2] ) , .p0 ( optlc_net_104 ) ) ;
mux_tree_tapbuf_size7_4_1 mux_left_track_7 (
    .in ( { chany_top_in[6] , chany_bottom_in[3] , chany_bottom_in[6] , 
        left_top_grid_pin_43_[0] , left_top_grid_pin_45_[0] , 
        left_top_grid_pin_47_[0] , left_top_grid_pin_49_[0] } ) ,
    .sram ( mux_tree_tapbuf_size7_6_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size7_6_sram_inv ) , 
    .out ( chanx_left_out[3] ) , .p0 ( optlc_net_106 ) ) ;
mux_tree_tapbuf_size7_mem_5_1 mem_top_track_16 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size8_mem_1_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size7_mem_0_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size7_0_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size7_0_sram_inv ) ) ;
mux_tree_tapbuf_size7_mem_8 mem_top_track_24 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size7_mem_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size7_mem_1_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size7_1_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size7_1_sram_inv ) ) ;
mux_tree_tapbuf_size7_mem_0_4 mem_bottom_track_17 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size8_mem_2_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size7_mem_2_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size7_2_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size7_2_sram_inv ) ) ;
mux_tree_tapbuf_size7_mem_1_4 mem_left_track_1 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size6_mem_2_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size7_mem_3_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size7_3_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size7_3_sram_inv ) ) ;
mux_tree_tapbuf_size7_mem_2_3 mem_left_track_3 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size7_mem_3_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size7_mem_4_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size7_4_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size7_4_sram_inv ) ) ;
mux_tree_tapbuf_size7_mem_3_1 mem_left_track_5 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size7_mem_4_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size7_mem_5_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size7_5_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size7_5_sram_inv ) ) ;
mux_tree_tapbuf_size7_mem_4_1 mem_left_track_7 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size7_mem_5_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size7_mem_6_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size7_6_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size7_6_sram_inv ) ) ;
mux_tree_tapbuf_size6_9 mux_top_track_32 (
    .in ( { top_left_grid_pin_37_[0] , top_left_grid_pin_41_[0] , 
        chany_bottom_in[10] , chanx_left_in[1] , chanx_left_in[8] , 
        chanx_left_in[15] } ) ,
    .sram ( mux_tree_tapbuf_size6_0_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size6_0_sram_inv ) , 
    .out ( chany_top_out[16] ) , .p0 ( optlc_net_105 ) ) ;
mux_tree_tapbuf_size6_0_5 mux_bottom_track_25 (
    .in ( { chany_top_in[9] , chany_top_in[18] , bottom_left_grid_pin_35_[0] , 
        bottom_left_grid_pin_39_[0] , chanx_left_in[6] , chanx_left_in[13] } ) ,
    .sram ( mux_tree_tapbuf_size6_1_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size6_1_sram_inv ) , 
    .out ( chany_bottom_out[12] ) , .p0 ( optlc_net_103 ) ) ;
mux_tree_tapbuf_size6_1_3 mux_bottom_track_33 (
    .in ( { chany_top_in[10] , bottom_left_grid_pin_36_[0] , 
        bottom_left_grid_pin_40_[0] , chanx_left_in[0] , chanx_left_in[7] , 
        chanx_left_in[14] } ) ,
    .sram ( mux_tree_tapbuf_size6_2_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size6_2_sram_inv ) , 
    .out ( chany_bottom_out[16] ) , .p0 ( optlc_net_105 ) ) ;
mux_tree_tapbuf_size6_mem_9 mem_top_track_32 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size7_mem_1_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size6_mem_0_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size6_0_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size6_0_sram_inv ) ) ;
mux_tree_tapbuf_size6_mem_0_5 mem_bottom_track_25 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size7_mem_2_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size6_mem_1_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size6_1_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size6_1_sram_inv ) ) ;
mux_tree_tapbuf_size6_mem_1_3 mem_bottom_track_33 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size6_mem_1_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size6_mem_2_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size6_2_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size6_2_sram_inv ) ) ;
mux_tree_tapbuf_size9_1 mux_bottom_track_3 (
    .in ( { chany_top_in[4] , chany_top_in[13] , bottom_left_grid_pin_34_[0] , 
        bottom_left_grid_pin_36_[0] , bottom_left_grid_pin_38_[0] , 
        bottom_left_grid_pin_40_[0] , chanx_left_in[2] , chanx_left_in[9] , 
        chanx_left_in[16] } ) ,
    .sram ( mux_tree_tapbuf_size9_0_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size9_0_sram_inv ) , 
    .out ( chany_bottom_out[1] ) , .p0 ( optlc_net_105 ) ) ;
mux_tree_tapbuf_size9_mem_1 mem_bottom_track_3 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size10_mem_1_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size9_mem_0_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size9_0_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size9_0_sram_inv ) ) ;
mux_tree_tapbuf_size4_8 mux_left_track_9 (
    .in ( { chany_top_in[8] , chany_bottom_in[7] , chany_bottom_in[8] , 
        left_top_grid_pin_42_[0] } ) ,
    .sram ( mux_tree_tapbuf_size4_0_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size4_0_sram_inv ) , 
    .out ( chanx_left_out[4] ) , .p0 ( optlc_net_103 ) ) ;
mux_tree_tapbuf_size4_0_3 mux_left_track_11 (
    .in ( { chany_top_in[9] , chany_bottom_in[9] , chany_bottom_in[11] , 
        left_top_grid_pin_43_[0] } ) ,
    .sram ( mux_tree_tapbuf_size4_1_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size4_1_sram_inv ) , 
    .out ( chanx_left_out[5] ) , .p0 ( optlc_net_103 ) ) ;
mux_tree_tapbuf_size4_1_2 mux_left_track_13 (
    .in ( { chany_top_in[10] , chany_bottom_in[10] , chany_bottom_in[15] , 
        left_top_grid_pin_44_[0] } ) ,
    .sram ( mux_tree_tapbuf_size4_2_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size4_2_sram_inv ) , 
    .out ( chanx_left_out[6] ) , .p0 ( optlc_net_103 ) ) ;
mux_tree_tapbuf_size4_2_2 mux_left_track_15 (
    .in ( { chany_top_in[12] , chany_bottom_in[12] , chany_bottom_in[19] , 
        left_top_grid_pin_45_[0] } ) ,
    .sram ( mux_tree_tapbuf_size4_3_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size4_3_sram_inv ) , 
    .out ( chanx_left_out[7] ) , .p0 ( optlc_net_103 ) ) ;
mux_tree_tapbuf_size4_mem_8 mem_left_track_9 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size7_mem_6_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size4_mem_0_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size4_0_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size4_0_sram_inv ) ) ;
mux_tree_tapbuf_size4_mem_0_3 mem_left_track_11 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size4_mem_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size4_mem_1_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size4_1_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size4_1_sram_inv ) ) ;
mux_tree_tapbuf_size4_mem_1_2 mem_left_track_13 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size4_mem_1_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size4_mem_2_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size4_2_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size4_2_sram_inv ) ) ;
mux_tree_tapbuf_size4_mem_2_2 mem_left_track_15 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size4_mem_2_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size4_mem_3_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size4_3_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size4_3_sram_inv ) ) ;
mux_tree_tapbuf_size3_0_5 mux_left_track_17 (
    .in ( { chany_top_in[13] , chany_bottom_in[13] , 
        left_top_grid_pin_46_[0] } ) ,
    .sram ( mux_tree_tapbuf_size3_0_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size3_0_sram_inv ) , 
    .out ( chanx_left_out[8] ) , .p0 ( optlc_net_104 ) ) ;
mux_tree_tapbuf_size3_1_4 mux_left_track_19 (
    .in ( { chany_top_in[14] , chany_bottom_in[14] , 
        left_top_grid_pin_47_[0] } ) ,
    .sram ( mux_tree_tapbuf_size3_1_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size3_1_sram_inv ) , 
    .out ( chanx_left_out[9] ) , .p0 ( optlc_net_106 ) ) ;
mux_tree_tapbuf_size3_2_4 mux_left_track_21 (
    .in ( { chany_top_in[16] , chany_bottom_in[16] , 
        left_top_grid_pin_48_[0] } ) ,
    .sram ( mux_tree_tapbuf_size3_2_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size3_2_sram_inv ) , 
    .out ( chanx_left_out[10] ) , .p0 ( optlc_net_106 ) ) ;
mux_tree_tapbuf_size3_3_3 mux_left_track_23 (
    .in ( { chany_top_in[17] , chany_bottom_in[17] , 
        left_top_grid_pin_49_[0] } ) ,
    .sram ( mux_tree_tapbuf_size3_3_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size3_3_sram_inv ) , 
    .out ( chanx_left_out[11] ) , .p0 ( optlc_net_106 ) ) ;
mux_tree_tapbuf_size3_10 mux_left_track_25 (
    .in ( { chany_top_in[18] , chany_bottom_in[18] , 
        left_top_grid_pin_42_[0] } ) ,
    .sram ( mux_tree_tapbuf_size3_4_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size3_4_sram_inv ) , 
    .out ( chanx_left_out[12] ) , .p0 ( optlc_net_104 ) ) ;
mux_tree_tapbuf_size3_mem_0_5 mem_left_track_17 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size4_mem_3_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size3_mem_0_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size3_0_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size3_0_sram_inv ) ) ;
mux_tree_tapbuf_size3_mem_1_4 mem_left_track_19 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size3_mem_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size3_mem_1_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size3_1_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size3_1_sram_inv ) ) ;
mux_tree_tapbuf_size3_mem_2_4 mem_left_track_21 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size3_mem_1_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size3_mem_2_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size3_2_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size3_2_sram_inv ) ) ;
mux_tree_tapbuf_size3_mem_3_3 mem_left_track_23 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size3_mem_2_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size3_mem_3_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size3_3_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size3_3_sram_inv ) ) ;
mux_tree_tapbuf_size3_mem_10 mem_left_track_25 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size3_mem_3_ccff_tail ) ,
    .ccff_tail ( { ropt_net_115 } ) ,
    .mem_out ( mux_tree_tapbuf_size3_4_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size3_4_sram_inv ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_1__0 ( .A ( chany_top_in[1] ) , 
    .X ( ropt_net_117 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_2__1 ( .A ( chany_top_in[2] ) , 
    .X ( ropt_net_125 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_97 ( .LO ( SYNOPSYS_UNCONNECTED_1 ) , 
    .HI ( optlc_net_103 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_4__3 ( .A ( chany_top_in[4] ) , 
    .X ( ropt_net_122 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_5__4 ( .A ( chany_top_in[5] ) , 
    .X ( ropt_net_116 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_99 ( .LO ( SYNOPSYS_UNCONNECTED_2 ) , 
    .HI ( optlc_net_104 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_7__6 ( .A ( chany_top_in[7] ) , 
    .X ( ropt_net_135 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_8__7 ( .A ( chany_top_in[8] ) , 
    .X ( ropt_net_123 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_9__8 ( .A ( chany_top_in[9] ) , 
    .X ( ropt_net_128 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_10__9 ( .A ( chany_top_in[10] ) , 
    .X ( chany_bottom_out[11] ) ) ;
sky130_fd_sc_hd__conb_1 optlc_101 ( .LO ( SYNOPSYS_UNCONNECTED_3 ) , 
    .HI ( optlc_net_105 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_12__11 ( .A ( chany_top_in[12] ) , 
    .X ( chany_bottom_out[13] ) ) ;
sky130_fd_sc_hd__conb_1 optlc_103 ( .LO ( SYNOPSYS_UNCONNECTED_4 ) , 
    .HI ( optlc_net_106 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_14__13 ( .A ( chany_top_in[14] ) , 
    .X ( ropt_net_127 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_741 ( .A ( ropt_net_137 ) , 
    .X ( chanx_left_out[1] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_16__15 ( .A ( chany_top_in[16] ) , 
    .X ( ropt_net_131 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_17__16 ( .A ( chany_top_in[17] ) , 
    .X ( ropt_net_133 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_18__17 ( .A ( chany_top_in[18] ) , 
    .X ( ropt_net_134 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_705 ( .A ( chany_top_in[11] ) , 
    .X ( ropt_net_140 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_20__19 ( .A ( chany_bottom_in[2] ) , 
    .X ( chany_top_out[3] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_706 ( .A ( ropt_net_108 ) , 
    .X ( ropt_net_137 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_22__21 ( .A ( chany_bottom_in[5] ) , 
    .X ( chany_top_out[6] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_707 ( .A ( chany_top_in[19] ) , 
    .X ( chanx_left_out[14] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_24__23 ( .A ( chany_bottom_in[8] ) , 
    .X ( chany_top_out[9] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_708 ( 
    .A ( left_top_grid_pin_43_[0] ) , .X ( chanx_left_out[13] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_709 ( .A ( chany_top_in[6] ) , 
    .X ( chany_bottom_out[7] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_27__26 ( .A ( chany_bottom_in[12] ) , 
    .X ( ropt_net_120 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_710 ( 
    .A ( chany_bottom_in[17] ) , .X ( chany_top_out[18] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_711 ( .A ( chany_top_in[15] ) , 
    .X ( chanx_left_out[15] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_30__29 ( .A ( chany_bottom_in[16] ) , 
    .X ( ropt_net_132 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_712 ( .A ( chany_top_in[3] ) , 
    .X ( ropt_net_148 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_714 ( .A ( ropt_net_115 ) , 
    .X ( ropt_net_141 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_715 ( .A ( ropt_net_116 ) , 
    .X ( chany_bottom_out[6] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_716 ( .A ( ropt_net_117 ) , 
    .X ( ropt_net_144 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_742 ( .A ( ropt_net_138 ) , 
    .X ( chanx_left_out[17] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_717 ( .A ( ropt_net_118 ) , 
    .X ( chany_top_out[5] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_RR_67 ( .A ( chany_bottom_in[4] ) , 
    .X ( ropt_net_118 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_RR_68 ( .A ( chany_bottom_in[6] ) , 
    .X ( ropt_net_129 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_RR_69 ( .A ( chany_bottom_in[9] ) , 
    .X ( ropt_net_119 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_RR_70 ( .A ( chany_bottom_in[10] ) , 
    .X ( ropt_net_121 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_71 ( .A ( chany_bottom_in[13] ) , 
    .X ( ropt_net_124 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_743 ( .A ( ropt_net_139 ) , 
    .X ( chany_top_out[14] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_RR_73 ( .A ( chany_bottom_in[18] ) , 
    .X ( chany_top_out[19] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_718 ( .A ( ropt_net_119 ) , 
    .X ( chany_top_out[10] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_719 ( .A ( ropt_net_120 ) , 
    .X ( ropt_net_146 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_720 ( .A ( ropt_net_121 ) , 
    .X ( chany_top_out[11] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_744 ( .A ( ropt_net_140 ) , 
    .X ( chanx_left_out[16] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_P_86 ( .A ( chany_top_in[13] ) , 
    .X ( ropt_net_126 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_P_87 ( .A ( chany_bottom_in[14] ) , 
    .X ( ropt_net_130 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_746 ( .A ( ropt_net_141 ) , 
    .X ( ccff_tail[0] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_747 ( .A ( ropt_net_142 ) , 
    .X ( chany_bottom_out[19] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_721 ( .A ( ropt_net_122 ) , 
    .X ( chany_bottom_out[5] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_748 ( .A ( ropt_net_143 ) , 
    .X ( chany_top_out[15] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_722 ( .A ( ropt_net_123 ) , 
    .X ( chany_bottom_out[9] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_723 ( .A ( ropt_net_124 ) , 
    .X ( ropt_net_139 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_724 ( .A ( ropt_net_125 ) , 
    .X ( chany_bottom_out[3] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_725 ( .A ( ropt_net_126 ) , 
    .X ( chany_bottom_out[14] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_726 ( .A ( ropt_net_127 ) , 
    .X ( chany_bottom_out[15] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_727 ( .A ( ropt_net_128 ) , 
    .X ( chany_bottom_out[10] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_728 ( .A ( ropt_net_129 ) , 
    .X ( chany_top_out[7] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_729 ( .A ( ropt_net_130 ) , 
    .X ( ropt_net_143 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_731 ( .A ( ropt_net_131 ) , 
    .X ( chany_bottom_out[17] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_732 ( .A ( ropt_net_132 ) , 
    .X ( ropt_net_145 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_733 ( .A ( ropt_net_133 ) , 
    .X ( ropt_net_147 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_737 ( .A ( ropt_net_134 ) , 
    .X ( ropt_net_142 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_740 ( .A ( ropt_net_135 ) , 
    .X ( ropt_net_138 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_749 ( .A ( ropt_net_144 ) , 
    .X ( chanx_left_out[19] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_751 ( .A ( ropt_net_145 ) , 
    .X ( chany_top_out[17] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_756 ( .A ( ropt_net_146 ) , 
    .X ( chany_top_out[13] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_759 ( .A ( ropt_net_147 ) , 
    .X ( chany_bottom_out[18] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_764 ( .A ( ropt_net_148 ) , 
    .X ( chanx_left_out[18] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_7_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_34__39 ( .A ( mem_out[1] ) , 
    .X ( net_net_62 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_87 ( .A ( net_net_62 ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_6_2 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_33__38 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_5_3 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_32__37 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_4_3 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_31__36 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_3_4 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_30__35 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_2_4 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_29__34 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_1_4 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_28__33 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_0_4 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_27__32 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_21 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_26__31 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_20 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_25__30 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_19 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_24__29 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_18 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_23__28 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_17 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_22__27 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_16 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_21__26 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_15 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_20__25 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_14 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_19__24 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_13 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_18__23 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_12 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_17__22 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_11 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_16__21 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_10_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_15__20 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_9_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_14__19 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_8_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_13__18 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_37 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_7_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_37 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
endmodule


module const1_32_1 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_6_2 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_32_1 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
endmodule


module const1_31_2 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_5_3 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_31_2 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
endmodule


module const1_30_3 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_4_3 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_30_3 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
endmodule


module const1_29_3 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_3_4 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_29_3 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_59 ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
endmodule


module const1_28_3 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_2_4 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_28_3 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
endmodule


module const1_27_3 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_1_4 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_27_3 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
endmodule


module const1_26_5 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_0_4 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_26_5 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
endmodule


module const1_25_5 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_21 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_25_5 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
endmodule


module const1_24_5 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_20 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_24_5 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
endmodule


module const1_23_5 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_19 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_23_5 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
endmodule


module const1_22_5 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_18 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_22_5 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_57 ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
endmodule


module const1_21_5 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_17 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;

const1_21_5 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_8 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , .X ( out[0] ) ) ;
endmodule


module const1_20_5 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_16 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_20_5 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_55 ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( BUF_net_55 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_P_93 ( .A ( BUF_net_55 ) , 
    .X ( out[0] ) ) ;
endmodule


module const1_19_5 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_15 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_19_5 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
endmodule


module const1_18_5 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_14 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_18_5 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_53 ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
endmodule


module const1_17_5 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_13 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;

const1_17_5 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_8 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , .X ( out[0] ) ) ;
endmodule


module const1_16_6 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_12 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_16_6 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
endmodule


module const1_15_6 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_11 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_15_6 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
endmodule


module const1_14_6 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_10_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_14_6 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
endmodule


module const1_13_6 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_9_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_13_6 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
endmodule


module const1_12_6 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_8_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_12_6 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
endmodule


module mux_tree_tapbuf_size3_mem_0_4 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_12__17 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size3_mem_1_3 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_11__16 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size3_mem_2_3 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_10__15 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size3_mem_9 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_9__14 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_11_6 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size3_0_4 ( in , sram , sram_inv , out , p0 ) ;
input  [0:2] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;

const1_11_6 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( p0 ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
endmodule


module const1_10_6 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size3_1_3 ( in , sram , sram_inv , out , p0 ) ;
input  [0:2] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;

const1_10_6 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( p0 ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
endmodule


module const1_9_6 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size3_2_3 ( in , sram , sram_inv , out , p0 ) ;
input  [0:2] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;

const1_9_6 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( p0 ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_46 ( 
    .A ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .X ( out[0] ) ) ;
endmodule


module const1_8_6 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size3_9 ( in , sram , sram_inv , out , p0 ) ;
input  [0:2] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;

const1_8_6 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( p0 ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_P_90 ( 
    .A ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .X ( out[0] ) ) ;
endmodule


module mux_tree_tapbuf_size5_mem_1_2 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_8__13 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size5_mem_0_3 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_7__12 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size5_mem_7 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_6__11 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size5_mem_2_2 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_5__10 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_7_6 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size5_1_2 ( in , sram , sram_inv , out , p0 ) ;
input  [0:4] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;

const1_7_6 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , .A1 ( in[4] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
endmodule


module const1_6_7 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size5_0_3 ( in , sram , sram_inv , out , p0 ) ;
input  [0:4] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;

const1_6_7 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , .A1 ( in[4] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
endmodule


module const1_5_7 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size5_7 ( in , sram , sram_inv , out , p0 ) ;
input  [0:4] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;

const1_5_7 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , .A1 ( in[4] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
endmodule


module const1_4_7 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size5_2_2 ( in , sram , sram_inv , out , p0 ) ;
input  [0:4] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;

const1_4_7 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , .A1 ( in[4] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
endmodule


module mux_tree_tapbuf_size6_mem_1_2 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_4__9 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size6_mem_0_4 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_3__8 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size6_mem_8 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_2__7 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size6_mem_2_2 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_1__6 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_3_7 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size6_1_2 ( in , sram , sram_inv , out , p0 ) ;
input  [0:5] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;

const1_3_7 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_42 ( 
    .A ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .X ( out[0] ) ) ;
endmodule


module const1_2_7 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size6_0_4 ( in , sram , sram_inv , out , p0 ) ;
input  [0:5] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;

const1_2_7 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
endmodule


module const1_1_7 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size6_8 ( in , sram , sram_inv , out , p0 ) ;
input  [0:5] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;

const1_1_7 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
endmodule


module const1_0_7 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size6_2_2 ( in , sram , sram_inv , out , p0 ) ;
input  [0:5] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;

const1_0_7 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_8 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , .X ( out[0] ) ) ;
endmodule


module sb_2__0_ ( prog_clk , chany_top_in , top_left_grid_pin_34_ , 
    top_left_grid_pin_35_ , top_left_grid_pin_36_ , top_left_grid_pin_37_ , 
    top_left_grid_pin_38_ , top_left_grid_pin_39_ , top_left_grid_pin_40_ , 
    top_left_grid_pin_41_ , top_right_grid_pin_1_ , chanx_left_in , 
    left_top_grid_pin_42_ , left_top_grid_pin_43_ , left_top_grid_pin_44_ , 
    left_top_grid_pin_45_ , left_top_grid_pin_46_ , left_top_grid_pin_47_ , 
    left_top_grid_pin_48_ , left_top_grid_pin_49_ , left_bottom_grid_pin_1_ , 
    ccff_head , chany_top_out , chanx_left_out , ccff_tail ) ;
input  [0:0] prog_clk ;
input  [0:19] chany_top_in ;
input  [0:0] top_left_grid_pin_34_ ;
input  [0:0] top_left_grid_pin_35_ ;
input  [0:0] top_left_grid_pin_36_ ;
input  [0:0] top_left_grid_pin_37_ ;
input  [0:0] top_left_grid_pin_38_ ;
input  [0:0] top_left_grid_pin_39_ ;
input  [0:0] top_left_grid_pin_40_ ;
input  [0:0] top_left_grid_pin_41_ ;
input  [0:0] top_right_grid_pin_1_ ;
input  [0:19] chanx_left_in ;
input  [0:0] left_top_grid_pin_42_ ;
input  [0:0] left_top_grid_pin_43_ ;
input  [0:0] left_top_grid_pin_44_ ;
input  [0:0] left_top_grid_pin_45_ ;
input  [0:0] left_top_grid_pin_46_ ;
input  [0:0] left_top_grid_pin_47_ ;
input  [0:0] left_top_grid_pin_48_ ;
input  [0:0] left_top_grid_pin_49_ ;
input  [0:0] left_bottom_grid_pin_1_ ;
input  [0:0] ccff_head ;
output [0:19] chany_top_out ;
output [0:19] chanx_left_out ;
output [0:0] ccff_tail ;

wire [0:1] mux_tree_tapbuf_size2_0_sram ;
wire [0:1] mux_tree_tapbuf_size2_0_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_10_sram ;
wire [0:1] mux_tree_tapbuf_size2_10_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_11_sram ;
wire [0:1] mux_tree_tapbuf_size2_11_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_12_sram ;
wire [0:1] mux_tree_tapbuf_size2_12_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_13_sram ;
wire [0:1] mux_tree_tapbuf_size2_13_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_14_sram ;
wire [0:1] mux_tree_tapbuf_size2_14_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_15_sram ;
wire [0:1] mux_tree_tapbuf_size2_15_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_16_sram ;
wire [0:1] mux_tree_tapbuf_size2_16_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_17_sram ;
wire [0:1] mux_tree_tapbuf_size2_17_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_18_sram ;
wire [0:1] mux_tree_tapbuf_size2_18_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_19_sram ;
wire [0:1] mux_tree_tapbuf_size2_19_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_1_sram ;
wire [0:1] mux_tree_tapbuf_size2_1_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_20_sram ;
wire [0:1] mux_tree_tapbuf_size2_20_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_21_sram ;
wire [0:1] mux_tree_tapbuf_size2_21_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_2_sram ;
wire [0:1] mux_tree_tapbuf_size2_2_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_3_sram ;
wire [0:1] mux_tree_tapbuf_size2_3_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_4_sram ;
wire [0:1] mux_tree_tapbuf_size2_4_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_5_sram ;
wire [0:1] mux_tree_tapbuf_size2_5_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_6_sram ;
wire [0:1] mux_tree_tapbuf_size2_6_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_7_sram ;
wire [0:1] mux_tree_tapbuf_size2_7_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_8_sram ;
wire [0:1] mux_tree_tapbuf_size2_8_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_9_sram ;
wire [0:1] mux_tree_tapbuf_size2_9_sram_inv ;
wire [0:0] mux_tree_tapbuf_size2_mem_0_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_10_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_11_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_12_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_13_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_14_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_15_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_16_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_17_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_18_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_19_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_1_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_20_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_2_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_3_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_4_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_5_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_6_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_7_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_8_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_9_ccff_tail ;
wire [0:1] mux_tree_tapbuf_size3_0_sram ;
wire [0:1] mux_tree_tapbuf_size3_0_sram_inv ;
wire [0:1] mux_tree_tapbuf_size3_1_sram ;
wire [0:1] mux_tree_tapbuf_size3_1_sram_inv ;
wire [0:1] mux_tree_tapbuf_size3_2_sram ;
wire [0:1] mux_tree_tapbuf_size3_2_sram_inv ;
wire [0:1] mux_tree_tapbuf_size3_3_sram ;
wire [0:1] mux_tree_tapbuf_size3_3_sram_inv ;
wire [0:0] mux_tree_tapbuf_size3_mem_0_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size3_mem_1_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size3_mem_2_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size3_mem_3_ccff_tail ;
wire [0:2] mux_tree_tapbuf_size5_0_sram ;
wire [0:2] mux_tree_tapbuf_size5_0_sram_inv ;
wire [0:2] mux_tree_tapbuf_size5_1_sram ;
wire [0:2] mux_tree_tapbuf_size5_1_sram_inv ;
wire [0:2] mux_tree_tapbuf_size5_2_sram ;
wire [0:2] mux_tree_tapbuf_size5_2_sram_inv ;
wire [0:2] mux_tree_tapbuf_size5_3_sram ;
wire [0:2] mux_tree_tapbuf_size5_3_sram_inv ;
wire [0:0] mux_tree_tapbuf_size5_mem_0_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size5_mem_1_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size5_mem_2_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size5_mem_3_ccff_tail ;
wire [0:2] mux_tree_tapbuf_size6_0_sram ;
wire [0:2] mux_tree_tapbuf_size6_0_sram_inv ;
wire [0:2] mux_tree_tapbuf_size6_1_sram ;
wire [0:2] mux_tree_tapbuf_size6_1_sram_inv ;
wire [0:2] mux_tree_tapbuf_size6_2_sram ;
wire [0:2] mux_tree_tapbuf_size6_2_sram_inv ;
wire [0:2] mux_tree_tapbuf_size6_3_sram ;
wire [0:2] mux_tree_tapbuf_size6_3_sram_inv ;
wire [0:0] mux_tree_tapbuf_size6_mem_0_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size6_mem_1_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size6_mem_2_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size6_mem_3_ccff_tail ;

mux_tree_tapbuf_size6_2_2 mux_top_track_0 (
    .in ( { top_left_grid_pin_34_[0] , top_left_grid_pin_36_[0] , 
        top_left_grid_pin_38_[0] , top_left_grid_pin_40_[0] , 
        top_right_grid_pin_1_[0] , chanx_left_in[0] } ) ,
    .sram ( mux_tree_tapbuf_size6_0_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size6_0_sram_inv ) , 
    .out ( chany_top_out[0] ) , .p0 ( optlc_net_111 ) ) ;
mux_tree_tapbuf_size6_8 mux_top_track_4 (
    .in ( { top_left_grid_pin_34_[0] , top_left_grid_pin_36_[0] , 
        top_left_grid_pin_38_[0] , top_left_grid_pin_40_[0] , 
        top_right_grid_pin_1_[0] , chanx_left_in[18] } ) ,
    .sram ( mux_tree_tapbuf_size6_1_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size6_1_sram_inv ) , 
    .out ( chany_top_out[2] ) , .p0 ( optlc_net_111 ) ) ;
mux_tree_tapbuf_size6_0_4 mux_left_track_1 (
    .in ( { chany_top_in[0] , left_top_grid_pin_42_[0] , 
        left_top_grid_pin_44_[0] , left_top_grid_pin_46_[0] , 
        left_top_grid_pin_48_[0] , left_bottom_grid_pin_1_[0] } ) ,
    .sram ( mux_tree_tapbuf_size6_2_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size6_2_sram_inv ) , 
    .out ( chanx_left_out[0] ) , .p0 ( optlc_net_113 ) ) ;
mux_tree_tapbuf_size6_1_2 mux_left_track_5 (
    .in ( { chany_top_in[18] , left_top_grid_pin_42_[0] , 
        left_top_grid_pin_44_[0] , left_top_grid_pin_46_[0] , 
        left_top_grid_pin_48_[0] , left_bottom_grid_pin_1_[0] } ) ,
    .sram ( mux_tree_tapbuf_size6_3_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size6_3_sram_inv ) ,
    .out ( { ropt_net_120 } ) ,
    .p0 ( optlc_net_113 ) ) ;
mux_tree_tapbuf_size6_mem_2_2 mem_top_track_0 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( ccff_head ) , 
    .ccff_tail ( mux_tree_tapbuf_size6_mem_0_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size6_0_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size6_0_sram_inv ) ) ;
mux_tree_tapbuf_size6_mem_8 mem_top_track_4 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size5_mem_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size6_mem_1_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size6_1_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size6_1_sram_inv ) ) ;
mux_tree_tapbuf_size6_mem_0_4 mem_left_track_1 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_13_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size6_mem_2_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size6_2_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size6_2_sram_inv ) ) ;
mux_tree_tapbuf_size6_mem_1_2 mem_left_track_5 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size5_mem_2_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size6_mem_3_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size6_3_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size6_3_sram_inv ) ) ;
mux_tree_tapbuf_size5_2_2 mux_top_track_2 (
    .in ( { top_left_grid_pin_35_[0] , top_left_grid_pin_37_[0] , 
        top_left_grid_pin_39_[0] , top_left_grid_pin_41_[0] , 
        chanx_left_in[19] } ) ,
    .sram ( mux_tree_tapbuf_size5_0_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size5_0_sram_inv ) , 
    .out ( chany_top_out[1] ) , .p0 ( optlc_net_111 ) ) ;
mux_tree_tapbuf_size5_7 mux_top_track_6 (
    .in ( { top_left_grid_pin_35_[0] , top_left_grid_pin_37_[0] , 
        top_left_grid_pin_39_[0] , top_left_grid_pin_41_[0] , 
        chanx_left_in[17] } ) ,
    .sram ( mux_tree_tapbuf_size5_1_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size5_1_sram_inv ) , 
    .out ( chany_top_out[3] ) , .p0 ( optlc_net_111 ) ) ;
mux_tree_tapbuf_size5_0_3 mux_left_track_3 (
    .in ( { chany_top_in[19] , left_top_grid_pin_43_[0] , 
        left_top_grid_pin_45_[0] , left_top_grid_pin_47_[0] , 
        left_top_grid_pin_49_[0] } ) ,
    .sram ( mux_tree_tapbuf_size5_2_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size5_2_sram_inv ) , 
    .out ( chanx_left_out[1] ) , .p0 ( optlc_net_113 ) ) ;
mux_tree_tapbuf_size5_1_2 mux_left_track_7 (
    .in ( { chany_top_in[17] , left_top_grid_pin_43_[0] , 
        left_top_grid_pin_45_[0] , left_top_grid_pin_47_[0] , 
        left_top_grid_pin_49_[0] } ) ,
    .sram ( mux_tree_tapbuf_size5_3_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size5_3_sram_inv ) , 
    .out ( chanx_left_out[3] ) , .p0 ( optlc_net_112 ) ) ;
mux_tree_tapbuf_size5_mem_2_2 mem_top_track_2 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size6_mem_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size5_mem_0_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size5_0_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size5_0_sram_inv ) ) ;
mux_tree_tapbuf_size5_mem_7 mem_top_track_6 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size6_mem_1_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size5_mem_1_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size5_1_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size5_1_sram_inv ) ) ;
mux_tree_tapbuf_size5_mem_0_3 mem_left_track_3 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size6_mem_2_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size5_mem_2_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size5_2_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size5_2_sram_inv ) ) ;
mux_tree_tapbuf_size5_mem_1_2 mem_left_track_7 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size6_mem_3_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size5_mem_3_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size5_3_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size5_3_sram_inv ) ) ;
mux_tree_tapbuf_size3_9 mux_top_track_8 (
    .in ( { top_left_grid_pin_34_[0] , top_right_grid_pin_1_[0] , 
        chanx_left_in[16] } ) ,
    .sram ( mux_tree_tapbuf_size3_0_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size3_0_sram_inv ) ,
    .out ( { ropt_net_122 } ) ,
    .p0 ( optlc_net_111 ) ) ;
mux_tree_tapbuf_size3_2_3 mux_top_track_24 (
    .in ( { top_left_grid_pin_34_[0] , top_right_grid_pin_1_[0] , 
        chanx_left_in[8] } ) ,
    .sram ( mux_tree_tapbuf_size3_1_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size3_1_sram_inv ) ,
    .out ( { ropt_net_123 } ) ,
    .p0 ( optlc_net_111 ) ) ;
mux_tree_tapbuf_size3_1_3 mux_left_track_9 (
    .in ( { chany_top_in[16] , left_top_grid_pin_42_[0] , 
        left_bottom_grid_pin_1_[0] } ) ,
    .sram ( mux_tree_tapbuf_size3_2_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size3_2_sram_inv ) , 
    .out ( chanx_left_out[4] ) , .p0 ( optlc_net_110 ) ) ;
mux_tree_tapbuf_size3_0_4 mux_left_track_25 (
    .in ( { chany_top_in[8] , left_top_grid_pin_42_[0] , 
        left_bottom_grid_pin_1_[0] } ) ,
    .sram ( mux_tree_tapbuf_size3_3_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size3_3_sram_inv ) , 
    .out ( chanx_left_out[12] ) , .p0 ( optlc_net_113 ) ) ;
mux_tree_tapbuf_size3_mem_9 mem_top_track_8 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size5_mem_1_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size3_mem_0_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size3_0_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size3_0_sram_inv ) ) ;
mux_tree_tapbuf_size3_mem_2_3 mem_top_track_24 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_6_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size3_mem_1_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size3_1_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size3_1_sram_inv ) ) ;
mux_tree_tapbuf_size3_mem_1_3 mem_left_track_9 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size5_mem_3_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size3_mem_2_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size3_2_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size3_2_sram_inv ) ) ;
mux_tree_tapbuf_size3_mem_0_4 mem_left_track_25 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_20_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size3_mem_3_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size3_3_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size3_3_sram_inv ) ) ;
mux_tree_tapbuf_size2_8_1 mux_top_track_10 (
    .in ( { top_left_grid_pin_35_[0] , chanx_left_in[15] } ) ,
    .sram ( mux_tree_tapbuf_size2_0_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_0_sram_inv ) , 
    .out ( chany_top_out[5] ) , .p0 ( optlc_net_111 ) ) ;
mux_tree_tapbuf_size2_9_1 mux_top_track_12 (
    .in ( { top_left_grid_pin_36_[0] , chanx_left_in[14] } ) ,
    .sram ( mux_tree_tapbuf_size2_1_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_1_sram_inv ) , 
    .out ( chany_top_out[6] ) , .p0 ( optlc_net_110 ) ) ;
mux_tree_tapbuf_size2_10_1 mux_top_track_14 (
    .in ( { top_left_grid_pin_37_[0] , chanx_left_in[13] } ) ,
    .sram ( mux_tree_tapbuf_size2_2_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_2_sram_inv ) , 
    .out ( chany_top_out[7] ) , .p0 ( optlc_net_110 ) ) ;
mux_tree_tapbuf_size2_11 mux_top_track_16 (
    .in ( { top_left_grid_pin_38_[0] , chanx_left_in[12] } ) ,
    .sram ( mux_tree_tapbuf_size2_3_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_3_sram_inv ) , 
    .out ( chany_top_out[8] ) , .p0 ( optlc_net_110 ) ) ;
mux_tree_tapbuf_size2_12 mux_top_track_18 (
    .in ( { top_left_grid_pin_39_[0] , chanx_left_in[11] } ) ,
    .sram ( mux_tree_tapbuf_size2_4_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_4_sram_inv ) , 
    .out ( chany_top_out[9] ) , .p0 ( optlc_net_110 ) ) ;
mux_tree_tapbuf_size2_13 mux_top_track_20 (
    .in ( { top_left_grid_pin_40_[0] , chanx_left_in[10] } ) ,
    .sram ( mux_tree_tapbuf_size2_5_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_5_sram_inv ) , 
    .out ( chany_top_out[10] ) , .p0 ( optlc_net_113 ) ) ;
mux_tree_tapbuf_size2_14 mux_top_track_22 (
    .in ( { top_left_grid_pin_41_[0] , chanx_left_in[9] } ) ,
    .sram ( mux_tree_tapbuf_size2_6_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_6_sram_inv ) ,
    .out ( { ropt_net_121 } ) ,
    .p0 ( optlc_net_113 ) ) ;
mux_tree_tapbuf_size2_15 mux_top_track_26 (
    .in ( { top_left_grid_pin_35_[0] , chanx_left_in[7] } ) ,
    .sram ( mux_tree_tapbuf_size2_7_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_7_sram_inv ) , 
    .out ( chany_top_out[13] ) , .p0 ( optlc_net_113 ) ) ;
mux_tree_tapbuf_size2_16 mux_top_track_28 (
    .in ( { top_left_grid_pin_36_[0] , chanx_left_in[6] } ) ,
    .sram ( mux_tree_tapbuf_size2_8_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_8_sram_inv ) ,
    .out ( { ropt_net_128 } ) ,
    .p0 ( optlc_net_110 ) ) ;
mux_tree_tapbuf_size2_17 mux_top_track_30 (
    .in ( { top_left_grid_pin_37_[0] , chanx_left_in[5] } ) ,
    .sram ( mux_tree_tapbuf_size2_9_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_9_sram_inv ) , 
    .out ( chany_top_out[15] ) , .p0 ( optlc_net_113 ) ) ;
mux_tree_tapbuf_size2_18 mux_top_track_32 (
    .in ( { top_left_grid_pin_38_[0] , chanx_left_in[4] } ) ,
    .sram ( mux_tree_tapbuf_size2_10_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_10_sram_inv ) ,
    .out ( { ropt_net_118 } ) ,
    .p0 ( optlc_net_110 ) ) ;
mux_tree_tapbuf_size2_19 mux_top_track_34 (
    .in ( { top_left_grid_pin_39_[0] , chanx_left_in[3] } ) ,
    .sram ( mux_tree_tapbuf_size2_11_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_11_sram_inv ) , 
    .out ( chany_top_out[17] ) , .p0 ( optlc_net_110 ) ) ;
mux_tree_tapbuf_size2_20 mux_top_track_36 (
    .in ( { top_left_grid_pin_40_[0] , chanx_left_in[2] } ) ,
    .sram ( mux_tree_tapbuf_size2_12_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_12_sram_inv ) , 
    .out ( chany_top_out[18] ) , .p0 ( optlc_net_113 ) ) ;
mux_tree_tapbuf_size2_21 mux_top_track_38 (
    .in ( { top_left_grid_pin_41_[0] , chanx_left_in[1] } ) ,
    .sram ( mux_tree_tapbuf_size2_13_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_13_sram_inv ) , 
    .out ( chany_top_out[19] ) , .p0 ( optlc_net_113 ) ) ;
mux_tree_tapbuf_size2_0_4 mux_left_track_11 (
    .in ( { chany_top_in[15] , left_top_grid_pin_43_[0] } ) ,
    .sram ( mux_tree_tapbuf_size2_14_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_14_sram_inv ) , 
    .out ( chanx_left_out[5] ) , .p0 ( optlc_net_110 ) ) ;
mux_tree_tapbuf_size2_1_4 mux_left_track_13 (
    .in ( { chany_top_in[14] , left_top_grid_pin_44_[0] } ) ,
    .sram ( mux_tree_tapbuf_size2_15_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_15_sram_inv ) , 
    .out ( chanx_left_out[6] ) , .p0 ( optlc_net_112 ) ) ;
mux_tree_tapbuf_size2_2_4 mux_left_track_15 (
    .in ( { chany_top_in[13] , left_top_grid_pin_45_[0] } ) ,
    .sram ( mux_tree_tapbuf_size2_16_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_16_sram_inv ) , 
    .out ( chanx_left_out[7] ) , .p0 ( optlc_net_112 ) ) ;
mux_tree_tapbuf_size2_3_4 mux_left_track_17 (
    .in ( { chany_top_in[12] , left_top_grid_pin_46_[0] } ) ,
    .sram ( mux_tree_tapbuf_size2_17_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_17_sram_inv ) ,
    .out ( { ropt_net_117 } ) ,
    .p0 ( optlc_net_112 ) ) ;
mux_tree_tapbuf_size2_4_3 mux_left_track_19 (
    .in ( { chany_top_in[11] , left_top_grid_pin_47_[0] } ) ,
    .sram ( mux_tree_tapbuf_size2_18_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_18_sram_inv ) , 
    .out ( chanx_left_out[9] ) , .p0 ( optlc_net_112 ) ) ;
mux_tree_tapbuf_size2_5_3 mux_left_track_21 (
    .in ( { chany_top_in[10] , left_top_grid_pin_48_[0] } ) ,
    .sram ( mux_tree_tapbuf_size2_19_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_19_sram_inv ) , 
    .out ( chanx_left_out[10] ) , .p0 ( optlc_net_112 ) ) ;
mux_tree_tapbuf_size2_6_2 mux_left_track_23 (
    .in ( { chany_top_in[9] , left_top_grid_pin_49_[0] } ) ,
    .sram ( mux_tree_tapbuf_size2_20_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_20_sram_inv ) , 
    .out ( chanx_left_out[11] ) , .p0 ( optlc_net_113 ) ) ;
mux_tree_tapbuf_size2_7_1 mux_left_track_27 (
    .in ( { chany_top_in[7] , left_top_grid_pin_43_[0] } ) ,
    .sram ( mux_tree_tapbuf_size2_21_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_21_sram_inv ) , 
    .out ( chanx_left_out[13] ) , .p0 ( optlc_net_110 ) ) ;
mux_tree_tapbuf_size2_mem_8_1 mem_top_track_10 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size3_mem_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_0_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_0_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_0_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem_9_1 mem_top_track_12 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_1_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_1_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_1_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem_10_1 mem_top_track_14 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_1_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_2_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_2_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_2_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem_11 mem_top_track_16 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_2_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_3_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_3_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_3_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem_12 mem_top_track_18 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_3_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_4_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_4_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_4_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem_13 mem_top_track_20 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_4_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_5_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_5_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_5_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem_14 mem_top_track_22 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_5_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_6_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_6_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_6_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem_15 mem_top_track_26 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size3_mem_1_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_7_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_7_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_7_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem_16 mem_top_track_28 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_7_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_8_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_8_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_8_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem_17 mem_top_track_30 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_8_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_9_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_9_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_9_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem_18 mem_top_track_32 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_9_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_10_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_10_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_10_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem_19 mem_top_track_34 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_10_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_11_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_11_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_11_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem_20 mem_top_track_36 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_11_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_12_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_12_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_12_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem_21 mem_top_track_38 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_12_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_13_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_13_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_13_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem_0_4 mem_left_track_11 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size3_mem_2_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_14_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_14_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_14_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem_1_4 mem_left_track_13 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_14_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_15_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_15_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_15_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem_2_4 mem_left_track_15 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_15_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_16_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_16_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_16_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem_3_4 mem_left_track_17 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_16_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_17_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_17_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_17_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem_4_3 mem_left_track_19 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_17_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_18_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_18_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_18_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem_5_3 mem_left_track_21 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_18_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_19_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_19_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_19_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem_6_2 mem_left_track_23 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_19_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_20_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_20_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_20_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem_7_1 mem_left_track_27 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size3_mem_3_ccff_tail ) ,
    .ccff_tail ( { ropt_net_129 } ) ,
    .mem_out ( mux_tree_tapbuf_size2_21_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_21_sram_inv ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_708 ( .A ( ropt_net_135 ) , 
    .X ( chanx_left_out[15] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_2__1 ( .A ( chany_top_in[2] ) , 
    .X ( chanx_left_out[18] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_709 ( .A ( ropt_net_136 ) , 
    .X ( chanx_left_out[19] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_710 ( .A ( ropt_net_137 ) , 
    .X ( chanx_left_out[16] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_711 ( .A ( ropt_net_138 ) , 
    .X ( chanx_left_out[14] ) ) ;
sky130_fd_sc_hd__conb_1 optlc_98 ( .LO ( SYNOPSYS_UNCONNECTED_1 ) , 
    .HI ( optlc_net_110 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_100 ( .LO ( SYNOPSYS_UNCONNECTED_2 ) , 
    .HI ( optlc_net_111 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_P_79 ( .A ( chany_top_in[6] ) , 
    .X ( ropt_net_127 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_P_86 ( .A ( chany_top_in[1] ) , 
    .X ( ropt_net_119 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_102 ( .LO ( SYNOPSYS_UNCONNECTED_3 ) , 
    .HI ( optlc_net_112 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_104 ( .LO ( SYNOPSYS_UNCONNECTED_4 ) , 
    .HI ( optlc_net_113 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_694 ( .A ( ropt_net_117 ) , 
    .X ( ropt_net_142 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_695 ( .A ( ropt_net_118 ) , 
    .X ( ropt_net_139 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_696 ( .A ( ropt_net_119 ) , 
    .X ( ropt_net_136 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_697 ( .A ( ropt_net_120 ) , 
    .X ( ropt_net_141 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_698 ( .A ( ropt_net_121 ) , 
    .X ( ropt_net_143 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_699 ( .A ( ropt_net_122 ) , 
    .X ( ropt_net_144 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_700 ( .A ( ropt_net_123 ) , 
    .X ( chany_top_out[12] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_701 ( .A ( chany_top_in[3] ) , 
    .X ( ropt_net_145 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_702 ( .A ( chany_top_in[4] ) , 
    .X ( ropt_net_137 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_703 ( .A ( chany_top_in[5] ) , 
    .X ( ropt_net_135 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_704 ( .A ( ropt_net_127 ) , 
    .X ( ropt_net_138 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_705 ( .A ( ropt_net_128 ) , 
    .X ( chany_top_out[14] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_706 ( .A ( ropt_net_129 ) , 
    .X ( ropt_net_140 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_712 ( .A ( ropt_net_139 ) , 
    .X ( chany_top_out[16] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_713 ( .A ( ropt_net_140 ) , 
    .X ( ccff_tail[0] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_714 ( .A ( ropt_net_141 ) , 
    .X ( chanx_left_out[2] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_715 ( .A ( ropt_net_142 ) , 
    .X ( chanx_left_out[8] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_716 ( .A ( ropt_net_143 ) , 
    .X ( chany_top_out[11] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_717 ( .A ( ropt_net_144 ) , 
    .X ( chany_top_out[4] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_718 ( .A ( ropt_net_145 ) , 
    .X ( chanx_left_out[17] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_14 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_34__59 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_5_2 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_33__58 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_4_2 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_32__57 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_3_3 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_31__56 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_2_3 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_30__55 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_1_3 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_29__54 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_0_3 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_28__53 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_36 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_14 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_36 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
endmodule


module const1_32 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_5_2 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_32 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
endmodule


module const1_31_1 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_4_2 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_31_1 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
endmodule


module const1_30_2 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_3_3 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_30_2 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
endmodule


module const1_29_2 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_2_3 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_29_2 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
endmodule


module const1_28_2 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_1_3 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_28_2 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
endmodule


module const1_27_2 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_0_3 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_27_2 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
endmodule


module mux_tree_tapbuf_size4_mem_7 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_27__52 ( .A ( mem_out[2] ) , 
    .X ( net_net_87 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_87 ( .A ( net_net_87 ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size4_mem_1_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_26__51 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size4_mem_0_2 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_25__50 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size4_mem_2_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_24__49 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_26_4 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size4_7 ( in , sram , sram_inv , out , p0 ) ;
input  [0:3] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;

const1_26_4 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( in[2] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , .A1 ( in[3] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
endmodule


module const1_25_4 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size4_1_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:3] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;

const1_25_4 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( in[2] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , .A1 ( in[3] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
endmodule


module const1_24_4 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size4_0_2 ( in , sram , sram_inv , out , p0 ) ;
input  [0:3] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;

const1_24_4 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( in[2] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , .A1 ( in[3] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
endmodule


module const1_23_4 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size4_2_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:3] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;

const1_23_4 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( in[2] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , .A1 ( in[3] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
endmodule


module mux_tree_tapbuf_size7_mem_7 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_23__48 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size7_mem_2_2 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_22__47 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size7_mem_1_3 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_21__46 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size7_mem_0_3 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_20__45 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_22_4 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size7_7 ( in , sram , sram_inv , out , p0 ) ;
input  [0:6] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;

const1_22_4 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_3_ ( .A0 ( p0 ) , .A1 ( in[6] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
endmodule


module const1_21_4 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size7_2_2 ( in , sram , sram_inv , out , p0 ) ;
input  [0:6] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;

const1_21_4 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_3_ ( .A0 ( p0 ) , .A1 ( in[6] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_66 ( 
    .A ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , .X ( BUF_net_66 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_118 ( .A ( BUF_net_66 ) , 
    .X ( out[0] ) ) ;
endmodule


module const1_20_4 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size7_1_3 ( in , sram , sram_inv , out , p0 ) ;
input  [0:6] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;

const1_20_4 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_3_ ( .A0 ( p0 ) , .A1 ( in[6] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
endmodule


module const1_19_4 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size7_0_3 ( in , sram , sram_inv , out , p0 ) ;
input  [0:6] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;

const1_19_4 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_3_ ( .A0 ( p0 ) , .A1 ( in[6] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
endmodule


module mux_tree_tapbuf_size3_mem_5_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_19__44 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size3_mem_4_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_18__43 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size3_mem_3_2 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_17__42 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size3_mem_2_2 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_16__41 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size3_mem_1_2 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_15__40 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size3_mem_0_3 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_14__39 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size3_mem_8 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_13__38 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_18_4 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size3_5_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:2] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;

const1_18_4 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( p0 ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
endmodule


module const1_17_4 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size3_4_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:2] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;

const1_17_4 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( p0 ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
endmodule


module const1_16_5 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size3_3_2 ( in , sram , sram_inv , out , p0 ) ;
input  [0:2] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;

const1_16_5 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( p0 ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
endmodule


module const1_15_5 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size3_2_2 ( in , sram , sram_inv , out , p0 ) ;
input  [0:2] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;

const1_15_5 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( p0 ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
endmodule


module const1_14_5 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size3_1_2 ( in , sram , sram_inv , out , p0 ) ;
input  [0:2] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;

const1_14_5 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( p0 ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
endmodule


module const1_13_5 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size3_0_3 ( in , sram , sram_inv , out , p0 ) ;
input  [0:2] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;

const1_13_5 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( p0 ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
endmodule


module const1_12_5 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size3_8 ( in , sram , sram_inv , out , p0 ) ;
input  [0:2] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;

const1_12_5 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( p0 ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
endmodule


module mux_tree_tapbuf_size5_mem_2_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_12__37 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size5_mem_1_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_11__36 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size5_mem_3_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_10__35 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size5_mem_0_2 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_9__34 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size5_mem_6 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_8__33 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size5_mem_4 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_7__32 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size5_mem_5 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_6__31 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_11_5 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size5_2_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:4] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;

const1_11_5 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , .A1 ( in[4] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_64 ( 
    .A ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .X ( out[0] ) ) ;
endmodule


module const1_10_5 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size5_1_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:4] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;

const1_10_5 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , .A1 ( in[4] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_63 ( 
    .A ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .X ( out[0] ) ) ;
endmodule


module const1_9_5 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size5_3_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:4] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;

const1_9_5 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , .A1 ( in[4] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
endmodule


module const1_8_5 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size5_0_2 ( in , sram , sram_inv , out , p0 ) ;
input  [0:4] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;

const1_8_5 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , .A1 ( in[4] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_8 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[2] ) , .X ( out[0] ) ) ;
endmodule


module const1_7_5 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size5_6 ( in , sram , sram_inv , out , p0 ) ;
input  [0:4] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;

const1_7_5 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , .A1 ( in[4] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
endmodule


module const1_6_6 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size5_4 ( in , sram , sram_inv , out , p0 ) ;
input  [0:4] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;

const1_6_6 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , .A1 ( in[4] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
endmodule


module const1_5_6 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size5_5 ( in , sram , sram_inv , out , p0 ) ;
input  [0:4] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;

const1_5_6 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , .A1 ( in[4] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
endmodule


module mux_tree_tapbuf_size6_mem_1_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_5__30 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size6_mem_0_3 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_4__29 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size6_mem_7 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_3__28 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size6_mem_3_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_2__27 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size6_mem_2_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_1__26 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_4_6 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size6_1_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:5] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;

const1_4_6 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
endmodule


module const1_3_6 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size6_0_3 ( in , sram , sram_inv , out , p0 ) ;
input  [0:5] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;

const1_3_6 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
endmodule


module const1_2_6 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size6_7 ( in , sram , sram_inv , out , p0 ) ;
input  [0:5] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;

const1_2_6 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_8 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , .X ( out[0] ) ) ;
endmodule


module const1_1_6 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size6_3_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:5] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;

const1_1_6 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
endmodule


module const1_0_6 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size6_2_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:5] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;

const1_0_6 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
endmodule


module sb_1__2_ ( prog_clk , chanx_right_in , right_top_grid_pin_1_ , 
    chany_bottom_in , bottom_left_grid_pin_34_ , bottom_left_grid_pin_35_ , 
    bottom_left_grid_pin_36_ , bottom_left_grid_pin_37_ , 
    bottom_left_grid_pin_38_ , bottom_left_grid_pin_39_ , 
    bottom_left_grid_pin_40_ , bottom_left_grid_pin_41_ , chanx_left_in , 
    left_top_grid_pin_1_ , ccff_head , chanx_right_out , chany_bottom_out , 
    chanx_left_out , ccff_tail ) ;
input  [0:0] prog_clk ;
input  [0:19] chanx_right_in ;
input  [0:0] right_top_grid_pin_1_ ;
input  [0:19] chany_bottom_in ;
input  [0:0] bottom_left_grid_pin_34_ ;
input  [0:0] bottom_left_grid_pin_35_ ;
input  [0:0] bottom_left_grid_pin_36_ ;
input  [0:0] bottom_left_grid_pin_37_ ;
input  [0:0] bottom_left_grid_pin_38_ ;
input  [0:0] bottom_left_grid_pin_39_ ;
input  [0:0] bottom_left_grid_pin_40_ ;
input  [0:0] bottom_left_grid_pin_41_ ;
input  [0:19] chanx_left_in ;
input  [0:0] left_top_grid_pin_1_ ;
input  [0:0] ccff_head ;
output [0:19] chanx_right_out ;
output [0:19] chany_bottom_out ;
output [0:19] chanx_left_out ;
output [0:0] ccff_tail ;

wire [0:1] mux_tree_tapbuf_size2_0_sram ;
wire [0:1] mux_tree_tapbuf_size2_0_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_1_sram ;
wire [0:1] mux_tree_tapbuf_size2_1_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_2_sram ;
wire [0:1] mux_tree_tapbuf_size2_2_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_3_sram ;
wire [0:1] mux_tree_tapbuf_size2_3_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_4_sram ;
wire [0:1] mux_tree_tapbuf_size2_4_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_5_sram ;
wire [0:1] mux_tree_tapbuf_size2_5_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_6_sram ;
wire [0:1] mux_tree_tapbuf_size2_6_sram_inv ;
wire [0:0] mux_tree_tapbuf_size2_mem_0_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_1_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_2_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_3_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_4_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_5_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_6_ccff_tail ;
wire [0:1] mux_tree_tapbuf_size3_0_sram ;
wire [0:1] mux_tree_tapbuf_size3_0_sram_inv ;
wire [0:1] mux_tree_tapbuf_size3_1_sram ;
wire [0:1] mux_tree_tapbuf_size3_1_sram_inv ;
wire [0:1] mux_tree_tapbuf_size3_2_sram ;
wire [0:1] mux_tree_tapbuf_size3_2_sram_inv ;
wire [0:1] mux_tree_tapbuf_size3_3_sram ;
wire [0:1] mux_tree_tapbuf_size3_3_sram_inv ;
wire [0:1] mux_tree_tapbuf_size3_4_sram ;
wire [0:1] mux_tree_tapbuf_size3_4_sram_inv ;
wire [0:1] mux_tree_tapbuf_size3_5_sram ;
wire [0:1] mux_tree_tapbuf_size3_5_sram_inv ;
wire [0:1] mux_tree_tapbuf_size3_6_sram ;
wire [0:1] mux_tree_tapbuf_size3_6_sram_inv ;
wire [0:0] mux_tree_tapbuf_size3_mem_0_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size3_mem_1_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size3_mem_2_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size3_mem_3_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size3_mem_4_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size3_mem_5_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size3_mem_6_ccff_tail ;
wire [0:2] mux_tree_tapbuf_size4_0_sram ;
wire [0:2] mux_tree_tapbuf_size4_0_sram_inv ;
wire [0:2] mux_tree_tapbuf_size4_1_sram ;
wire [0:2] mux_tree_tapbuf_size4_1_sram_inv ;
wire [0:2] mux_tree_tapbuf_size4_2_sram ;
wire [0:2] mux_tree_tapbuf_size4_2_sram_inv ;
wire [0:2] mux_tree_tapbuf_size4_3_sram ;
wire [0:2] mux_tree_tapbuf_size4_3_sram_inv ;
wire [0:0] mux_tree_tapbuf_size4_mem_0_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size4_mem_1_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size4_mem_2_ccff_tail ;
wire [0:2] mux_tree_tapbuf_size5_0_sram ;
wire [0:2] mux_tree_tapbuf_size5_0_sram_inv ;
wire [0:2] mux_tree_tapbuf_size5_1_sram ;
wire [0:2] mux_tree_tapbuf_size5_1_sram_inv ;
wire [0:2] mux_tree_tapbuf_size5_2_sram ;
wire [0:2] mux_tree_tapbuf_size5_2_sram_inv ;
wire [0:2] mux_tree_tapbuf_size5_3_sram ;
wire [0:2] mux_tree_tapbuf_size5_3_sram_inv ;
wire [0:2] mux_tree_tapbuf_size5_4_sram ;
wire [0:2] mux_tree_tapbuf_size5_4_sram_inv ;
wire [0:2] mux_tree_tapbuf_size5_5_sram ;
wire [0:2] mux_tree_tapbuf_size5_5_sram_inv ;
wire [0:2] mux_tree_tapbuf_size5_6_sram ;
wire [0:2] mux_tree_tapbuf_size5_6_sram_inv ;
wire [0:0] mux_tree_tapbuf_size5_mem_0_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size5_mem_1_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size5_mem_2_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size5_mem_3_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size5_mem_4_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size5_mem_5_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size5_mem_6_ccff_tail ;
wire [0:2] mux_tree_tapbuf_size6_0_sram ;
wire [0:2] mux_tree_tapbuf_size6_0_sram_inv ;
wire [0:2] mux_tree_tapbuf_size6_1_sram ;
wire [0:2] mux_tree_tapbuf_size6_1_sram_inv ;
wire [0:2] mux_tree_tapbuf_size6_2_sram ;
wire [0:2] mux_tree_tapbuf_size6_2_sram_inv ;
wire [0:2] mux_tree_tapbuf_size6_3_sram ;
wire [0:2] mux_tree_tapbuf_size6_3_sram_inv ;
wire [0:2] mux_tree_tapbuf_size6_4_sram ;
wire [0:2] mux_tree_tapbuf_size6_4_sram_inv ;
wire [0:0] mux_tree_tapbuf_size6_mem_0_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size6_mem_1_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size6_mem_2_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size6_mem_3_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size6_mem_4_ccff_tail ;
wire [0:2] mux_tree_tapbuf_size7_0_sram ;
wire [0:2] mux_tree_tapbuf_size7_0_sram_inv ;
wire [0:2] mux_tree_tapbuf_size7_1_sram ;
wire [0:2] mux_tree_tapbuf_size7_1_sram_inv ;
wire [0:2] mux_tree_tapbuf_size7_2_sram ;
wire [0:2] mux_tree_tapbuf_size7_2_sram_inv ;
wire [0:2] mux_tree_tapbuf_size7_3_sram ;
wire [0:2] mux_tree_tapbuf_size7_3_sram_inv ;
wire [0:0] mux_tree_tapbuf_size7_mem_0_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size7_mem_1_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size7_mem_2_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size7_mem_3_ccff_tail ;

mux_tree_tapbuf_size6_2_1 mux_right_track_0 (
    .in ( { right_top_grid_pin_1_[0] , chany_bottom_in[5] , 
        chany_bottom_in[12] , chany_bottom_in[19] , chanx_left_in[2] , 
        chanx_left_in[12] } ) ,
    .sram ( mux_tree_tapbuf_size6_0_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size6_0_sram_inv ) , 
    .out ( chanx_right_out[0] ) , .p0 ( optlc_net_135 ) ) ;
mux_tree_tapbuf_size6_3_1 mux_right_track_4 (
    .in ( { right_top_grid_pin_1_[0] , chany_bottom_in[3] , 
        chany_bottom_in[10] , chany_bottom_in[17] , chanx_left_in[5] , 
        chanx_left_in[14] } ) ,
    .sram ( mux_tree_tapbuf_size6_1_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size6_1_sram_inv ) , 
    .out ( chanx_right_out[2] ) , .p0 ( optlc_net_135 ) ) ;
mux_tree_tapbuf_size6_7 mux_right_track_8 (
    .in ( { right_top_grid_pin_1_[0] , chany_bottom_in[2] , 
        chany_bottom_in[9] , chany_bottom_in[16] , chanx_left_in[6] , 
        chanx_left_in[16] } ) ,
    .sram ( mux_tree_tapbuf_size6_2_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size6_2_sram_inv ) , 
    .out ( chanx_right_out[4] ) , .p0 ( optlc_net_135 ) ) ;
mux_tree_tapbuf_size6_0_3 mux_left_track_5 (
    .in ( { chanx_right_in[5] , chanx_right_in[14] , chany_bottom_in[1] , 
        chany_bottom_in[8] , chany_bottom_in[15] , left_top_grid_pin_1_[0] } ) ,
    .sram ( mux_tree_tapbuf_size6_3_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size6_3_sram_inv ) , 
    .out ( chanx_left_out[2] ) , .p0 ( optlc_net_136 ) ) ;
mux_tree_tapbuf_size6_1_1 mux_left_track_9 (
    .in ( { chanx_right_in[6] , chanx_right_in[16] , chany_bottom_in[2] , 
        chany_bottom_in[9] , chany_bottom_in[16] , left_top_grid_pin_1_[0] } ) ,
    .sram ( mux_tree_tapbuf_size6_4_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size6_4_sram_inv ) , 
    .out ( chanx_left_out[4] ) , .p0 ( optlc_net_136 ) ) ;
mux_tree_tapbuf_size6_mem_2_1 mem_right_track_0 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( ccff_head ) , 
    .ccff_tail ( mux_tree_tapbuf_size6_mem_0_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size6_0_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size6_0_sram_inv ) ) ;
mux_tree_tapbuf_size6_mem_3_1 mem_right_track_4 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size5_mem_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size6_mem_1_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size6_1_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size6_1_sram_inv ) ) ;
mux_tree_tapbuf_size6_mem_7 mem_right_track_8 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size6_mem_1_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size6_mem_2_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size6_2_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size6_2_sram_inv ) ) ;
mux_tree_tapbuf_size6_mem_0_3 mem_left_track_5 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size5_mem_4_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size6_mem_3_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size6_3_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size6_3_sram_inv ) ) ;
mux_tree_tapbuf_size6_mem_1_1 mem_left_track_9 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size6_mem_3_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size6_mem_4_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size6_4_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size6_4_sram_inv ) ) ;
mux_tree_tapbuf_size5_5 mux_right_track_2 (
    .in ( { chany_bottom_in[4] , chany_bottom_in[11] , chany_bottom_in[18] , 
        chanx_left_in[4] , chanx_left_in[13] } ) ,
    .sram ( mux_tree_tapbuf_size5_0_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size5_0_sram_inv ) , 
    .out ( chanx_right_out[1] ) , .p0 ( optlc_net_135 ) ) ;
mux_tree_tapbuf_size5_4 mux_right_track_16 (
    .in ( { chany_bottom_in[1] , chany_bottom_in[8] , chany_bottom_in[15] , 
        chanx_left_in[8] , chanx_left_in[17] } ) ,
    .sram ( mux_tree_tapbuf_size5_1_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size5_1_sram_inv ) , 
    .out ( chanx_right_out[8] ) , .p0 ( optlc_net_136 ) ) ;
mux_tree_tapbuf_size5_6 mux_right_track_24 (
    .in ( { chany_bottom_in[0] , chany_bottom_in[7] , chany_bottom_in[14] , 
        chanx_left_in[9] , chanx_left_in[18] } ) ,
    .sram ( mux_tree_tapbuf_size5_2_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size5_2_sram_inv ) , 
    .out ( chanx_right_out[12] ) , .p0 ( optlc_net_135 ) ) ;
mux_tree_tapbuf_size5_0_2 mux_left_track_1 (
    .in ( { chanx_right_in[2] , chanx_right_in[12] , chany_bottom_in[6] , 
        chany_bottom_in[13] , left_top_grid_pin_1_[0] } ) ,
    .sram ( mux_tree_tapbuf_size5_3_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size5_3_sram_inv ) , 
    .out ( chanx_left_out[0] ) , .p0 ( optlc_net_136 ) ) ;
mux_tree_tapbuf_size5_3_1 mux_left_track_3 (
    .in ( { chanx_right_in[4] , chanx_right_in[13] , chany_bottom_in[0] , 
        chany_bottom_in[7] , chany_bottom_in[14] } ) ,
    .sram ( mux_tree_tapbuf_size5_4_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size5_4_sram_inv ) , 
    .out ( chanx_left_out[1] ) , .p0 ( optlc_net_137 ) ) ;
mux_tree_tapbuf_size5_1_1 mux_left_track_17 (
    .in ( { chanx_right_in[8] , chanx_right_in[17] , chany_bottom_in[3] , 
        chany_bottom_in[10] , chany_bottom_in[17] } ) ,
    .sram ( mux_tree_tapbuf_size5_5_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size5_5_sram_inv ) ,
    .out ( { ropt_net_140 } ) ,
    .p0 ( optlc_net_135 ) ) ;
mux_tree_tapbuf_size5_2_1 mux_left_track_25 (
    .in ( { chanx_right_in[9] , chanx_right_in[18] , chany_bottom_in[4] , 
        chany_bottom_in[11] , chany_bottom_in[18] } ) ,
    .sram ( mux_tree_tapbuf_size5_6_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size5_6_sram_inv ) ,
    .out ( { ropt_net_139 } ) ,
    .p0 ( optlc_net_135 ) ) ;
mux_tree_tapbuf_size5_mem_5 mem_right_track_2 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size6_mem_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size5_mem_0_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size5_0_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size5_0_sram_inv ) ) ;
mux_tree_tapbuf_size5_mem_4 mem_right_track_16 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size6_mem_2_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size5_mem_1_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size5_1_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size5_1_sram_inv ) ) ;
mux_tree_tapbuf_size5_mem_6 mem_right_track_24 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size5_mem_1_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size5_mem_2_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size5_2_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size5_2_sram_inv ) ) ;
mux_tree_tapbuf_size5_mem_0_2 mem_left_track_1 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_6_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size5_mem_3_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size5_3_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size5_3_sram_inv ) ) ;
mux_tree_tapbuf_size5_mem_3_1 mem_left_track_3 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size5_mem_3_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size5_mem_4_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size5_4_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size5_4_sram_inv ) ) ;
mux_tree_tapbuf_size5_mem_1_1 mem_left_track_17 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size6_mem_4_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size5_mem_5_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size5_5_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size5_5_sram_inv ) ) ;
mux_tree_tapbuf_size5_mem_2_1 mem_left_track_25 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size5_mem_5_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size5_mem_6_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size5_6_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size5_6_sram_inv ) ) ;
mux_tree_tapbuf_size3_8 mux_right_track_32 (
    .in ( { chany_bottom_in[6] , chany_bottom_in[13] , chanx_left_in[10] } ) ,
    .sram ( mux_tree_tapbuf_size3_0_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size3_0_sram_inv ) , 
    .out ( chanx_right_out[16] ) , .p0 ( optlc_net_137 ) ) ;
mux_tree_tapbuf_size3_0_3 mux_bottom_track_13 (
    .in ( { chanx_right_in[10] , bottom_left_grid_pin_36_[0] , 
        chanx_left_in[10] } ) ,
    .sram ( mux_tree_tapbuf_size3_1_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size3_1_sram_inv ) , 
    .out ( chany_bottom_out[6] ) , .p0 ( optlc_net_137 ) ) ;
mux_tree_tapbuf_size3_1_2 mux_bottom_track_15 (
    .in ( { chanx_right_in[12] , bottom_left_grid_pin_37_[0] , 
        chanx_left_in[12] } ) ,
    .sram ( mux_tree_tapbuf_size3_2_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size3_2_sram_inv ) , 
    .out ( chany_bottom_out[7] ) , .p0 ( optlc_net_137 ) ) ;
mux_tree_tapbuf_size3_2_2 mux_bottom_track_17 (
    .in ( { chanx_right_in[13] , bottom_left_grid_pin_38_[0] , 
        chanx_left_in[13] } ) ,
    .sram ( mux_tree_tapbuf_size3_3_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size3_3_sram_inv ) , 
    .out ( chany_bottom_out[8] ) , .p0 ( optlc_net_137 ) ) ;
mux_tree_tapbuf_size3_3_2 mux_bottom_track_19 (
    .in ( { chanx_right_in[14] , bottom_left_grid_pin_39_[0] , 
        chanx_left_in[14] } ) ,
    .sram ( mux_tree_tapbuf_size3_4_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size3_4_sram_inv ) , 
    .out ( chany_bottom_out[9] ) , .p0 ( optlc_net_137 ) ) ;
mux_tree_tapbuf_size3_4_1 mux_bottom_track_21 (
    .in ( { chanx_right_in[16] , bottom_left_grid_pin_40_[0] , 
        chanx_left_in[16] } ) ,
    .sram ( mux_tree_tapbuf_size3_5_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size3_5_sram_inv ) , 
    .out ( chany_bottom_out[10] ) , .p0 ( optlc_net_135 ) ) ;
mux_tree_tapbuf_size3_5_1 mux_bottom_track_23 (
    .in ( { chanx_right_in[17] , bottom_left_grid_pin_41_[0] , 
        chanx_left_in[17] } ) ,
    .sram ( mux_tree_tapbuf_size3_6_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size3_6_sram_inv ) , 
    .out ( chany_bottom_out[11] ) , .p0 ( optlc_net_138 ) ) ;
mux_tree_tapbuf_size3_mem_8 mem_right_track_32 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size5_mem_2_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size3_mem_0_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size3_0_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size3_0_sram_inv ) ) ;
mux_tree_tapbuf_size3_mem_0_3 mem_bottom_track_13 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size4_mem_1_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size3_mem_1_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size3_1_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size3_1_sram_inv ) ) ;
mux_tree_tapbuf_size3_mem_1_2 mem_bottom_track_15 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size3_mem_1_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size3_mem_2_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size3_2_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size3_2_sram_inv ) ) ;
mux_tree_tapbuf_size3_mem_2_2 mem_bottom_track_17 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size3_mem_2_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size3_mem_3_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size3_3_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size3_3_sram_inv ) ) ;
mux_tree_tapbuf_size3_mem_3_2 mem_bottom_track_19 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size3_mem_3_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size3_mem_4_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size3_4_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size3_4_sram_inv ) ) ;
mux_tree_tapbuf_size3_mem_4_1 mem_bottom_track_21 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size3_mem_4_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size3_mem_5_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size3_5_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size3_5_sram_inv ) ) ;
mux_tree_tapbuf_size3_mem_5_1 mem_bottom_track_23 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size3_mem_5_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size3_mem_6_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size3_6_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size3_6_sram_inv ) ) ;
mux_tree_tapbuf_size7_0_3 mux_bottom_track_1 (
    .in ( { chanx_right_in[2] , bottom_left_grid_pin_34_[0] , 
        bottom_left_grid_pin_36_[0] , bottom_left_grid_pin_38_[0] , 
        bottom_left_grid_pin_40_[0] , chanx_left_in[1] , chanx_left_in[2] } ) ,
    .sram ( mux_tree_tapbuf_size7_0_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size7_0_sram_inv ) , 
    .out ( chany_bottom_out[0] ) , .p0 ( optlc_net_137 ) ) ;
mux_tree_tapbuf_size7_1_3 mux_bottom_track_3 (
    .in ( { chanx_right_in[4] , bottom_left_grid_pin_35_[0] , 
        bottom_left_grid_pin_37_[0] , bottom_left_grid_pin_39_[0] , 
        bottom_left_grid_pin_41_[0] , chanx_left_in[3] , chanx_left_in[4] } ) ,
    .sram ( mux_tree_tapbuf_size7_1_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size7_1_sram_inv ) , 
    .out ( chany_bottom_out[1] ) , .p0 ( optlc_net_136 ) ) ;
mux_tree_tapbuf_size7_2_2 mux_bottom_track_5 (
    .in ( { chanx_right_in[5] , bottom_left_grid_pin_34_[0] , 
        bottom_left_grid_pin_36_[0] , bottom_left_grid_pin_38_[0] , 
        bottom_left_grid_pin_40_[0] , chanx_left_in[5] , chanx_left_in[7] } ) ,
    .sram ( mux_tree_tapbuf_size7_2_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size7_2_sram_inv ) ,
    .out ( { ropt_net_145 } ) ,
    .p0 ( optlc_net_136 ) ) ;
mux_tree_tapbuf_size7_7 mux_bottom_track_7 (
    .in ( { chanx_right_in[6] , bottom_left_grid_pin_35_[0] , 
        bottom_left_grid_pin_37_[0] , bottom_left_grid_pin_39_[0] , 
        bottom_left_grid_pin_41_[0] , chanx_left_in[6] , chanx_left_in[11] } ) ,
    .sram ( mux_tree_tapbuf_size7_3_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size7_3_sram_inv ) , 
    .out ( chany_bottom_out[3] ) , .p0 ( optlc_net_136 ) ) ;
mux_tree_tapbuf_size7_mem_0_3 mem_bottom_track_1 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size3_mem_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size7_mem_0_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size7_0_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size7_0_sram_inv ) ) ;
mux_tree_tapbuf_size7_mem_1_3 mem_bottom_track_3 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size7_mem_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size7_mem_1_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size7_1_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size7_1_sram_inv ) ) ;
mux_tree_tapbuf_size7_mem_2_2 mem_bottom_track_5 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size7_mem_1_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size7_mem_2_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size7_2_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size7_2_sram_inv ) ) ;
mux_tree_tapbuf_size7_mem_7 mem_bottom_track_7 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size7_mem_2_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size7_mem_3_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size7_3_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size7_3_sram_inv ) ) ;
mux_tree_tapbuf_size4_2_1 mux_bottom_track_9 (
    .in ( { chanx_right_in[8] , bottom_left_grid_pin_34_[0] , 
        chanx_left_in[8] , chanx_left_in[15] } ) ,
    .sram ( mux_tree_tapbuf_size4_0_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size4_0_sram_inv ) , 
    .out ( chany_bottom_out[4] ) , .p0 ( optlc_net_136 ) ) ;
mux_tree_tapbuf_size4_0_2 mux_bottom_track_11 (
    .in ( { chanx_right_in[9] , bottom_left_grid_pin_35_[0] , 
        chanx_left_in[9] , chanx_left_in[19] } ) ,
    .sram ( mux_tree_tapbuf_size4_1_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size4_1_sram_inv ) , 
    .out ( chany_bottom_out[5] ) , .p0 ( optlc_net_136 ) ) ;
mux_tree_tapbuf_size4_1_1 mux_bottom_track_25 (
    .in ( { chanx_right_in[18] , chanx_right_in[19] , 
        bottom_left_grid_pin_34_[0] , chanx_left_in[18] } ) ,
    .sram ( mux_tree_tapbuf_size4_2_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size4_2_sram_inv ) , 
    .out ( chany_bottom_out[12] ) , .p0 ( optlc_net_138 ) ) ;
mux_tree_tapbuf_size4_7 mux_left_track_33 (
    .in ( { chanx_right_in[10] , chany_bottom_in[5] , chany_bottom_in[12] , 
        chany_bottom_in[19] } ) ,
    .sram ( mux_tree_tapbuf_size4_3_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size4_3_sram_inv ) , 
    .out ( chanx_left_out[16] ) , .p0 ( optlc_net_135 ) ) ;
mux_tree_tapbuf_size4_mem_2_1 mem_bottom_track_9 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size7_mem_3_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size4_mem_0_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size4_0_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size4_0_sram_inv ) ) ;
mux_tree_tapbuf_size4_mem_0_2 mem_bottom_track_11 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size4_mem_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size4_mem_1_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size4_1_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size4_1_sram_inv ) ) ;
mux_tree_tapbuf_size4_mem_1_1 mem_bottom_track_25 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size3_mem_6_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size4_mem_2_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size4_2_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size4_2_sram_inv ) ) ;
mux_tree_tapbuf_size4_mem_7 mem_left_track_33 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size5_mem_6_ccff_tail ) ,
    .ccff_tail ( { ropt_net_152 } ) ,
    .mem_out ( mux_tree_tapbuf_size4_3_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size4_3_sram_inv ) ) ;
mux_tree_tapbuf_size2_0_3 mux_bottom_track_27 (
    .in ( { chanx_right_in[15] , bottom_left_grid_pin_35_[0] } ) ,
    .sram ( mux_tree_tapbuf_size2_0_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_0_sram_inv ) , 
    .out ( chany_bottom_out[13] ) , .p0 ( optlc_net_138 ) ) ;
mux_tree_tapbuf_size2_1_3 mux_bottom_track_29 (
    .in ( { chanx_right_in[11] , bottom_left_grid_pin_36_[0] } ) ,
    .sram ( mux_tree_tapbuf_size2_1_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_1_sram_inv ) , 
    .out ( chany_bottom_out[14] ) , .p0 ( optlc_net_138 ) ) ;
mux_tree_tapbuf_size2_2_3 mux_bottom_track_31 (
    .in ( { chanx_right_in[7] , bottom_left_grid_pin_37_[0] } ) ,
    .sram ( mux_tree_tapbuf_size2_2_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_2_sram_inv ) , 
    .out ( chany_bottom_out[15] ) , .p0 ( optlc_net_137 ) ) ;
mux_tree_tapbuf_size2_3_3 mux_bottom_track_33 (
    .in ( { chanx_right_in[3] , bottom_left_grid_pin_38_[0] } ) ,
    .sram ( mux_tree_tapbuf_size2_3_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_3_sram_inv ) , 
    .out ( chany_bottom_out[16] ) , .p0 ( optlc_net_138 ) ) ;
mux_tree_tapbuf_size2_4_2 mux_bottom_track_35 (
    .in ( { chanx_right_in[1] , bottom_left_grid_pin_39_[0] } ) ,
    .sram ( mux_tree_tapbuf_size2_4_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_4_sram_inv ) , 
    .out ( chany_bottom_out[17] ) , .p0 ( optlc_net_138 ) ) ;
mux_tree_tapbuf_size2_5_2 mux_bottom_track_37 (
    .in ( { chanx_right_in[0] , bottom_left_grid_pin_40_[0] } ) ,
    .sram ( mux_tree_tapbuf_size2_5_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_5_sram_inv ) , 
    .out ( chany_bottom_out[18] ) , .p0 ( optlc_net_138 ) ) ;
mux_tree_tapbuf_size2_14 mux_bottom_track_39 (
    .in ( { bottom_left_grid_pin_41_[0] , chanx_left_in[0] } ) ,
    .sram ( mux_tree_tapbuf_size2_6_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_6_sram_inv ) , 
    .out ( chany_bottom_out[19] ) , .p0 ( optlc_net_137 ) ) ;
mux_tree_tapbuf_size2_mem_0_3 mem_bottom_track_27 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size4_mem_2_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_0_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_0_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_0_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem_1_3 mem_bottom_track_29 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_1_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_1_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_1_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem_2_3 mem_bottom_track_31 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_1_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_2_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_2_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_2_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem_3_3 mem_bottom_track_33 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_2_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_3_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_3_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_3_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem_4_2 mem_bottom_track_35 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_3_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_4_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_4_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_4_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem_5_2 mem_bottom_track_37 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_4_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_5_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_5_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_5_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem_14 mem_bottom_track_39 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_5_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_6_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_6_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_6_sram_inv ) ) ;
sky130_fd_sc_hd__conb_1 optlc_124 ( .LO ( SYNOPSYS_UNCONNECTED_1 ) , 
    .HI ( optlc_net_135 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_2__1 ( .A ( chanx_right_in[4] ) , 
    .X ( ropt_net_157 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_3__2 ( .A ( chanx_right_in[5] ) , 
    .X ( ropt_net_155 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_4__3 ( .A ( chanx_right_in[6] ) , 
    .X ( ropt_net_158 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_759 ( .A ( ropt_net_167 ) , 
    .X ( chanx_left_out[3] ) ) ;
sky130_fd_sc_hd__conb_1 optlc_126 ( .LO ( SYNOPSYS_UNCONNECTED_2 ) , 
    .HI ( optlc_net_136 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_760 ( .A ( ropt_net_168 ) , 
    .X ( chanx_left_out[12] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_725 ( .A ( ropt_net_139 ) , 
    .X ( ropt_net_168 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_761 ( .A ( ropt_net_169 ) , 
    .X ( ccff_tail[0] ) ) ;
sky130_fd_sc_hd__conb_1 optlc_128 ( .LO ( SYNOPSYS_UNCONNECTED_3 ) , 
    .HI ( optlc_net_137 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_130 ( .LO ( SYNOPSYS_UNCONNECTED_4 ) , 
    .HI ( optlc_net_138 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_762 ( .A ( ropt_net_170 ) , 
    .X ( chanx_left_out[5] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_13__12 ( .A ( chanx_right_in[18] ) , 
    .X ( ropt_net_182 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_14__13 ( .A ( chanx_left_in[2] ) , 
    .X ( ropt_net_162 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_726 ( .A ( ropt_net_140 ) , 
    .X ( ropt_net_175 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_727 ( .A ( chanx_right_in[14] ) , 
    .X ( chanx_left_out[15] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_728 ( .A ( chanx_left_in[10] ) , 
    .X ( chanx_right_out[11] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_729 ( .A ( ropt_net_143 ) , 
    .X ( ropt_net_172 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_730 ( .A ( chanx_right_in[2] ) , 
    .X ( ropt_net_167 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_731 ( .A ( ropt_net_145 ) , 
    .X ( ropt_net_171 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_21__20 ( .A ( chanx_left_in[12] ) , 
    .X ( ropt_net_161 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_22__21 ( .A ( chanx_left_in[13] ) , 
    .X ( ropt_net_183 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_732 ( .A ( chanx_right_in[10] ) , 
    .X ( chanx_left_out[11] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_733 ( .A ( chanx_right_in[16] ) , 
    .X ( chanx_left_out[17] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_25__24 ( .A ( chanx_left_in[17] ) , 
    .X ( ropt_net_163 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_26__25 ( .A ( chanx_left_in[18] ) , 
    .X ( ropt_net_159 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_734 ( .A ( chanx_right_in[8] ) , 
    .X ( chanx_left_out[9] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_735 ( .A ( chanx_right_in[17] ) , 
    .X ( chanx_left_out[18] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_736 ( .A ( ropt_net_150 ) , 
    .X ( ropt_net_174 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_763 ( .A ( ropt_net_171 ) , 
    .X ( chany_bottom_out[2] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_764 ( .A ( ropt_net_172 ) , 
    .X ( chanx_left_out[14] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_765 ( .A ( ropt_net_173 ) , 
    .X ( chanx_right_out[17] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_766 ( .A ( ropt_net_174 ) , 
    .X ( chanx_right_out[7] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_767 ( .A ( ropt_net_175 ) , 
    .X ( chanx_left_out[8] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_79 ( .A ( chanx_left_in[5] ) , 
    .X ( ropt_net_153 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_80 ( .A ( chanx_left_in[6] ) , 
    .X ( ropt_net_150 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_737 ( .A ( chanx_left_in[4] ) , 
    .X ( chanx_right_out[5] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_82 ( .A ( chanx_left_in[9] ) , 
    .X ( ropt_net_154 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_768 ( .A ( ropt_net_176 ) , 
    .X ( chanx_right_out[10] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_RR_84 ( .A ( chanx_left_in[14] ) , 
    .X ( chanx_right_out[15] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_85 ( .A ( chanx_left_in[16] ) , 
    .X ( ropt_net_160 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_769 ( .A ( ropt_net_177 ) , 
    .X ( chanx_right_out[13] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_738 ( .A ( ropt_net_152 ) , 
    .X ( ropt_net_169 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_739 ( .A ( ropt_net_153 ) , 
    .X ( ropt_net_180 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_101 ( .A ( chanx_left_in[8] ) , 
    .X ( ropt_net_156 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_740 ( .A ( ropt_net_154 ) , 
    .X ( ropt_net_176 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_770 ( .A ( ropt_net_178 ) , 
    .X ( chanx_right_out[9] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_P_108 ( .A ( chanx_right_in[9] ) , 
    .X ( chanx_left_out[10] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_771 ( .A ( ropt_net_179 ) , 
    .X ( chanx_left_out[6] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_P_111 ( .A ( chanx_right_in[12] ) , 
    .X ( chanx_left_out[13] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_P_112 ( .A ( chanx_right_in[13] ) , 
    .X ( ropt_net_143 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_772 ( .A ( ropt_net_180 ) , 
    .X ( chanx_right_out[6] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_742 ( .A ( ropt_net_155 ) , 
    .X ( ropt_net_179 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_773 ( .A ( ropt_net_181 ) , 
    .X ( chanx_left_out[7] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_777 ( .A ( ropt_net_182 ) , 
    .X ( chanx_left_out[19] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_743 ( .A ( ropt_net_156 ) , 
    .X ( ropt_net_178 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_744 ( .A ( ropt_net_157 ) , 
    .X ( ropt_net_170 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_745 ( .A ( ropt_net_158 ) , 
    .X ( ropt_net_181 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_746 ( .A ( ropt_net_159 ) , 
    .X ( chanx_right_out[19] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_747 ( .A ( ropt_net_160 ) , 
    .X ( ropt_net_173 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_749 ( .A ( ropt_net_161 ) , 
    .X ( ropt_net_177 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_750 ( .A ( ropt_net_162 ) , 
    .X ( chanx_right_out[3] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_753 ( .A ( ropt_net_163 ) , 
    .X ( chanx_right_out[18] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_780 ( .A ( ropt_net_183 ) , 
    .X ( chanx_right_out[14] ) ) ;
endmodule


module mux_tree_tapbuf_size7_mem_1_2 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd1_1 FTB_28__79 ( .A ( mem_out[2] ) , 
    .X ( net_net_91 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 BUFT_RR_91 ( .A ( net_net_91 ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size7_mem_0_2 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_27__78 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size7_mem_2_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_26__77 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size7_mem_6 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_25__76 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_35 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size7_1_2 ( in , sram , sram_inv , out , p0 ) ;
input  [0:6] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;

const1_35 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_3_ ( .A0 ( p0 ) , .A1 ( in[6] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
endmodule


module const1_26_3 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size7_0_2 ( in , sram , sram_inv , out , p0 ) ;
input  [0:6] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;

const1_26_3 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_3_ ( .A0 ( p0 ) , .A1 ( in[6] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
endmodule


module const1_25_3 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size7_2_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:6] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;

const1_25_3 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_3_ ( .A0 ( p0 ) , .A1 ( in[6] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
endmodule


module const1_24_3 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size7_6 ( in , sram , sram_inv , out , p0 ) ;
input  [0:6] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;

const1_24_3 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_3_ ( .A0 ( p0 ) , .A1 ( in[6] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
endmodule


module mux_tree_tapbuf_size10_mem_4 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_24__75 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size10_mem_3 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_23__74 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size10_mem_5 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_22__73 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size10_mem_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_21__72 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size10_mem_0 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_20__71 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size10_mem_2 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_19__70 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size10_mem_7 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_18__69 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size10_mem_6 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_17__68 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size10_mem_8 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_16__67 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size10_mem_10 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_15__66 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size10_mem_9 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_14__65 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size10_mem_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_13__64 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_23_3 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size10_4 ( in , sram , sram_inv , out , p0 ) ;
input  [0:9] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

const1_23_3 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[6] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[8] ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[9] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
endmodule


module const1_22_3 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size10_3 ( in , sram , sram_inv , out , p0 ) ;
input  [0:9] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

const1_22_3 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[6] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[8] ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[9] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
endmodule


module const1_21_3 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size10_5 ( in , sram , sram_inv , out , p0 ) ;
input  [0:9] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

const1_21_3 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[6] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[8] ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[9] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
endmodule


module const1_20_3 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size10_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:9] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

const1_20_3 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[6] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[8] ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[9] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
endmodule


module const1_19_3 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size10_0 ( in , sram , sram_inv , out , p0 ) ;
input  [0:9] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

const1_19_3 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[6] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[8] ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[9] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
endmodule


module const1_18_3 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size10_2 ( in , sram , sram_inv , out , p0 ) ;
input  [0:9] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

const1_18_3 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[6] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[8] ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[9] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
endmodule


module const1_17_3 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size10_7 ( in , sram , sram_inv , out , p0 ) ;
input  [0:9] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;

const1_17_3 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[6] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[8] ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[9] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_4 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .S ( sram[3] ) , .X ( out[0] ) ) ;
endmodule


module const1_16_4 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size10_6 ( in , sram , sram_inv , out , p0 ) ;
input  [0:9] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

const1_16_4 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[6] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[8] ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[9] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
endmodule


module const1_15_4 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size10_8 ( in , sram , sram_inv , out , p0 ) ;
input  [0:9] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

const1_15_4 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[6] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[8] ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[9] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
endmodule


module const1_14_4 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size10_10 ( in , sram , sram_inv , out , p0 ) ;
input  [0:9] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

const1_14_4 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[6] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[8] ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[9] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
endmodule


module const1_13_4 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size10_9 ( in , sram , sram_inv , out , p0 ) ;
input  [0:9] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

const1_13_4 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[6] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[8] ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[9] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
endmodule


module const1_12_4 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size10_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:9] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

const1_12_4 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[6] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[8] ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[9] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
endmodule


module mux_tree_tapbuf_size16_mem_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:4] mem_out ;
output [0:4] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_4_ ( .D ( mem_out[3] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[4] ) , .Q_N ( mem_outb[4] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_12__63 ( .A ( mem_out[4] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size16_mem_0 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:4] mem_out ;
output [0:4] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_4_ ( .D ( mem_out[3] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[4] ) , .Q_N ( mem_outb[4] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_11__62 ( .A ( mem_out[4] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size16_mem_2 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:4] mem_out ;
output [0:4] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_4_ ( .D ( mem_out[3] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[4] ) , .Q_N ( mem_outb[4] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_10__61 ( .A ( mem_out[4] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size16_mem ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:4] mem_out ;
output [0:4] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_4_ ( .D ( mem_out[3] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[4] ) , .Q_N ( mem_outb[4] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_9__60 ( .A ( mem_out[4] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_11_4 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size16_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:15] in ;
input  [0:4] sram ;
input  [0:4] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_10_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_11_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_12_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_13_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_14_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_15_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

const1_11_4 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_15_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( in[2] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[4] ) , .A1 ( in[3] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[6] ) , .A1 ( in[5] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( in[8] ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_4_ ( .A0 ( in[10] ) , .A1 ( in[9] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_5_ ( .A0 ( in[12] ) , .A1 ( in[11] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_6_ ( .A0 ( in[14] ) , .A1 ( in[13] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_7_ ( .A0 ( p0 ) , .A1 ( in[15] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_10_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_2_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_11_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_3_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_12_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_10_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_13_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_12_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_11_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_14_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l5_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_14_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_13_X[0] ) , .S ( sram[4] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_15_X[0] ) ) ;
endmodule


module const1_10_4 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size16_0 ( in , sram , sram_inv , out , p0 ) ;
input  [0:15] in ;
input  [0:4] sram ;
input  [0:4] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_10_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_11_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_12_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_13_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_14_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_15_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

const1_10_4 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( in[2] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[4] ) , .A1 ( in[3] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[6] ) , .A1 ( in[5] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( in[8] ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_4_ ( .A0 ( in[10] ) , .A1 ( in[9] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_5_ ( .A0 ( in[12] ) , .A1 ( in[11] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_6_ ( .A0 ( in[14] ) , .A1 ( in[13] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_7_ ( .A0 ( p0 ) , .A1 ( in[15] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_10_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_2_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_11_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_3_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_12_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_10_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_13_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_12_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_11_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_14_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l5_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_14_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_13_X[0] ) , .S ( sram[4] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_15_X[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_81 ( 
    .A ( sky130_fd_sc_hd__mux2_1_15_X[0] ) , .X ( BUF_net_81 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 BUFT_RR_99 ( .A ( BUF_net_81 ) , 
    .X ( out[0] ) ) ;
endmodule


module const1_9_4 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size16_2 ( in , sram , sram_inv , out , p0 ) ;
input  [0:15] in ;
input  [0:4] sram ;
input  [0:4] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_10_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_11_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_12_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_13_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_14_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_15_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

const1_9_4 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_15_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( in[2] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[4] ) , .A1 ( in[3] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[6] ) , .A1 ( in[5] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( in[8] ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_4_ ( .A0 ( in[10] ) , .A1 ( in[9] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_5_ ( .A0 ( in[12] ) , .A1 ( in[11] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_6_ ( .A0 ( in[14] ) , .A1 ( in[13] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_7_ ( .A0 ( p0 ) , .A1 ( in[15] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_10_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_2_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_11_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_3_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_12_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_10_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_13_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_12_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_11_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_14_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l5_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_14_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_13_X[0] ) , .S ( sram[4] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_15_X[0] ) ) ;
endmodule


module const1_8_4 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size16 ( in , sram , sram_inv , out , p0 ) ;
input  [0:15] in ;
input  [0:4] sram ;
input  [0:4] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_10_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_11_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_12_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_13_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_14_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_15_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

const1_8_4 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_15_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( in[2] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[4] ) , .A1 ( in[3] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[6] ) , .A1 ( in[5] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( in[8] ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_4_ ( .A0 ( in[10] ) , .A1 ( in[9] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_5_ ( .A0 ( in[12] ) , .A1 ( in[11] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_6_ ( .A0 ( in[14] ) , .A1 ( in[13] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_7_ ( .A0 ( p0 ) , .A1 ( in[15] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_10_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_2_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_11_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_3_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_12_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_10_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_13_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_12_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_11_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_14_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l5_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_14_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_13_X[0] ) , .S ( sram[4] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_15_X[0] ) ) ;
endmodule


module mux_tree_tapbuf_size12_mem_3 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_8__59 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size12_mem_2 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_7__58 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size12_mem_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_6__57 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size12_mem_0 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_5__56 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size12_mem_5 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_4__55 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size12_mem_4 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_3__54 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size12_mem ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_2__53 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size12_mem_6 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_1__52 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_7_4 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size12_3 ( in , sram , sram_inv , out , p0 ) ;
input  [0:11] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_10_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_11_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

const1_7_4 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_11_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_3_ ( .A0 ( in[7] ) , .A1 ( in[6] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_4_ ( .A0 ( in[9] ) , .A1 ( in[8] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[10] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[11] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_10_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_10_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_11_X[0] ) ) ;
endmodule


module const1_6_5 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size12_2 ( in , sram , sram_inv , out , p0 ) ;
input  [0:11] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_10_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_11_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

const1_6_5 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_11_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_3_ ( .A0 ( in[7] ) , .A1 ( in[6] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_4_ ( .A0 ( in[9] ) , .A1 ( in[8] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[10] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[11] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_10_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_10_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_11_X[0] ) ) ;
endmodule


module const1_5_5 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size12_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:11] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_10_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_11_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

const1_5_5 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_11_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_3_ ( .A0 ( in[7] ) , .A1 ( in[6] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_4_ ( .A0 ( in[9] ) , .A1 ( in[8] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[10] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[11] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_10_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_10_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_11_X[0] ) ) ;
endmodule


module const1_4_5 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size12_0 ( in , sram , sram_inv , out , p0 ) ;
input  [0:11] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_10_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_11_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

const1_4_5 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_11_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_3_ ( .A0 ( in[7] ) , .A1 ( in[6] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_4_ ( .A0 ( in[9] ) , .A1 ( in[8] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[10] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[11] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_10_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_10_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_11_X[0] ) ) ;
endmodule


module const1_3_5 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size12_5 ( in , sram , sram_inv , out , p0 ) ;
input  [0:11] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_10_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_11_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

const1_3_5 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_11_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_3_ ( .A0 ( in[7] ) , .A1 ( in[6] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_4_ ( .A0 ( in[9] ) , .A1 ( in[8] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[10] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[11] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_10_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_10_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_11_X[0] ) ) ;
endmodule


module const1_2_5 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size12_4 ( in , sram , sram_inv , out , p0 ) ;
input  [0:11] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_10_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_11_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

const1_2_5 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_11_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_3_ ( .A0 ( in[7] ) , .A1 ( in[6] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_4_ ( .A0 ( in[9] ) , .A1 ( in[8] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[10] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[11] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_10_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_10_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_11_X[0] ) ) ;
endmodule


module const1_1_5 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size12 ( in , sram , sram_inv , out , p0 ) ;
input  [0:11] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_10_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_11_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

const1_1_5 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_11_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_3_ ( .A0 ( in[7] ) , .A1 ( in[6] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_4_ ( .A0 ( in[9] ) , .A1 ( in[8] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[10] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[11] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_10_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_10_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_11_X[0] ) ) ;
endmodule


module const1_0_5 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size12_6 ( in , sram , sram_inv , out , p0 ) ;
input  [0:11] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_10_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_11_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

const1_0_5 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_11_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_3_ ( .A0 ( in[7] ) , .A1 ( in[6] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_4_ ( .A0 ( in[9] ) , .A1 ( in[8] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[10] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[11] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_10_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_10_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_11_X[0] ) ) ;
endmodule


module sb_1__1_ ( prog_clk , chany_top_in , top_left_grid_pin_34_ , 
    top_left_grid_pin_35_ , top_left_grid_pin_36_ , top_left_grid_pin_37_ , 
    top_left_grid_pin_38_ , top_left_grid_pin_39_ , top_left_grid_pin_40_ , 
    top_left_grid_pin_41_ , chanx_right_in , right_top_grid_pin_42_ , 
    right_top_grid_pin_43_ , right_top_grid_pin_44_ , right_top_grid_pin_45_ , 
    right_top_grid_pin_46_ , right_top_grid_pin_47_ , right_top_grid_pin_48_ , 
    right_top_grid_pin_49_ , chany_bottom_in , bottom_left_grid_pin_34_ , 
    bottom_left_grid_pin_35_ , bottom_left_grid_pin_36_ , 
    bottom_left_grid_pin_37_ , bottom_left_grid_pin_38_ , 
    bottom_left_grid_pin_39_ , bottom_left_grid_pin_40_ , 
    bottom_left_grid_pin_41_ , chanx_left_in , left_top_grid_pin_42_ , 
    left_top_grid_pin_43_ , left_top_grid_pin_44_ , left_top_grid_pin_45_ , 
    left_top_grid_pin_46_ , left_top_grid_pin_47_ , left_top_grid_pin_48_ , 
    left_top_grid_pin_49_ , ccff_head , chany_top_out , chanx_right_out , 
    chany_bottom_out , chanx_left_out , ccff_tail ) ;
input  [0:0] prog_clk ;
input  [0:19] chany_top_in ;
input  [0:0] top_left_grid_pin_34_ ;
input  [0:0] top_left_grid_pin_35_ ;
input  [0:0] top_left_grid_pin_36_ ;
input  [0:0] top_left_grid_pin_37_ ;
input  [0:0] top_left_grid_pin_38_ ;
input  [0:0] top_left_grid_pin_39_ ;
input  [0:0] top_left_grid_pin_40_ ;
input  [0:0] top_left_grid_pin_41_ ;
input  [0:19] chanx_right_in ;
input  [0:0] right_top_grid_pin_42_ ;
input  [0:0] right_top_grid_pin_43_ ;
input  [0:0] right_top_grid_pin_44_ ;
input  [0:0] right_top_grid_pin_45_ ;
input  [0:0] right_top_grid_pin_46_ ;
input  [0:0] right_top_grid_pin_47_ ;
input  [0:0] right_top_grid_pin_48_ ;
input  [0:0] right_top_grid_pin_49_ ;
input  [0:19] chany_bottom_in ;
input  [0:0] bottom_left_grid_pin_34_ ;
input  [0:0] bottom_left_grid_pin_35_ ;
input  [0:0] bottom_left_grid_pin_36_ ;
input  [0:0] bottom_left_grid_pin_37_ ;
input  [0:0] bottom_left_grid_pin_38_ ;
input  [0:0] bottom_left_grid_pin_39_ ;
input  [0:0] bottom_left_grid_pin_40_ ;
input  [0:0] bottom_left_grid_pin_41_ ;
input  [0:19] chanx_left_in ;
input  [0:0] left_top_grid_pin_42_ ;
input  [0:0] left_top_grid_pin_43_ ;
input  [0:0] left_top_grid_pin_44_ ;
input  [0:0] left_top_grid_pin_45_ ;
input  [0:0] left_top_grid_pin_46_ ;
input  [0:0] left_top_grid_pin_47_ ;
input  [0:0] left_top_grid_pin_48_ ;
input  [0:0] left_top_grid_pin_49_ ;
input  [0:0] ccff_head ;
output [0:19] chany_top_out ;
output [0:19] chanx_right_out ;
output [0:19] chany_bottom_out ;
output [0:19] chanx_left_out ;
output [0:0] ccff_tail ;

wire [0:3] mux_tree_tapbuf_size10_0_sram ;
wire [0:3] mux_tree_tapbuf_size10_0_sram_inv ;
wire [0:3] mux_tree_tapbuf_size10_10_sram ;
wire [0:3] mux_tree_tapbuf_size10_10_sram_inv ;
wire [0:3] mux_tree_tapbuf_size10_11_sram ;
wire [0:3] mux_tree_tapbuf_size10_11_sram_inv ;
wire [0:3] mux_tree_tapbuf_size10_1_sram ;
wire [0:3] mux_tree_tapbuf_size10_1_sram_inv ;
wire [0:3] mux_tree_tapbuf_size10_2_sram ;
wire [0:3] mux_tree_tapbuf_size10_2_sram_inv ;
wire [0:3] mux_tree_tapbuf_size10_3_sram ;
wire [0:3] mux_tree_tapbuf_size10_3_sram_inv ;
wire [0:3] mux_tree_tapbuf_size10_4_sram ;
wire [0:3] mux_tree_tapbuf_size10_4_sram_inv ;
wire [0:3] mux_tree_tapbuf_size10_5_sram ;
wire [0:3] mux_tree_tapbuf_size10_5_sram_inv ;
wire [0:3] mux_tree_tapbuf_size10_6_sram ;
wire [0:3] mux_tree_tapbuf_size10_6_sram_inv ;
wire [0:3] mux_tree_tapbuf_size10_7_sram ;
wire [0:3] mux_tree_tapbuf_size10_7_sram_inv ;
wire [0:3] mux_tree_tapbuf_size10_8_sram ;
wire [0:3] mux_tree_tapbuf_size10_8_sram_inv ;
wire [0:3] mux_tree_tapbuf_size10_9_sram ;
wire [0:3] mux_tree_tapbuf_size10_9_sram_inv ;
wire [0:0] mux_tree_tapbuf_size10_mem_0_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size10_mem_10_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size10_mem_11_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size10_mem_1_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size10_mem_2_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size10_mem_3_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size10_mem_4_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size10_mem_5_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size10_mem_6_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size10_mem_7_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size10_mem_8_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size10_mem_9_ccff_tail ;
wire [0:3] mux_tree_tapbuf_size12_0_sram ;
wire [0:3] mux_tree_tapbuf_size12_0_sram_inv ;
wire [0:3] mux_tree_tapbuf_size12_1_sram ;
wire [0:3] mux_tree_tapbuf_size12_1_sram_inv ;
wire [0:3] mux_tree_tapbuf_size12_2_sram ;
wire [0:3] mux_tree_tapbuf_size12_2_sram_inv ;
wire [0:3] mux_tree_tapbuf_size12_3_sram ;
wire [0:3] mux_tree_tapbuf_size12_3_sram_inv ;
wire [0:3] mux_tree_tapbuf_size12_4_sram ;
wire [0:3] mux_tree_tapbuf_size12_4_sram_inv ;
wire [0:3] mux_tree_tapbuf_size12_5_sram ;
wire [0:3] mux_tree_tapbuf_size12_5_sram_inv ;
wire [0:3] mux_tree_tapbuf_size12_6_sram ;
wire [0:3] mux_tree_tapbuf_size12_6_sram_inv ;
wire [0:3] mux_tree_tapbuf_size12_7_sram ;
wire [0:3] mux_tree_tapbuf_size12_7_sram_inv ;
wire [0:0] mux_tree_tapbuf_size12_mem_0_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size12_mem_1_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size12_mem_2_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size12_mem_3_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size12_mem_4_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size12_mem_5_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size12_mem_6_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size12_mem_7_ccff_tail ;
wire [0:4] mux_tree_tapbuf_size16_0_sram ;
wire [0:4] mux_tree_tapbuf_size16_0_sram_inv ;
wire [0:4] mux_tree_tapbuf_size16_1_sram ;
wire [0:4] mux_tree_tapbuf_size16_1_sram_inv ;
wire [0:4] mux_tree_tapbuf_size16_2_sram ;
wire [0:4] mux_tree_tapbuf_size16_2_sram_inv ;
wire [0:4] mux_tree_tapbuf_size16_3_sram ;
wire [0:4] mux_tree_tapbuf_size16_3_sram_inv ;
wire [0:0] mux_tree_tapbuf_size16_mem_0_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size16_mem_1_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size16_mem_2_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size16_mem_3_ccff_tail ;
wire [0:2] mux_tree_tapbuf_size7_0_sram ;
wire [0:2] mux_tree_tapbuf_size7_0_sram_inv ;
wire [0:2] mux_tree_tapbuf_size7_1_sram ;
wire [0:2] mux_tree_tapbuf_size7_1_sram_inv ;
wire [0:2] mux_tree_tapbuf_size7_2_sram ;
wire [0:2] mux_tree_tapbuf_size7_2_sram_inv ;
wire [0:2] mux_tree_tapbuf_size7_3_sram ;
wire [0:2] mux_tree_tapbuf_size7_3_sram_inv ;
wire [0:0] mux_tree_tapbuf_size7_mem_0_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size7_mem_1_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size7_mem_2_ccff_tail ;

mux_tree_tapbuf_size12_6 mux_top_track_0 (
    .in ( { top_left_grid_pin_34_[0] , top_left_grid_pin_36_[0] , 
        top_left_grid_pin_38_[0] , top_left_grid_pin_40_[0] , 
        chanx_right_in[1] , chanx_right_in[2] , chanx_right_in[12] , 
        chany_bottom_in[2] , chany_bottom_in[12] , chanx_left_in[0] , 
        chanx_left_in[2] , chanx_left_in[12] } ) ,
    .sram ( mux_tree_tapbuf_size12_0_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size12_0_sram_inv ) , 
    .out ( chany_top_out[0] ) , .p0 ( optlc_net_127 ) ) ;
mux_tree_tapbuf_size12 mux_top_track_2 (
    .in ( { top_left_grid_pin_35_[0] , top_left_grid_pin_37_[0] , 
        top_left_grid_pin_39_[0] , top_left_grid_pin_41_[0] , 
        chanx_right_in[3] , chanx_right_in[4] , chanx_right_in[13] , 
        chany_bottom_in[4] , chany_bottom_in[13] , chanx_left_in[4] , 
        chanx_left_in[13] , chanx_left_in[19] } ) ,
    .sram ( mux_tree_tapbuf_size12_1_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size12_1_sram_inv ) , 
    .out ( chany_top_out[1] ) , .p0 ( optlc_net_125 ) ) ;
mux_tree_tapbuf_size12_4 mux_right_track_0 (
    .in ( { chany_top_in[2] , chany_top_in[12] , chany_top_in[19] , 
        right_top_grid_pin_42_[0] , right_top_grid_pin_44_[0] , 
        right_top_grid_pin_46_[0] , right_top_grid_pin_48_[0] , 
        chany_bottom_in[2] , chany_bottom_in[12] , chany_bottom_in[15] , 
        chanx_left_in[2] , chanx_left_in[12] } ) ,
    .sram ( mux_tree_tapbuf_size12_2_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size12_2_sram_inv ) , 
    .out ( chanx_right_out[0] ) , .p0 ( optlc_net_126 ) ) ;
mux_tree_tapbuf_size12_5 mux_right_track_2 (
    .in ( { chany_top_in[0] , chany_top_in[4] , chany_top_in[13] , 
        right_top_grid_pin_43_[0] , right_top_grid_pin_45_[0] , 
        right_top_grid_pin_47_[0] , right_top_grid_pin_49_[0] , 
        chany_bottom_in[4] , chany_bottom_in[11] , chany_bottom_in[13] , 
        chanx_left_in[4] , chanx_left_in[13] } ) ,
    .sram ( mux_tree_tapbuf_size12_3_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size12_3_sram_inv ) , 
    .out ( chanx_right_out[1] ) , .p0 ( optlc_net_126 ) ) ;
mux_tree_tapbuf_size12_0 mux_bottom_track_1 (
    .in ( { chany_top_in[2] , chany_top_in[12] , chanx_right_in[2] , 
        chanx_right_in[12] , chanx_right_in[15] , 
        bottom_left_grid_pin_34_[0] , bottom_left_grid_pin_36_[0] , 
        bottom_left_grid_pin_38_[0] , bottom_left_grid_pin_40_[0] , 
        chanx_left_in[1] , chanx_left_in[2] , chanx_left_in[12] } ) ,
    .sram ( mux_tree_tapbuf_size12_4_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size12_4_sram_inv ) , 
    .out ( chany_bottom_out[0] ) , .p0 ( optlc_net_126 ) ) ;
mux_tree_tapbuf_size12_1 mux_bottom_track_3 (
    .in ( { chany_top_in[4] , chany_top_in[13] , chanx_right_in[4] , 
        chanx_right_in[11] , chanx_right_in[13] , 
        bottom_left_grid_pin_35_[0] , bottom_left_grid_pin_37_[0] , 
        bottom_left_grid_pin_39_[0] , bottom_left_grid_pin_41_[0] , 
        chanx_left_in[3] , chanx_left_in[4] , chanx_left_in[13] } ) ,
    .sram ( mux_tree_tapbuf_size12_5_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size12_5_sram_inv ) , 
    .out ( chany_bottom_out[1] ) , .p0 ( optlc_net_125 ) ) ;
mux_tree_tapbuf_size12_2 mux_left_track_1 (
    .in ( { chany_top_in[0] , chany_top_in[2] , chany_top_in[12] , 
        chanx_right_in[2] , chanx_right_in[12] , chany_bottom_in[2] , 
        chany_bottom_in[12] , chany_bottom_in[19] , left_top_grid_pin_42_[0] , 
        left_top_grid_pin_44_[0] , left_top_grid_pin_46_[0] , 
        left_top_grid_pin_48_[0] } ) ,
    .sram ( mux_tree_tapbuf_size12_6_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size12_6_sram_inv ) , 
    .out ( chanx_left_out[0] ) , .p0 ( optlc_net_127 ) ) ;
mux_tree_tapbuf_size12_3 mux_left_track_3 (
    .in ( { chany_top_in[4] , chany_top_in[13] , chany_top_in[19] , 
        chanx_right_in[4] , chanx_right_in[13] , chany_bottom_in[0] , 
        chany_bottom_in[4] , chany_bottom_in[13] , left_top_grid_pin_43_[0] , 
        left_top_grid_pin_45_[0] , left_top_grid_pin_47_[0] , 
        left_top_grid_pin_49_[0] } ) ,
    .sram ( mux_tree_tapbuf_size12_7_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size12_7_sram_inv ) , 
    .out ( chanx_left_out[1] ) , .p0 ( optlc_net_127 ) ) ;
mux_tree_tapbuf_size12_mem_6 mem_top_track_0 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( ccff_head ) , 
    .ccff_tail ( mux_tree_tapbuf_size12_mem_0_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size12_0_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size12_0_sram_inv ) ) ;
mux_tree_tapbuf_size12_mem mem_top_track_2 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size12_mem_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size12_mem_1_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size12_1_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size12_1_sram_inv ) ) ;
mux_tree_tapbuf_size12_mem_4 mem_right_track_0 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size7_mem_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size12_mem_2_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size12_2_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size12_2_sram_inv ) ) ;
mux_tree_tapbuf_size12_mem_5 mem_right_track_2 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size12_mem_2_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size12_mem_3_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size12_3_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size12_3_sram_inv ) ) ;
mux_tree_tapbuf_size12_mem_0 mem_bottom_track_1 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size7_mem_1_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size12_mem_4_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size12_4_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size12_4_sram_inv ) ) ;
mux_tree_tapbuf_size12_mem_1 mem_bottom_track_3 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size12_mem_4_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size12_mem_5_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size12_5_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size12_5_sram_inv ) ) ;
mux_tree_tapbuf_size12_mem_2 mem_left_track_1 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size7_mem_2_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size12_mem_6_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size12_6_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size12_6_sram_inv ) ) ;
mux_tree_tapbuf_size12_mem_3 mem_left_track_3 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size12_mem_6_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size12_mem_7_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size12_7_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size12_7_sram_inv ) ) ;
mux_tree_tapbuf_size16 mux_top_track_4 (
    .in ( { top_left_grid_pin_34_[0] , top_left_grid_pin_35_[0] , 
        top_left_grid_pin_36_[0] , top_left_grid_pin_37_[0] , 
        top_left_grid_pin_38_[0] , top_left_grid_pin_39_[0] , 
        top_left_grid_pin_40_[0] , top_left_grid_pin_41_[0] , 
        chanx_right_in[5] , chanx_right_in[7] , chanx_right_in[14] , 
        chany_bottom_in[5] , chany_bottom_in[14] , chanx_left_in[5] , 
        chanx_left_in[14] , chanx_left_in[15] } ) ,
    .sram ( mux_tree_tapbuf_size16_0_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size16_0_sram_inv ) , 
    .out ( chany_top_out[2] ) , .p0 ( optlc_net_125 ) ) ;
mux_tree_tapbuf_size16_2 mux_right_track_4 (
    .in ( { chany_top_in[1] , chany_top_in[5] , chany_top_in[14] , 
        right_top_grid_pin_42_[0] , right_top_grid_pin_43_[0] , 
        right_top_grid_pin_44_[0] , right_top_grid_pin_45_[0] , 
        right_top_grid_pin_46_[0] , right_top_grid_pin_47_[0] , 
        right_top_grid_pin_48_[0] , right_top_grid_pin_49_[0] , 
        chany_bottom_in[5] , chany_bottom_in[7] , chany_bottom_in[14] , 
        chanx_left_in[5] , chanx_left_in[14] } ) ,
    .sram ( mux_tree_tapbuf_size16_1_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size16_1_sram_inv ) , 
    .out ( chanx_right_out[2] ) , .p0 ( optlc_net_128 ) ) ;
mux_tree_tapbuf_size16_0 mux_bottom_track_5 (
    .in ( { chany_top_in[5] , chany_top_in[14] , chanx_right_in[5] , 
        chanx_right_in[7] , chanx_right_in[14] , bottom_left_grid_pin_34_[0] , 
        bottom_left_grid_pin_35_[0] , bottom_left_grid_pin_36_[0] , 
        bottom_left_grid_pin_37_[0] , bottom_left_grid_pin_38_[0] , 
        bottom_left_grid_pin_39_[0] , bottom_left_grid_pin_40_[0] , 
        bottom_left_grid_pin_41_[0] , chanx_left_in[5] , chanx_left_in[7] , 
        chanx_left_in[14] } ) ,
    .sram ( mux_tree_tapbuf_size16_2_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size16_2_sram_inv ) , 
    .out ( chany_bottom_out[2] ) , .p0 ( optlc_net_125 ) ) ;
mux_tree_tapbuf_size16_1 mux_left_track_5 (
    .in ( { chany_top_in[5] , chany_top_in[14] , chany_top_in[15] , 
        chanx_right_in[5] , chanx_right_in[14] , chany_bottom_in[1] , 
        chany_bottom_in[5] , chany_bottom_in[14] , left_top_grid_pin_42_[0] , 
        left_top_grid_pin_43_[0] , left_top_grid_pin_44_[0] , 
        left_top_grid_pin_45_[0] , left_top_grid_pin_46_[0] , 
        left_top_grid_pin_47_[0] , left_top_grid_pin_48_[0] , 
        left_top_grid_pin_49_[0] } ) ,
    .sram ( mux_tree_tapbuf_size16_3_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size16_3_sram_inv ) , 
    .out ( chanx_left_out[2] ) , .p0 ( optlc_net_127 ) ) ;
mux_tree_tapbuf_size16_mem mem_top_track_4 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size12_mem_1_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size16_mem_0_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size16_0_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size16_0_sram_inv ) ) ;
mux_tree_tapbuf_size16_mem_2 mem_right_track_4 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size12_mem_3_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size16_mem_1_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size16_1_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size16_1_sram_inv ) ) ;
mux_tree_tapbuf_size16_mem_0 mem_bottom_track_5 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size12_mem_5_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size16_mem_2_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size16_2_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size16_2_sram_inv ) ) ;
mux_tree_tapbuf_size16_mem_1 mem_left_track_5 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size12_mem_7_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size16_mem_3_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size16_3_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size16_3_sram_inv ) ) ;
mux_tree_tapbuf_size10_1 mux_top_track_8 (
    .in ( { top_left_grid_pin_34_[0] , top_left_grid_pin_38_[0] , 
        chanx_right_in[6] , chanx_right_in[11] , chanx_right_in[16] , 
        chany_bottom_in[6] , chany_bottom_in[16] , chanx_left_in[6] , 
        chanx_left_in[11] , chanx_left_in[16] } ) ,
    .sram ( mux_tree_tapbuf_size10_0_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size10_0_sram_inv ) , 
    .out ( chany_top_out[4] ) , .p0 ( optlc_net_129 ) ) ;
mux_tree_tapbuf_size10_9 mux_top_track_16 (
    .in ( { top_left_grid_pin_35_[0] , top_left_grid_pin_39_[0] , 
        chanx_right_in[8] , chanx_right_in[15] , chanx_right_in[17] , 
        chany_bottom_in[8] , chany_bottom_in[17] , chanx_left_in[7] , 
        chanx_left_in[8] , chanx_left_in[17] } ) ,
    .sram ( mux_tree_tapbuf_size10_1_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size10_1_sram_inv ) , 
    .out ( chany_top_out[8] ) , .p0 ( optlc_net_129 ) ) ;
mux_tree_tapbuf_size10_10 mux_top_track_24 (
    .in ( { top_left_grid_pin_36_[0] , top_left_grid_pin_40_[0] , 
        chanx_right_in[9] , chanx_right_in[18] , chanx_right_in[19] , 
        chany_bottom_in[9] , chany_bottom_in[18] , chanx_left_in[3] , 
        chanx_left_in[9] , chanx_left_in[18] } ) ,
    .sram ( mux_tree_tapbuf_size10_2_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size10_2_sram_inv ) , 
    .out ( chany_top_out[12] ) , .p0 ( optlc_net_129 ) ) ;
mux_tree_tapbuf_size10_8 mux_right_track_8 (
    .in ( { chany_top_in[3] , chany_top_in[6] , chany_top_in[16] , 
        right_top_grid_pin_42_[0] , right_top_grid_pin_46_[0] , 
        chany_bottom_in[3] , chany_bottom_in[6] , chany_bottom_in[16] , 
        chanx_left_in[6] , chanx_left_in[16] } ) ,
    .sram ( mux_tree_tapbuf_size10_3_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size10_3_sram_inv ) , 
    .out ( chanx_right_out[4] ) , .p0 ( optlc_net_128 ) ) ;
mux_tree_tapbuf_size10_6 mux_right_track_16 (
    .in ( { chany_top_in[7] , chany_top_in[8] , chany_top_in[17] , 
        right_top_grid_pin_43_[0] , right_top_grid_pin_47_[0] , 
        chany_bottom_in[1] , chany_bottom_in[8] , chany_bottom_in[17] , 
        chanx_left_in[8] , chanx_left_in[17] } ) ,
    .sram ( mux_tree_tapbuf_size10_4_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size10_4_sram_inv ) , 
    .out ( chanx_right_out[8] ) , .p0 ( optlc_net_128 ) ) ;
mux_tree_tapbuf_size10_7 mux_right_track_24 (
    .in ( { chany_top_in[9] , chany_top_in[11] , chany_top_in[18] , 
        right_top_grid_pin_44_[0] , right_top_grid_pin_48_[0] , 
        chany_bottom_in[0] , chany_bottom_in[9] , chany_bottom_in[18] , 
        chanx_left_in[9] , chanx_left_in[18] } ) ,
    .sram ( mux_tree_tapbuf_size10_5_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size10_5_sram_inv ) , 
    .out ( chanx_right_out[12] ) , .p0 ( optlc_net_128 ) ) ;
mux_tree_tapbuf_size10_2 mux_bottom_track_9 (
    .in ( { chany_top_in[6] , chany_top_in[16] , chanx_right_in[3] , 
        chanx_right_in[6] , chanx_right_in[16] , bottom_left_grid_pin_34_[0] , 
        bottom_left_grid_pin_38_[0] , chanx_left_in[6] , chanx_left_in[11] , 
        chanx_left_in[16] } ) ,
    .sram ( mux_tree_tapbuf_size10_6_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size10_6_sram_inv ) , 
    .out ( chany_bottom_out[4] ) , .p0 ( optlc_net_127 ) ) ;
mux_tree_tapbuf_size10_0 mux_bottom_track_17 (
    .in ( { chany_top_in[8] , chany_top_in[17] , chanx_right_in[1] , 
        chanx_right_in[8] , chanx_right_in[17] , bottom_left_grid_pin_35_[0] , 
        bottom_left_grid_pin_39_[0] , chanx_left_in[8] , chanx_left_in[15] , 
        chanx_left_in[17] } ) ,
    .sram ( mux_tree_tapbuf_size10_7_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size10_7_sram_inv ) , 
    .out ( chany_bottom_out[8] ) , .p0 ( optlc_net_126 ) ) ;
mux_tree_tapbuf_size10_1 mux_bottom_track_25 (
    .in ( { chany_top_in[9] , chany_top_in[18] , chanx_right_in[0] , 
        chanx_right_in[9] , chanx_right_in[18] , bottom_left_grid_pin_36_[0] , 
        bottom_left_grid_pin_40_[0] , chanx_left_in[9] , chanx_left_in[18] , 
        chanx_left_in[19] } ) ,
    .sram ( mux_tree_tapbuf_size10_8_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size10_8_sram_inv ) , 
    .out ( chany_bottom_out[12] ) , .p0 ( optlc_net_126 ) ) ;
mux_tree_tapbuf_size10_5 mux_left_track_9 (
    .in ( { chany_top_in[6] , chany_top_in[11] , chany_top_in[16] , 
        chanx_right_in[6] , chanx_right_in[16] , chany_bottom_in[3] , 
        chany_bottom_in[6] , chany_bottom_in[16] , left_top_grid_pin_42_[0] , 
        left_top_grid_pin_46_[0] } ) ,
    .sram ( mux_tree_tapbuf_size10_9_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size10_9_sram_inv ) , 
    .out ( chanx_left_out[4] ) , .p0 ( optlc_net_129 ) ) ;
mux_tree_tapbuf_size10_3 mux_left_track_17 (
    .in ( { chany_top_in[7] , chany_top_in[8] , chany_top_in[17] , 
        chanx_right_in[8] , chanx_right_in[17] , chany_bottom_in[7] , 
        chany_bottom_in[8] , chany_bottom_in[17] , left_top_grid_pin_43_[0] , 
        left_top_grid_pin_47_[0] } ) ,
    .sram ( mux_tree_tapbuf_size10_10_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size10_10_sram_inv ) , 
    .out ( chanx_left_out[8] ) , .p0 ( optlc_net_129 ) ) ;
mux_tree_tapbuf_size10_4 mux_left_track_25 (
    .in ( { chany_top_in[3] , chany_top_in[9] , chany_top_in[18] , 
        chanx_right_in[9] , chanx_right_in[18] , chany_bottom_in[9] , 
        chany_bottom_in[11] , chany_bottom_in[18] , left_top_grid_pin_44_[0] , 
        left_top_grid_pin_48_[0] } ) ,
    .sram ( mux_tree_tapbuf_size10_11_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size10_11_sram_inv ) , 
    .out ( chanx_left_out[12] ) , .p0 ( optlc_net_129 ) ) ;
mux_tree_tapbuf_size10_mem_1 mem_top_track_8 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size16_mem_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size10_mem_0_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size10_0_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size10_0_sram_inv ) ) ;
mux_tree_tapbuf_size10_mem_9 mem_top_track_16 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size10_mem_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size10_mem_1_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size10_1_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size10_1_sram_inv ) ) ;
mux_tree_tapbuf_size10_mem_10 mem_top_track_24 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size10_mem_1_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size10_mem_2_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size10_2_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size10_2_sram_inv ) ) ;
mux_tree_tapbuf_size10_mem_8 mem_right_track_8 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size16_mem_1_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size10_mem_3_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size10_3_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size10_3_sram_inv ) ) ;
mux_tree_tapbuf_size10_mem_6 mem_right_track_16 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size10_mem_3_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size10_mem_4_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size10_4_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size10_4_sram_inv ) ) ;
mux_tree_tapbuf_size10_mem_7 mem_right_track_24 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size10_mem_4_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size10_mem_5_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size10_5_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size10_5_sram_inv ) ) ;
mux_tree_tapbuf_size10_mem_2 mem_bottom_track_9 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size16_mem_2_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size10_mem_6_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size10_6_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size10_6_sram_inv ) ) ;
mux_tree_tapbuf_size10_mem_0 mem_bottom_track_17 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size10_mem_6_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size10_mem_7_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size10_7_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size10_7_sram_inv ) ) ;
mux_tree_tapbuf_size10_mem_1 mem_bottom_track_25 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size10_mem_7_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size10_mem_8_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size10_8_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size10_8_sram_inv ) ) ;
mux_tree_tapbuf_size10_mem_5 mem_left_track_9 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size16_mem_3_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size10_mem_9_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size10_9_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size10_9_sram_inv ) ) ;
mux_tree_tapbuf_size10_mem_3 mem_left_track_17 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size10_mem_9_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size10_mem_10_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size10_10_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size10_10_sram_inv ) ) ;
mux_tree_tapbuf_size10_mem_4 mem_left_track_25 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size10_mem_10_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size10_mem_11_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size10_11_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size10_11_sram_inv ) ) ;
mux_tree_tapbuf_size7_6 mux_top_track_32 (
    .in ( { top_left_grid_pin_37_[0] , top_left_grid_pin_41_[0] , 
        chanx_right_in[0] , chanx_right_in[10] , chany_bottom_in[10] , 
        chanx_left_in[1] , chanx_left_in[10] } ) ,
    .sram ( mux_tree_tapbuf_size7_0_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size7_0_sram_inv ) , 
    .out ( chany_top_out[16] ) , .p0 ( optlc_net_126 ) ) ;
mux_tree_tapbuf_size7_2_1 mux_right_track_32 (
    .in ( { chany_top_in[10] , chany_top_in[15] , right_top_grid_pin_45_[0] , 
        right_top_grid_pin_49_[0] , chany_bottom_in[10] , 
        chany_bottom_in[19] , chanx_left_in[10] } ) ,
    .sram ( mux_tree_tapbuf_size7_1_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size7_1_sram_inv ) , 
    .out ( chanx_right_out[16] ) , .p0 ( optlc_net_126 ) ) ;
mux_tree_tapbuf_size7_0_2 mux_bottom_track_33 (
    .in ( { chany_top_in[10] , chanx_right_in[10] , chanx_right_in[19] , 
        bottom_left_grid_pin_37_[0] , bottom_left_grid_pin_41_[0] , 
        chanx_left_in[0] , chanx_left_in[10] } ) ,
    .sram ( mux_tree_tapbuf_size7_2_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size7_2_sram_inv ) , 
    .out ( chany_bottom_out[16] ) , .p0 ( optlc_net_126 ) ) ;
mux_tree_tapbuf_size7_1_2 mux_left_track_33 (
    .in ( { chany_top_in[1] , chany_top_in[10] , chanx_right_in[10] , 
        chany_bottom_in[10] , chany_bottom_in[15] , left_top_grid_pin_45_[0] , 
        left_top_grid_pin_49_[0] } ) ,
    .sram ( mux_tree_tapbuf_size7_3_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size7_3_sram_inv ) , 
    .out ( chanx_left_out[16] ) , .p0 ( optlc_net_127 ) ) ;
mux_tree_tapbuf_size7_mem_6 mem_top_track_32 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size10_mem_2_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size7_mem_0_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size7_0_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size7_0_sram_inv ) ) ;
mux_tree_tapbuf_size7_mem_2_1 mem_right_track_32 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size10_mem_5_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size7_mem_1_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size7_1_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size7_1_sram_inv ) ) ;
mux_tree_tapbuf_size7_mem_0_2 mem_bottom_track_33 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size10_mem_8_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size7_mem_2_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size7_2_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size7_2_sram_inv ) ) ;
mux_tree_tapbuf_size7_mem_1_2 mem_left_track_33 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size10_mem_11_ccff_tail ) ,
    .ccff_tail ( { ropt_net_135 } ) ,
    .mem_out ( mux_tree_tapbuf_size7_3_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size7_3_sram_inv ) ) ;
sky130_fd_sc_hd__conb_1 optlc_121 ( .LO ( SYNOPSYS_UNCONNECTED_1 ) , 
    .HI ( optlc_net_125 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_2__1 ( .A ( chany_top_in[4] ) , 
    .X ( chany_bottom_out[5] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_3__2 ( .A ( chany_top_in[5] ) , 
    .X ( chany_bottom_out[6] ) ) ;
sky130_fd_sc_hd__conb_1 optlc_124 ( .LO ( SYNOPSYS_UNCONNECTED_2 ) , 
    .HI ( optlc_net_126 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_126 ( .LO ( SYNOPSYS_UNCONNECTED_3 ) , 
    .HI ( optlc_net_127 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_6__5 ( .A ( chany_top_in[9] ) , 
    .X ( chany_bottom_out[10] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_7__6 ( .A ( chany_top_in[10] ) , 
    .X ( ropt_net_139 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_8__7 ( .A ( chany_top_in[12] ) , 
    .X ( chany_bottom_out[13] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_9__8 ( .A ( chany_top_in[13] ) , 
    .X ( chany_bottom_out[14] ) ) ;
sky130_fd_sc_hd__conb_1 optlc_128 ( .LO ( SYNOPSYS_UNCONNECTED_4 ) , 
    .HI ( optlc_net_128 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_11__10 ( .A ( chany_top_in[16] ) , 
    .X ( chany_bottom_out[17] ) ) ;
sky130_fd_sc_hd__conb_1 optlc_130 ( .LO ( SYNOPSYS_UNCONNECTED_5 ) , 
    .HI ( optlc_net_129 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_13__12 ( .A ( chany_top_in[18] ) , 
    .X ( chany_bottom_out[19] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_737 ( .A ( ropt_net_131 ) , 
    .X ( chany_top_out[5] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_738 ( .A ( chany_top_in[8] ) , 
    .X ( chany_bottom_out[9] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_739 ( .A ( chanx_right_in[8] ) , 
    .X ( chanx_left_out[9] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_17__16 ( .A ( chanx_right_in[6] ) , 
    .X ( chanx_left_out[7] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_749 ( .A ( ropt_net_138 ) , 
    .X ( chanx_right_out[10] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_19__18 ( .A ( chanx_right_in[9] ) , 
    .X ( chanx_left_out[10] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_20__19 ( .A ( chanx_right_in[10] ) , 
    .X ( aps_rename_1_ ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_21__20 ( .A ( chanx_right_in[12] ) , 
    .X ( aps_rename_2_ ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_22__21 ( .A ( chanx_right_in[13] ) , 
    .X ( chanx_left_out[14] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_23__22 ( .A ( chanx_right_in[14] ) , 
    .X ( chanx_left_out[15] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_24__23 ( .A ( chanx_right_in[16] ) , 
    .X ( chanx_left_out[17] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_25__24 ( .A ( chanx_right_in[17] ) , 
    .X ( chanx_left_out[18] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_740 ( 
    .A ( chany_bottom_in[17] ) , .X ( chany_top_out[18] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_27__26 ( .A ( chany_bottom_in[2] ) , 
    .X ( chany_top_out[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd1_1 FTB_28__27 ( .A ( chany_bottom_in[4] ) , 
    .X ( ropt_net_131 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_744 ( .A ( ropt_net_135 ) , 
    .X ( ccff_tail[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd1_1 FTB_30__29 ( .A ( chany_bottom_in[6] ) , 
    .X ( chany_top_out[7] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_31__30 ( .A ( chany_bottom_in[8] ) , 
    .X ( chany_top_out[9] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_745 ( .A ( ropt_net_136 ) , 
    .X ( ropt_net_138 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_33__32 ( .A ( chany_bottom_in[10] ) , 
    .X ( chany_top_out[11] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_34__33 ( .A ( chany_bottom_in[12] ) , 
    .X ( chany_top_out[13] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_746 ( .A ( ropt_net_137 ) , 
    .X ( chanx_right_out[13] ) ) ;
sky130_fd_sc_hd__dlygate4sd1_1 FTB_36__35 ( .A ( chany_bottom_in[14] ) , 
    .X ( chany_top_out[15] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_37__36 ( .A ( chany_bottom_in[16] ) , 
    .X ( chany_top_out[17] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_763 ( .A ( ropt_net_139 ) , 
    .X ( chany_bottom_out[11] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_42__41 ( .A ( chanx_left_in[5] ) , 
    .X ( chanx_right_out[6] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_44__43 ( .A ( chanx_left_in[8] ) , 
    .X ( chanx_right_out[9] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_45__44 ( .A ( chanx_left_in[9] ) , 
    .X ( ropt_net_136 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_50__49 ( .A ( chanx_left_in[16] ) , 
    .X ( chanx_right_out[17] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_52__51 ( .A ( chanx_left_in[18] ) , 
    .X ( chanx_right_out[19] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_RR_84 ( .A ( chanx_right_in[4] ) , 
    .X ( chanx_left_out[5] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_RR_89 ( .A ( chanx_left_in[13] ) , 
    .X ( chanx_right_out[14] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_RR_90 ( .A ( chanx_left_in[17] ) , 
    .X ( chanx_right_out[18] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_RR_93 ( .A ( chanx_right_in[2] ) , 
    .X ( chanx_left_out[3] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_RR_94 ( .A ( chanx_right_in[5] ) , 
    .X ( chanx_left_out[6] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_RR_95 ( .A ( chany_bottom_in[9] ) , 
    .X ( chany_top_out[10] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_RR_96 ( .A ( chanx_left_in[6] ) , 
    .X ( chanx_right_out[7] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_RR_97 ( .A ( chanx_left_in[12] ) , 
    .X ( ropt_net_137 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_RR_98 ( .A ( chanx_left_in[14] ) , 
    .X ( chanx_right_out[15] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 BUFT_RR_100 ( .A ( aps_rename_2_ ) , 
    .X ( chanx_left_out[13] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_RR_101 ( .A ( chanx_left_in[2] ) , 
    .X ( chanx_right_out[3] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_RR_102 ( .A ( chanx_left_in[4] ) , 
    .X ( chanx_right_out[5] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_P_107 ( .A ( chany_top_in[2] ) , 
    .X ( chany_bottom_out[3] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_P_108 ( .A ( chany_top_in[6] ) , 
    .X ( chany_bottom_out[7] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_P_109 ( .A ( chany_top_in[14] ) , 
    .X ( chany_bottom_out[15] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_P_110 ( .A ( chany_top_in[17] ) , 
    .X ( chany_bottom_out[18] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_P_111 ( .A ( chanx_right_in[18] ) , 
    .X ( chanx_left_out[19] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_P_112 ( .A ( chany_bottom_in[5] ) , 
    .X ( chany_top_out[6] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_P_113 ( .A ( chany_bottom_in[13] ) , 
    .X ( chany_top_out[14] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_P_114 ( .A ( chany_bottom_in[18] ) , 
    .X ( chany_top_out[19] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_P_115 ( .A ( chanx_left_in[10] ) , 
    .X ( chanx_right_out[11] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 BUFT_P_117 ( .A ( aps_rename_1_ ) , 
    .X ( chanx_left_out[11] ) ) ;
endmodule


module mux_tree_tapbuf_size10_mem ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_33__59 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_34 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size10 ( in , sram , sram_inv , out , p0 ) ;
input  [0:9] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

const1_34 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[6] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[8] ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[9] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
endmodule


module mux_tree_tapbuf_size6_mem_0_2 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd1_1 FTB_32__58 ( .A ( mem_out[2] ) , 
    .X ( net_net_93 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 BUFT_RR_93 ( .A ( net_net_93 ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size6_mem_6 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_31__57 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_31 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size6_0_2 ( in , sram , sram_inv , out , p0 ) ;
input  [0:5] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;

const1_31 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
endmodule


module const1_30_1 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size6_6 ( in , sram , sram_inv , out , p0 ) ;
input  [0:5] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;

const1_30_1 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
endmodule


module mux_tree_tapbuf_size14_mem_0 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_30__56 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size14_mem ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_29__55 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_29_1 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size14_0 ( in , sram , sram_inv , out , p0 ) ;
input  [0:13] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_10_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_11_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_12_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_13_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

const1_29_1 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_13_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_3_ ( .A0 ( in[7] ) , .A1 ( in[6] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_4_ ( .A0 ( in[9] ) , .A1 ( in[8] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_5_ ( .A0 ( in[11] ) , .A1 ( in[10] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_6_ ( .A0 ( in[13] ) , .A1 ( in[12] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_10_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_11_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_10_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_12_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_12_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_11_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_13_X[0] ) ) ;
endmodule


module const1_28_1 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size14 ( in , sram , sram_inv , out , p0 ) ;
input  [0:13] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_10_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_11_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_12_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_13_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

const1_28_1 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_13_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_3_ ( .A0 ( in[7] ) , .A1 ( in[6] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_4_ ( .A0 ( in[9] ) , .A1 ( in[8] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_5_ ( .A0 ( in[11] ) , .A1 ( in[10] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_6_ ( .A0 ( in[13] ) , .A1 ( in[12] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_10_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_11_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_10_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_12_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_12_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_11_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_13_X[0] ) ) ;
endmodule


module mux_tree_tapbuf_size9_mem ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_28__54 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size9_mem_0 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_27__53 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_27_1 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size9 ( in , sram , sram_inv , out , p0 ) ;
input  [0:8] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;

const1_27_1 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[7] ) , .A1 ( in[6] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[8] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
endmodule


module const1_26_2 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size9_0 ( in , sram , sram_inv , out , p0 ) ;
input  [0:8] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;

const1_26_2 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[7] ) , .A1 ( in[6] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[8] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_13 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_26__52 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_3_2 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_25__51 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_2_2 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_24__50 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_1_2 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_23__49 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_0_2 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_22__48 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_25_2 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_13 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_25_2 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
endmodule


module const1_24_2 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_3_2 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_24_2 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
endmodule


module const1_23_2 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_2_2 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_23_2 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
endmodule


module const1_22_2 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_1_2 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_22_2 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
endmodule


module const1_21_2 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_0_2 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_21_2 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_62 ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
endmodule


module mux_tree_tapbuf_size3_mem_7 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_21__47 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size3_mem_6 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_20__46 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size3_mem_5 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_19__45 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size3_mem_4 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_18__44 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size3_mem_3_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_17__43 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size3_mem_2_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_16__42 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size3_mem_1_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_15__41 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size3_mem_0_2 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_14__40 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_20_2 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size3_7 ( in , sram , sram_inv , out , p0 ) ;
input  [0:2] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;

const1_20_2 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( p0 ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
endmodule


module const1_19_2 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size3_6 ( in , sram , sram_inv , out , p0 ) ;
input  [0:2] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;

const1_19_2 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( p0 ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
endmodule


module const1_18_2 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size3_5 ( in , sram , sram_inv , out , p0 ) ;
input  [0:2] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;

const1_18_2 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( p0 ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
endmodule


module const1_17_2 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size3_4 ( in , sram , sram_inv , out , p0 ) ;
input  [0:2] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;

const1_17_2 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( p0 ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
endmodule


module const1_16_3 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size3_3_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:2] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;

const1_16_3 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( p0 ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
endmodule


module const1_15_3 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size3_2_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:2] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;

const1_15_3 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( p0 ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
endmodule


module const1_14_3 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size3_1_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:2] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;

const1_14_3 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( p0 ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
endmodule


module const1_13_3 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size3_0_2 ( in , sram , sram_inv , out , p0 ) ;
input  [0:2] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;

const1_13_3 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( p0 ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
endmodule


module mux_tree_tapbuf_size4_mem_0_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_13__39 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size4_mem_6 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_12__38 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_12_3 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size4_0_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:3] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;

const1_12_3 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( in[2] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , .A1 ( in[3] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
endmodule


module const1_11_3 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size4_6 ( in , sram , sram_inv , out , p0 ) ;
input  [0:3] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;

const1_11_3 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( in[2] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , .A1 ( in[3] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
endmodule


module mux_tree_tapbuf_size7_mem_1_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_11__37 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size7_mem_0_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_10__36 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size7_mem_3 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_9__35 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size7_mem_2 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_8__34 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size7_mem_2 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_7__33 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size7_mem_5 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_6__32 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size7_mem_4 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_5__31 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_10_3 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size7_1_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:6] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;

const1_10_3 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_3_ ( .A0 ( p0 ) , .A1 ( in[6] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
endmodule


module const1_9_3 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size7_0_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:6] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;

const1_9_3 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_3_ ( .A0 ( p0 ) , .A1 ( in[6] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
endmodule


module const1_8_3 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size7_3 ( in , sram , sram_inv , out , p0 ) ;
input  [0:6] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;

const1_8_3 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_3_ ( .A0 ( p0 ) , .A1 ( in[6] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
endmodule


module const1_7_3 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size7_2 ( in , sram , sram_inv , out , p0 ) ;
input  [0:6] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;

const1_7_3 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_3_ ( .A0 ( p0 ) , .A1 ( in[6] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
endmodule


module const1_6_4 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size7_2 ( in , sram , sram_inv , out , p0 ) ;
input  [0:6] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;

const1_6_4 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_3_ ( .A0 ( p0 ) , .A1 ( in[6] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
endmodule


module const1_5_4 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size7_5 ( in , sram , sram_inv , out , p0 ) ;
input  [0:6] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;

const1_5_4 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_3_ ( .A0 ( p0 ) , .A1 ( in[6] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
endmodule


module const1_4_4 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size7_4 ( in , sram , sram_inv , out , p0 ) ;
input  [0:6] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;

const1_4_4 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_3_ ( .A0 ( p0 ) , .A1 ( in[6] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
endmodule


module mux_tree_tapbuf_size8_mem_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_4__30 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size8_mem_0 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_3__29 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size8_mem_2 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_2__28 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size8_mem ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_1__27 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_3_4 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size8_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:7] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;

const1_3_4 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( in[2] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[4] ) , .A1 ( in[3] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[6] ) , .A1 ( in[5] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
endmodule


module const1_2_4 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size8_0 ( in , sram , sram_inv , out , p0 ) ;
input  [0:7] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;

const1_2_4 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( in[2] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[4] ) , .A1 ( in[3] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[6] ) , .A1 ( in[5] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
endmodule


module const1_1_4 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size8_2 ( in , sram , sram_inv , out , p0 ) ;
input  [0:7] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;

const1_1_4 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( in[2] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[4] ) , .A1 ( in[3] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[6] ) , .A1 ( in[5] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
endmodule


module const1_0_4 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size8 ( in , sram , sram_inv , out , p0 ) ;
input  [0:7] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;

const1_0_4 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( in[2] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[4] ) , .A1 ( in[3] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[6] ) , .A1 ( in[5] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
endmodule


module sb_1__0_ ( prog_clk , chany_top_in , top_left_grid_pin_34_ , 
    top_left_grid_pin_35_ , top_left_grid_pin_36_ , top_left_grid_pin_37_ , 
    top_left_grid_pin_38_ , top_left_grid_pin_39_ , top_left_grid_pin_40_ , 
    top_left_grid_pin_41_ , chanx_right_in , right_top_grid_pin_42_ , 
    right_top_grid_pin_43_ , right_top_grid_pin_44_ , right_top_grid_pin_45_ , 
    right_top_grid_pin_46_ , right_top_grid_pin_47_ , right_top_grid_pin_48_ , 
    right_top_grid_pin_49_ , right_bottom_grid_pin_1_ , chanx_left_in , 
    left_top_grid_pin_42_ , left_top_grid_pin_43_ , left_top_grid_pin_44_ , 
    left_top_grid_pin_45_ , left_top_grid_pin_46_ , left_top_grid_pin_47_ , 
    left_top_grid_pin_48_ , left_top_grid_pin_49_ , left_bottom_grid_pin_1_ , 
    ccff_head , chany_top_out , chanx_right_out , chanx_left_out , ccff_tail ) ;
input  [0:0] prog_clk ;
input  [0:19] chany_top_in ;
input  [0:0] top_left_grid_pin_34_ ;
input  [0:0] top_left_grid_pin_35_ ;
input  [0:0] top_left_grid_pin_36_ ;
input  [0:0] top_left_grid_pin_37_ ;
input  [0:0] top_left_grid_pin_38_ ;
input  [0:0] top_left_grid_pin_39_ ;
input  [0:0] top_left_grid_pin_40_ ;
input  [0:0] top_left_grid_pin_41_ ;
input  [0:19] chanx_right_in ;
input  [0:0] right_top_grid_pin_42_ ;
input  [0:0] right_top_grid_pin_43_ ;
input  [0:0] right_top_grid_pin_44_ ;
input  [0:0] right_top_grid_pin_45_ ;
input  [0:0] right_top_grid_pin_46_ ;
input  [0:0] right_top_grid_pin_47_ ;
input  [0:0] right_top_grid_pin_48_ ;
input  [0:0] right_top_grid_pin_49_ ;
input  [0:0] right_bottom_grid_pin_1_ ;
input  [0:19] chanx_left_in ;
input  [0:0] left_top_grid_pin_42_ ;
input  [0:0] left_top_grid_pin_43_ ;
input  [0:0] left_top_grid_pin_44_ ;
input  [0:0] left_top_grid_pin_45_ ;
input  [0:0] left_top_grid_pin_46_ ;
input  [0:0] left_top_grid_pin_47_ ;
input  [0:0] left_top_grid_pin_48_ ;
input  [0:0] left_top_grid_pin_49_ ;
input  [0:0] left_bottom_grid_pin_1_ ;
input  [0:0] ccff_head ;
output [0:19] chany_top_out ;
output [0:19] chanx_right_out ;
output [0:19] chanx_left_out ;
output [0:0] ccff_tail ;

wire [0:3] mux_tree_tapbuf_size10_0_sram ;
wire [0:3] mux_tree_tapbuf_size10_0_sram_inv ;
wire [0:0] mux_tree_tapbuf_size10_mem_0_ccff_tail ;
wire [0:3] mux_tree_tapbuf_size14_0_sram ;
wire [0:3] mux_tree_tapbuf_size14_0_sram_inv ;
wire [0:3] mux_tree_tapbuf_size14_1_sram ;
wire [0:3] mux_tree_tapbuf_size14_1_sram_inv ;
wire [0:0] mux_tree_tapbuf_size14_mem_0_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size14_mem_1_ccff_tail ;
wire [0:1] mux_tree_tapbuf_size2_0_sram ;
wire [0:1] mux_tree_tapbuf_size2_0_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_1_sram ;
wire [0:1] mux_tree_tapbuf_size2_1_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_2_sram ;
wire [0:1] mux_tree_tapbuf_size2_2_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_3_sram ;
wire [0:1] mux_tree_tapbuf_size2_3_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_4_sram ;
wire [0:1] mux_tree_tapbuf_size2_4_sram_inv ;
wire [0:0] mux_tree_tapbuf_size2_mem_0_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_1_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_2_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_3_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_4_ccff_tail ;
wire [0:1] mux_tree_tapbuf_size3_0_sram ;
wire [0:1] mux_tree_tapbuf_size3_0_sram_inv ;
wire [0:1] mux_tree_tapbuf_size3_1_sram ;
wire [0:1] mux_tree_tapbuf_size3_1_sram_inv ;
wire [0:1] mux_tree_tapbuf_size3_2_sram ;
wire [0:1] mux_tree_tapbuf_size3_2_sram_inv ;
wire [0:1] mux_tree_tapbuf_size3_3_sram ;
wire [0:1] mux_tree_tapbuf_size3_3_sram_inv ;
wire [0:1] mux_tree_tapbuf_size3_4_sram ;
wire [0:1] mux_tree_tapbuf_size3_4_sram_inv ;
wire [0:1] mux_tree_tapbuf_size3_5_sram ;
wire [0:1] mux_tree_tapbuf_size3_5_sram_inv ;
wire [0:1] mux_tree_tapbuf_size3_6_sram ;
wire [0:1] mux_tree_tapbuf_size3_6_sram_inv ;
wire [0:1] mux_tree_tapbuf_size3_7_sram ;
wire [0:1] mux_tree_tapbuf_size3_7_sram_inv ;
wire [0:0] mux_tree_tapbuf_size3_mem_0_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size3_mem_1_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size3_mem_2_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size3_mem_3_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size3_mem_4_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size3_mem_5_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size3_mem_6_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size3_mem_7_ccff_tail ;
wire [0:2] mux_tree_tapbuf_size4_0_sram ;
wire [0:2] mux_tree_tapbuf_size4_0_sram_inv ;
wire [0:2] mux_tree_tapbuf_size4_1_sram ;
wire [0:2] mux_tree_tapbuf_size4_1_sram_inv ;
wire [0:0] mux_tree_tapbuf_size4_mem_0_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size4_mem_1_ccff_tail ;
wire [0:2] mux_tree_tapbuf_size6_0_sram ;
wire [0:2] mux_tree_tapbuf_size6_0_sram_inv ;
wire [0:2] mux_tree_tapbuf_size6_1_sram ;
wire [0:2] mux_tree_tapbuf_size6_1_sram_inv ;
wire [0:0] mux_tree_tapbuf_size6_mem_0_ccff_tail ;
wire [0:2] mux_tree_tapbuf_size7_0_sram ;
wire [0:2] mux_tree_tapbuf_size7_0_sram_inv ;
wire [0:2] mux_tree_tapbuf_size7_1_sram ;
wire [0:2] mux_tree_tapbuf_size7_1_sram_inv ;
wire [0:2] mux_tree_tapbuf_size7_2_sram ;
wire [0:2] mux_tree_tapbuf_size7_2_sram_inv ;
wire [0:2] mux_tree_tapbuf_size7_3_sram ;
wire [0:2] mux_tree_tapbuf_size7_3_sram_inv ;
wire [0:2] mux_tree_tapbuf_size7_4_sram ;
wire [0:2] mux_tree_tapbuf_size7_4_sram_inv ;
wire [0:2] mux_tree_tapbuf_size7_5_sram ;
wire [0:2] mux_tree_tapbuf_size7_5_sram_inv ;
wire [0:2] mux_tree_tapbuf_size7_6_sram ;
wire [0:2] mux_tree_tapbuf_size7_6_sram_inv ;
wire [0:0] mux_tree_tapbuf_size7_mem_0_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size7_mem_1_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size7_mem_2_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size7_mem_3_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size7_mem_4_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size7_mem_5_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size7_mem_6_ccff_tail ;
wire [0:3] mux_tree_tapbuf_size8_0_sram ;
wire [0:3] mux_tree_tapbuf_size8_0_sram_inv ;
wire [0:3] mux_tree_tapbuf_size8_1_sram ;
wire [0:3] mux_tree_tapbuf_size8_1_sram_inv ;
wire [0:3] mux_tree_tapbuf_size8_2_sram ;
wire [0:3] mux_tree_tapbuf_size8_2_sram_inv ;
wire [0:3] mux_tree_tapbuf_size8_3_sram ;
wire [0:3] mux_tree_tapbuf_size8_3_sram_inv ;
wire [0:0] mux_tree_tapbuf_size8_mem_0_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size8_mem_1_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size8_mem_2_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size8_mem_3_ccff_tail ;
wire [0:3] mux_tree_tapbuf_size9_0_sram ;
wire [0:3] mux_tree_tapbuf_size9_0_sram_inv ;
wire [0:3] mux_tree_tapbuf_size9_1_sram ;
wire [0:3] mux_tree_tapbuf_size9_1_sram_inv ;
wire [0:0] mux_tree_tapbuf_size9_mem_0_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size9_mem_1_ccff_tail ;

mux_tree_tapbuf_size8 mux_top_track_0 (
    .in ( { top_left_grid_pin_34_[0] , top_left_grid_pin_36_[0] , 
        top_left_grid_pin_38_[0] , top_left_grid_pin_40_[0] , 
        chanx_right_in[1] , chanx_right_in[2] , chanx_left_in[0] , 
        chanx_left_in[2] } ) ,
    .sram ( mux_tree_tapbuf_size8_0_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size8_0_sram_inv ) , 
    .out ( chany_top_out[0] ) , .p0 ( optlc_net_114 ) ) ;
mux_tree_tapbuf_size8_2 mux_right_track_8 (
    .in ( { chany_top_in[2] , chany_top_in[9] , chany_top_in[16] , 
        right_top_grid_pin_42_[0] , right_top_grid_pin_46_[0] , 
        right_bottom_grid_pin_1_[0] , chanx_left_in[6] , chanx_left_in[16] } ) ,
    .sram ( mux_tree_tapbuf_size8_1_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size8_1_sram_inv ) , 
    .out ( chanx_right_out[4] ) , .p0 ( optlc_net_118 ) ) ;
mux_tree_tapbuf_size8_0 mux_left_track_3 (
    .in ( { chany_top_in[6] , chany_top_in[13] , chanx_right_in[4] , 
        chanx_right_in[13] , left_top_grid_pin_43_[0] , 
        left_top_grid_pin_45_[0] , left_top_grid_pin_47_[0] , 
        left_top_grid_pin_49_[0] } ) ,
    .sram ( mux_tree_tapbuf_size8_2_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size8_2_sram_inv ) , 
    .out ( chanx_left_out[1] ) , .p0 ( optlc_net_116 ) ) ;
mux_tree_tapbuf_size8_1 mux_left_track_9 (
    .in ( { chany_top_in[4] , chany_top_in[11] , chany_top_in[18] , 
        chanx_right_in[6] , chanx_right_in[16] , left_top_grid_pin_42_[0] , 
        left_top_grid_pin_46_[0] , left_bottom_grid_pin_1_[0] } ) ,
    .sram ( mux_tree_tapbuf_size8_3_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size8_3_sram_inv ) , 
    .out ( chanx_left_out[4] ) , .p0 ( optlc_net_114 ) ) ;
mux_tree_tapbuf_size8_mem mem_top_track_0 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( ccff_head ) , 
    .ccff_tail ( mux_tree_tapbuf_size8_mem_0_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size8_0_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size8_0_sram_inv ) ) ;
mux_tree_tapbuf_size8_mem_2 mem_right_track_8 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size14_mem_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size8_mem_1_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size8_1_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size8_1_sram_inv ) ) ;
mux_tree_tapbuf_size8_mem_0 mem_left_track_3 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size10_mem_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size8_mem_2_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size8_2_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size8_2_sram_inv ) ) ;
mux_tree_tapbuf_size8_mem_1 mem_left_track_9 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size14_mem_1_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size8_mem_3_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size8_3_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size8_3_sram_inv ) ) ;
mux_tree_tapbuf_size7_4 mux_top_track_2 (
    .in ( { top_left_grid_pin_35_[0] , top_left_grid_pin_37_[0] , 
        top_left_grid_pin_39_[0] , top_left_grid_pin_41_[0] , 
        chanx_right_in[3] , chanx_right_in[4] , chanx_left_in[4] } ) ,
    .sram ( mux_tree_tapbuf_size7_0_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size7_0_sram_inv ) , 
    .out ( chany_top_out[1] ) , .p0 ( optlc_net_115 ) ) ;
mux_tree_tapbuf_size7_5 mux_top_track_4 (
    .in ( { top_left_grid_pin_34_[0] , top_left_grid_pin_36_[0] , 
        top_left_grid_pin_38_[0] , top_left_grid_pin_40_[0] , 
        chanx_right_in[5] , chanx_right_in[7] , chanx_left_in[5] } ) ,
    .sram ( mux_tree_tapbuf_size7_1_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size7_1_sram_inv ) , 
    .out ( chany_top_out[2] ) , .p0 ( optlc_net_117 ) ) ;
mux_tree_tapbuf_size7_2 mux_top_track_6 (
    .in ( { top_left_grid_pin_35_[0] , top_left_grid_pin_37_[0] , 
        top_left_grid_pin_39_[0] , top_left_grid_pin_41_[0] , 
        chanx_right_in[6] , chanx_right_in[11] , chanx_left_in[6] } ) ,
    .sram ( mux_tree_tapbuf_size7_2_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size7_2_sram_inv ) , 
    .out ( chany_top_out[3] ) , .p0 ( optlc_net_117 ) ) ;
mux_tree_tapbuf_size7_2 mux_right_track_16 (
    .in ( { chany_top_in[3] , chany_top_in[10] , chany_top_in[17] , 
        right_top_grid_pin_43_[0] , right_top_grid_pin_47_[0] , 
        chanx_left_in[8] , chanx_left_in[17] } ) ,
    .sram ( mux_tree_tapbuf_size7_3_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size7_3_sram_inv ) , 
    .out ( chanx_right_out[8] ) , .p0 ( optlc_net_118 ) ) ;
mux_tree_tapbuf_size7_3 mux_right_track_24 (
    .in ( { chany_top_in[4] , chany_top_in[11] , chany_top_in[18] , 
        right_top_grid_pin_44_[0] , right_top_grid_pin_48_[0] , 
        chanx_left_in[9] , chanx_left_in[18] } ) ,
    .sram ( mux_tree_tapbuf_size7_4_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size7_4_sram_inv ) , 
    .out ( chanx_right_out[12] ) , .p0 ( optlc_net_117 ) ) ;
mux_tree_tapbuf_size7_0_1 mux_left_track_17 (
    .in ( { chany_top_in[3] , chany_top_in[10] , chany_top_in[17] , 
        chanx_right_in[8] , chanx_right_in[17] , left_top_grid_pin_43_[0] , 
        left_top_grid_pin_47_[0] } ) ,
    .sram ( mux_tree_tapbuf_size7_5_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size7_5_sram_inv ) , 
    .out ( chanx_left_out[8] ) , .p0 ( optlc_net_116 ) ) ;
mux_tree_tapbuf_size7_1_1 mux_left_track_25 (
    .in ( { chany_top_in[2] , chany_top_in[9] , chany_top_in[16] , 
        chanx_right_in[9] , chanx_right_in[18] , left_top_grid_pin_44_[0] , 
        left_top_grid_pin_48_[0] } ) ,
    .sram ( mux_tree_tapbuf_size7_6_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size7_6_sram_inv ) , 
    .out ( chanx_left_out[12] ) , .p0 ( optlc_net_116 ) ) ;
mux_tree_tapbuf_size7_mem_4 mem_top_track_2 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size8_mem_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size7_mem_0_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size7_0_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size7_0_sram_inv ) ) ;
mux_tree_tapbuf_size7_mem_5 mem_top_track_4 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size7_mem_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size7_mem_1_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size7_1_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size7_1_sram_inv ) ) ;
mux_tree_tapbuf_size7_mem_2 mem_top_track_6 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size7_mem_1_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size7_mem_2_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size7_2_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size7_2_sram_inv ) ) ;
mux_tree_tapbuf_size7_mem_2 mem_right_track_16 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size8_mem_1_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size7_mem_3_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size7_3_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size7_3_sram_inv ) ) ;
mux_tree_tapbuf_size7_mem_3 mem_right_track_24 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size7_mem_3_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size7_mem_4_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size7_4_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size7_4_sram_inv ) ) ;
mux_tree_tapbuf_size7_mem_0_1 mem_left_track_17 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size8_mem_3_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size7_mem_5_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size7_5_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size7_5_sram_inv ) ) ;
mux_tree_tapbuf_size7_mem_1_1 mem_left_track_25 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size7_mem_5_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size7_mem_6_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size7_6_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size7_6_sram_inv ) ) ;
mux_tree_tapbuf_size4_6 mux_top_track_8 (
    .in ( { top_left_grid_pin_34_[0] , chanx_right_in[8] , 
        chanx_right_in[15] , chanx_left_in[8] } ) ,
    .sram ( mux_tree_tapbuf_size4_0_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size4_0_sram_inv ) , 
    .out ( chany_top_out[4] ) , .p0 ( optlc_net_119 ) ) ;
mux_tree_tapbuf_size4_0_1 mux_top_track_10 (
    .in ( { top_left_grid_pin_35_[0] , chanx_right_in[9] , 
        chanx_right_in[19] , chanx_left_in[9] } ) ,
    .sram ( mux_tree_tapbuf_size4_1_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size4_1_sram_inv ) , 
    .out ( chany_top_out[5] ) , .p0 ( optlc_net_119 ) ) ;
mux_tree_tapbuf_size4_mem_6 mem_top_track_8 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size7_mem_2_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size4_mem_0_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size4_0_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size4_0_sram_inv ) ) ;
mux_tree_tapbuf_size4_mem_0_1 mem_top_track_10 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size4_mem_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size4_mem_1_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size4_1_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size4_1_sram_inv ) ) ;
mux_tree_tapbuf_size3_0_2 mux_top_track_12 (
    .in ( { top_left_grid_pin_36_[0] , chanx_right_in[10] , 
        chanx_left_in[10] } ) ,
    .sram ( mux_tree_tapbuf_size3_0_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size3_0_sram_inv ) , 
    .out ( chany_top_out[6] ) , .p0 ( optlc_net_117 ) ) ;
mux_tree_tapbuf_size3_1_1 mux_top_track_14 (
    .in ( { top_left_grid_pin_37_[0] , chanx_right_in[12] , 
        chanx_left_in[12] } ) ,
    .sram ( mux_tree_tapbuf_size3_1_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size3_1_sram_inv ) , 
    .out ( chany_top_out[7] ) , .p0 ( optlc_net_117 ) ) ;
mux_tree_tapbuf_size3_2_1 mux_top_track_16 (
    .in ( { top_left_grid_pin_38_[0] , chanx_right_in[13] , 
        chanx_left_in[13] } ) ,
    .sram ( mux_tree_tapbuf_size3_2_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size3_2_sram_inv ) , 
    .out ( chany_top_out[8] ) , .p0 ( optlc_net_114 ) ) ;
mux_tree_tapbuf_size3_3_1 mux_top_track_18 (
    .in ( { top_left_grid_pin_39_[0] , chanx_right_in[14] , 
        chanx_left_in[14] } ) ,
    .sram ( mux_tree_tapbuf_size3_3_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size3_3_sram_inv ) , 
    .out ( chany_top_out[9] ) , .p0 ( optlc_net_117 ) ) ;
mux_tree_tapbuf_size3_4 mux_top_track_20 (
    .in ( { top_left_grid_pin_40_[0] , chanx_right_in[16] , 
        chanx_left_in[16] } ) ,
    .sram ( mux_tree_tapbuf_size3_4_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size3_4_sram_inv ) , 
    .out ( chany_top_out[10] ) , .p0 ( optlc_net_117 ) ) ;
mux_tree_tapbuf_size3_5 mux_top_track_22 (
    .in ( { top_left_grid_pin_41_[0] , chanx_right_in[17] , 
        chanx_left_in[17] } ) ,
    .sram ( mux_tree_tapbuf_size3_5_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size3_5_sram_inv ) , 
    .out ( chany_top_out[11] ) , .p0 ( optlc_net_117 ) ) ;
mux_tree_tapbuf_size3_6 mux_top_track_24 (
    .in ( { top_left_grid_pin_34_[0] , chanx_right_in[18] , 
        chanx_left_in[18] } ) ,
    .sram ( mux_tree_tapbuf_size3_6_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size3_6_sram_inv ) , 
    .out ( chany_top_out[12] ) , .p0 ( optlc_net_116 ) ) ;
mux_tree_tapbuf_size3_7 mux_top_track_38 (
    .in ( { top_left_grid_pin_41_[0] , chanx_right_in[0] , chanx_left_in[1] } ) ,
    .sram ( mux_tree_tapbuf_size3_7_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size3_7_sram_inv ) , 
    .out ( chany_top_out[19] ) , .p0 ( optlc_net_115 ) ) ;
mux_tree_tapbuf_size3_mem_0_2 mem_top_track_12 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size4_mem_1_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size3_mem_0_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size3_0_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size3_0_sram_inv ) ) ;
mux_tree_tapbuf_size3_mem_1_1 mem_top_track_14 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size3_mem_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size3_mem_1_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size3_1_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size3_1_sram_inv ) ) ;
mux_tree_tapbuf_size3_mem_2_1 mem_top_track_16 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size3_mem_1_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size3_mem_2_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size3_2_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size3_2_sram_inv ) ) ;
mux_tree_tapbuf_size3_mem_3_1 mem_top_track_18 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size3_mem_2_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size3_mem_3_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size3_3_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size3_3_sram_inv ) ) ;
mux_tree_tapbuf_size3_mem_4 mem_top_track_20 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size3_mem_3_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size3_mem_4_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size3_4_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size3_4_sram_inv ) ) ;
mux_tree_tapbuf_size3_mem_5 mem_top_track_22 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size3_mem_4_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size3_mem_5_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size3_5_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size3_5_sram_inv ) ) ;
mux_tree_tapbuf_size3_mem_6 mem_top_track_24 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size3_mem_5_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size3_mem_6_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size3_6_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size3_6_sram_inv ) ) ;
mux_tree_tapbuf_size3_mem_7 mem_top_track_38 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_4_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size3_mem_7_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size3_7_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size3_7_sram_inv ) ) ;
mux_tree_tapbuf_size2_0_2 mux_top_track_28 (
    .in ( { top_left_grid_pin_36_[0] , chanx_left_in[19] } ) ,
    .sram ( mux_tree_tapbuf_size2_0_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_0_sram_inv ) ,
    .out ( { ropt_net_124 } ) ,
    .p0 ( optlc_net_114 ) ) ;
mux_tree_tapbuf_size2_1_2 mux_top_track_30 (
    .in ( { top_left_grid_pin_37_[0] , chanx_left_in[15] } ) ,
    .sram ( mux_tree_tapbuf_size2_1_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_1_sram_inv ) , 
    .out ( chany_top_out[15] ) , .p0 ( optlc_net_114 ) ) ;
mux_tree_tapbuf_size2_2_2 mux_top_track_32 (
    .in ( { top_left_grid_pin_38_[0] , chanx_left_in[11] } ) ,
    .sram ( mux_tree_tapbuf_size2_2_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_2_sram_inv ) , 
    .out ( chany_top_out[16] ) , .p0 ( optlc_net_114 ) ) ;
mux_tree_tapbuf_size2_3_2 mux_top_track_34 (
    .in ( { top_left_grid_pin_39_[0] , chanx_left_in[7] } ) ,
    .sram ( mux_tree_tapbuf_size2_3_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_3_sram_inv ) , 
    .out ( chany_top_out[17] ) , .p0 ( optlc_net_114 ) ) ;
mux_tree_tapbuf_size2_13 mux_top_track_36 (
    .in ( { top_left_grid_pin_40_[0] , chanx_left_in[3] } ) ,
    .sram ( mux_tree_tapbuf_size2_4_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_4_sram_inv ) , 
    .out ( chany_top_out[18] ) , .p0 ( optlc_net_115 ) ) ;
mux_tree_tapbuf_size2_mem_0_2 mem_top_track_28 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size3_mem_6_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_0_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_0_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_0_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem_1_2 mem_top_track_30 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_1_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_1_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_1_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem_2_2 mem_top_track_32 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_1_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_2_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_2_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_2_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem_3_2 mem_top_track_34 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_2_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_3_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_3_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_3_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem_13 mem_top_track_36 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_3_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_4_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_4_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_4_sram_inv ) ) ;
mux_tree_tapbuf_size9_0 mux_right_track_0 (
    .in ( { chany_top_in[6] , chany_top_in[13] , right_top_grid_pin_42_[0] , 
        right_top_grid_pin_44_[0] , right_top_grid_pin_46_[0] , 
        right_top_grid_pin_48_[0] , right_bottom_grid_pin_1_[0] , 
        chanx_left_in[2] , chanx_left_in[12] } ) ,
    .sram ( mux_tree_tapbuf_size9_0_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size9_0_sram_inv ) , 
    .out ( chanx_right_out[0] ) , .p0 ( optlc_net_119 ) ) ;
mux_tree_tapbuf_size9 mux_right_track_2 (
    .in ( { chany_top_in[0] , chany_top_in[7] , chany_top_in[14] , 
        right_top_grid_pin_43_[0] , right_top_grid_pin_45_[0] , 
        right_top_grid_pin_47_[0] , right_top_grid_pin_49_[0] , 
        chanx_left_in[4] , chanx_left_in[13] } ) ,
    .sram ( mux_tree_tapbuf_size9_1_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size9_1_sram_inv ) , 
    .out ( chanx_right_out[1] ) , .p0 ( optlc_net_119 ) ) ;
mux_tree_tapbuf_size9_mem_0 mem_right_track_0 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size3_mem_7_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size9_mem_0_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size9_0_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size9_0_sram_inv ) ) ;
mux_tree_tapbuf_size9_mem mem_right_track_2 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size9_mem_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size9_mem_1_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size9_1_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size9_1_sram_inv ) ) ;
mux_tree_tapbuf_size14 mux_right_track_4 (
    .in ( { chany_top_in[1] , chany_top_in[8] , chany_top_in[15] , 
        right_top_grid_pin_42_[0] , right_top_grid_pin_43_[0] , 
        right_top_grid_pin_44_[0] , right_top_grid_pin_45_[0] , 
        right_top_grid_pin_46_[0] , right_top_grid_pin_47_[0] , 
        right_top_grid_pin_48_[0] , right_top_grid_pin_49_[0] , 
        right_bottom_grid_pin_1_[0] , chanx_left_in[5] , chanx_left_in[14] } ) ,
    .sram ( mux_tree_tapbuf_size14_0_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size14_0_sram_inv ) , 
    .out ( chanx_right_out[2] ) , .p0 ( optlc_net_118 ) ) ;
mux_tree_tapbuf_size14_0 mux_left_track_5 (
    .in ( { chany_top_in[5] , chany_top_in[12] , chany_top_in[19] , 
        chanx_right_in[5] , chanx_right_in[14] , left_top_grid_pin_42_[0] , 
        left_top_grid_pin_43_[0] , left_top_grid_pin_44_[0] , 
        left_top_grid_pin_45_[0] , left_top_grid_pin_46_[0] , 
        left_top_grid_pin_47_[0] , left_top_grid_pin_48_[0] , 
        left_top_grid_pin_49_[0] , left_bottom_grid_pin_1_[0] } ) ,
    .sram ( mux_tree_tapbuf_size14_1_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size14_1_sram_inv ) , 
    .out ( chanx_left_out[2] ) , .p0 ( optlc_net_116 ) ) ;
mux_tree_tapbuf_size14_mem mem_right_track_4 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size9_mem_1_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size14_mem_0_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size14_0_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size14_0_sram_inv ) ) ;
mux_tree_tapbuf_size14_mem_0 mem_left_track_5 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size8_mem_2_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size14_mem_1_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size14_1_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size14_1_sram_inv ) ) ;
mux_tree_tapbuf_size6_6 mux_right_track_32 (
    .in ( { chany_top_in[5] , chany_top_in[12] , chany_top_in[19] , 
        right_top_grid_pin_45_[0] , right_top_grid_pin_49_[0] , 
        chanx_left_in[10] } ) ,
    .sram ( mux_tree_tapbuf_size6_0_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size6_0_sram_inv ) , 
    .out ( chanx_right_out[16] ) , .p0 ( optlc_net_118 ) ) ;
mux_tree_tapbuf_size6_0_2 mux_left_track_33 (
    .in ( { chany_top_in[1] , chany_top_in[8] , chany_top_in[15] , 
        chanx_right_in[10] , left_top_grid_pin_45_[0] , 
        left_top_grid_pin_49_[0] } ) ,
    .sram ( mux_tree_tapbuf_size6_1_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size6_1_sram_inv ) , 
    .out ( chanx_left_out[16] ) , .p0 ( optlc_net_116 ) ) ;
mux_tree_tapbuf_size6_mem_6 mem_right_track_32 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size7_mem_4_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size6_mem_0_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size6_0_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size6_0_sram_inv ) ) ;
mux_tree_tapbuf_size6_mem_0_2 mem_left_track_33 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size7_mem_6_ccff_tail ) , 
    .ccff_tail ( ccff_tail ) , .mem_out ( mux_tree_tapbuf_size6_1_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size6_1_sram_inv ) ) ;
mux_tree_tapbuf_size10 mux_left_track_1 (
    .in ( { chany_top_in[0] , chany_top_in[7] , chany_top_in[14] , 
        chanx_right_in[2] , chanx_right_in[12] , left_top_grid_pin_42_[0] , 
        left_top_grid_pin_44_[0] , left_top_grid_pin_46_[0] , 
        left_top_grid_pin_48_[0] , left_bottom_grid_pin_1_[0] } ) ,
    .sram ( mux_tree_tapbuf_size10_0_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size10_0_sram_inv ) , 
    .out ( chanx_left_out[0] ) , .p0 ( optlc_net_116 ) ) ;
mux_tree_tapbuf_size10_mem mem_left_track_1 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size6_mem_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size10_mem_0_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size10_0_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size10_0_sram_inv ) ) ;
sky130_fd_sc_hd__conb_1 optlc_109 ( .LO ( SYNOPSYS_UNCONNECTED_1 ) , 
    .HI ( optlc_net_114 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_111 ( .LO ( SYNOPSYS_UNCONNECTED_2 ) , 
    .HI ( optlc_net_115 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_3__2 ( .A ( chanx_right_in[4] ) , 
    .X ( ropt_net_133 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_113 ( .LO ( SYNOPSYS_UNCONNECTED_3 ) , 
    .HI ( optlc_net_116 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_117 ( .LO ( SYNOPSYS_UNCONNECTED_4 ) , 
    .HI ( optlc_net_117 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_742 ( .A ( ropt_net_138 ) , 
    .X ( chanx_left_out[7] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_745 ( .A ( ropt_net_139 ) , 
    .X ( chanx_left_out[5] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_716 ( .A ( chanx_right_in[17] ) , 
    .X ( chanx_left_out[18] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_746 ( .A ( ropt_net_140 ) , 
    .X ( chanx_right_out[18] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_10__9 ( .A ( chanx_right_in[13] ) , 
    .X ( ropt_net_148 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_11__10 ( .A ( chanx_right_in[14] ) , 
    .X ( chanx_left_out[15] ) ) ;
sky130_fd_sc_hd__conb_1 optlc_119 ( .LO ( SYNOPSYS_UNCONNECTED_5 ) , 
    .HI ( optlc_net_118 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_121 ( .LO ( SYNOPSYS_UNCONNECTED_6 ) , 
    .HI ( optlc_net_119 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_14__13 ( .A ( chanx_right_in[18] ) , 
    .X ( chanx_left_out[19] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_15__14 ( .A ( chanx_left_in[2] ) , 
    .X ( ropt_net_136 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_16__15 ( .A ( chanx_left_in[4] ) , 
    .X ( ropt_net_134 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_17__16 ( .A ( chanx_left_in[5] ) , 
    .X ( ropt_net_132 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_717 ( .A ( chanx_right_in[2] ) , 
    .X ( ropt_net_146 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_718 ( .A ( chanx_right_in[16] ) , 
    .X ( chanx_left_out[17] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_20__19 ( .A ( chanx_left_in[9] ) , 
    .X ( ropt_net_135 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_719 ( .A ( chanx_right_in[6] ) , 
    .X ( ropt_net_138 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_22__21 ( .A ( chanx_left_in[12] ) , 
    .X ( chanx_right_out[13] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_23__22 ( .A ( chanx_left_in[13] ) , 
    .X ( ropt_net_131 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_720 ( .A ( ropt_net_124 ) , 
    .X ( ropt_net_143 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_722 ( .A ( ropt_net_125 ) , 
    .X ( ropt_net_141 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_723 ( .A ( chanx_right_in[9] ) , 
    .X ( ropt_net_149 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_724 ( .A ( chanx_right_in[8] ) , 
    .X ( chanx_left_out[9] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_65 ( .A ( top_left_grid_pin_35_[0] ) , 
    .X ( BUF_net_65 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_725 ( .A ( chanx_right_in[12] ) , 
    .X ( ropt_net_147 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_67 ( .A ( chanx_right_in[5] ) , 
    .X ( BUF_net_67 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_747 ( .A ( ropt_net_141 ) , 
    .X ( chanx_right_out[7] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_748 ( .A ( ropt_net_142 ) , 
    .X ( chanx_left_out[6] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_749 ( .A ( ropt_net_143 ) , 
    .X ( chany_top_out[14] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_726 ( .A ( chanx_left_in[18] ) , 
    .X ( chanx_right_out[19] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_727 ( .A ( ropt_net_130 ) , 
    .X ( ropt_net_140 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_750 ( .A ( ropt_net_144 ) , 
    .X ( chanx_right_out[6] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_751 ( .A ( ropt_net_145 ) , 
    .X ( chanx_right_out[3] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_RR_75 ( .A ( chanx_left_in[8] ) , 
    .X ( chanx_right_out[9] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_RR_76 ( .A ( chanx_left_in[10] ) , 
    .X ( chanx_right_out[11] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_RR_77 ( .A ( chanx_left_in[14] ) , 
    .X ( chanx_right_out[15] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_78 ( .A ( chanx_left_in[17] ) , 
    .X ( ropt_net_130 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_752 ( .A ( ropt_net_146 ) , 
    .X ( chanx_left_out[3] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_728 ( .A ( ropt_net_131 ) , 
    .X ( chanx_right_out[14] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_729 ( .A ( ropt_net_132 ) , 
    .X ( ropt_net_144 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_730 ( .A ( ropt_net_133 ) , 
    .X ( ropt_net_139 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_732 ( .A ( ropt_net_134 ) , 
    .X ( chanx_right_out[5] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_734 ( .A ( ropt_net_135 ) , 
    .X ( chanx_right_out[10] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_735 ( .A ( ropt_net_136 ) , 
    .X ( ropt_net_145 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_753 ( .A ( ropt_net_147 ) , 
    .X ( chanx_left_out[13] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_P_92 ( .A ( chanx_left_in[16] ) , 
    .X ( chanx_right_out[17] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_754 ( .A ( ropt_net_148 ) , 
    .X ( chanx_left_out[14] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_756 ( .A ( ropt_net_149 ) , 
    .X ( chanx_left_out[10] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_P_98 ( .A ( chanx_right_in[10] ) , 
    .X ( chanx_left_out[11] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 BUFT_P_100 ( .A ( BUF_net_65 ) , 
    .X ( chany_top_out[13] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 BUFT_P_102 ( .A ( BUF_net_67 ) , 
    .X ( ropt_net_142 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_P_106 ( .A ( chanx_left_in[6] ) , 
    .X ( ropt_net_125 ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_1_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_8__39 ( .A ( mem_out[1] ) , 
    .X ( net_net_72 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_95 ( .A ( net_net_72 ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_3_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_7__38 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_2_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_6__37 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_0_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_5__36 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_5_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_4__35 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_12 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_3__34 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_6_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_2__33 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_4_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_1__32 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_33 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_1_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_33 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
endmodule


module const1_6_3 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_3_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_6_3 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
endmodule


module const1_5_3 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_2_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_5_3 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
endmodule


module const1_4_3 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_0_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_4_3 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
endmodule


module const1_3_3 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_5_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_3_3 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
endmodule


module const1_2_3 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_12 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_2_3 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
endmodule


module const1_1_3 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_6_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_1_3 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
endmodule


module const1_0_3 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_4_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_0_3 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
endmodule


module sb_0__2_ ( prog_clk , chanx_right_in , right_top_grid_pin_1_ , 
    chany_bottom_in , bottom_left_grid_pin_1_ , ccff_head , chanx_right_out , 
    chany_bottom_out , ccff_tail ) ;
input  [0:0] prog_clk ;
input  [0:19] chanx_right_in ;
input  [0:0] right_top_grid_pin_1_ ;
input  [0:19] chany_bottom_in ;
input  [0:0] bottom_left_grid_pin_1_ ;
input  [0:0] ccff_head ;
output [0:19] chanx_right_out ;
output [0:19] chany_bottom_out ;
output [0:0] ccff_tail ;

wire [0:1] mux_tree_tapbuf_size2_0_sram ;
wire [0:1] mux_tree_tapbuf_size2_0_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_1_sram ;
wire [0:1] mux_tree_tapbuf_size2_1_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_2_sram ;
wire [0:1] mux_tree_tapbuf_size2_2_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_3_sram ;
wire [0:1] mux_tree_tapbuf_size2_3_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_4_sram ;
wire [0:1] mux_tree_tapbuf_size2_4_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_5_sram ;
wire [0:1] mux_tree_tapbuf_size2_5_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_6_sram ;
wire [0:1] mux_tree_tapbuf_size2_6_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_7_sram ;
wire [0:1] mux_tree_tapbuf_size2_7_sram_inv ;
wire [0:0] mux_tree_tapbuf_size2_mem_0_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_1_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_2_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_3_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_4_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_5_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_6_ccff_tail ;

mux_tree_tapbuf_size2_4_1 mux_right_track_0 (
    .in ( { right_top_grid_pin_1_[0] , chany_bottom_in[18] } ) ,
    .sram ( mux_tree_tapbuf_size2_0_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_0_sram_inv ) , 
    .out ( chanx_right_out[0] ) , .p0 ( optlc_net_110 ) ) ;
mux_tree_tapbuf_size2_6_1 mux_right_track_4 (
    .in ( { right_top_grid_pin_1_[0] , chany_bottom_in[16] } ) ,
    .sram ( mux_tree_tapbuf_size2_1_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_1_sram_inv ) , 
    .out ( chanx_right_out[2] ) , .p0 ( optlc_net_110 ) ) ;
mux_tree_tapbuf_size2_12 mux_right_track_8 (
    .in ( { right_top_grid_pin_1_[0] , chany_bottom_in[14] } ) ,
    .sram ( mux_tree_tapbuf_size2_2_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_2_sram_inv ) , 
    .out ( chanx_right_out[4] ) , .p0 ( optlc_net_110 ) ) ;
mux_tree_tapbuf_size2_5_1 mux_right_track_24 (
    .in ( { right_top_grid_pin_1_[0] , chany_bottom_in[6] } ) ,
    .sram ( mux_tree_tapbuf_size2_3_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_3_sram_inv ) , 
    .out ( chanx_right_out[12] ) , .p0 ( optlc_net_110 ) ) ;
mux_tree_tapbuf_size2_0_1 mux_bottom_track_1 (
    .in ( { chanx_right_in[18] , bottom_left_grid_pin_1_[0] } ) ,
    .sram ( mux_tree_tapbuf_size2_4_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_4_sram_inv ) , 
    .out ( chany_bottom_out[0] ) , .p0 ( optlc_net_109 ) ) ;
mux_tree_tapbuf_size2_2_1 mux_bottom_track_5 (
    .in ( { chanx_right_in[16] , bottom_left_grid_pin_1_[0] } ) ,
    .sram ( mux_tree_tapbuf_size2_5_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_5_sram_inv ) , 
    .out ( chany_bottom_out[2] ) , .p0 ( optlc_net_109 ) ) ;
mux_tree_tapbuf_size2_3_1 mux_bottom_track_9 (
    .in ( { chanx_right_in[14] , bottom_left_grid_pin_1_[0] } ) ,
    .sram ( mux_tree_tapbuf_size2_6_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_6_sram_inv ) , 
    .out ( chany_bottom_out[4] ) , .p0 ( optlc_net_109 ) ) ;
mux_tree_tapbuf_size2_1_1 mux_bottom_track_25 (
    .in ( { chanx_right_in[6] , bottom_left_grid_pin_1_[0] } ) ,
    .sram ( mux_tree_tapbuf_size2_7_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_7_sram_inv ) , 
    .out ( chany_bottom_out[12] ) , .p0 ( optlc_net_109 ) ) ;
mux_tree_tapbuf_size2_mem_4_1 mem_right_track_0 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( ccff_head ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_0_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_0_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_0_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem_6_1 mem_right_track_4 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_1_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_1_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_1_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem_12 mem_right_track_8 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_1_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_2_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_2_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_2_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem_5_1 mem_right_track_24 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_2_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_3_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_3_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_3_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem_0_1 mem_bottom_track_1 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_3_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_4_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_4_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_4_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem_2_1 mem_bottom_track_5 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_4_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_5_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_5_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_5_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem_3_1 mem_bottom_track_9 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_5_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_6_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_6_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_6_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem_1_1 mem_bottom_track_25 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_6_ccff_tail ) ,
    .ccff_tail ( { ropt_net_138 } ) ,
    .mem_out ( mux_tree_tapbuf_size2_7_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_7_sram_inv ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_730 ( .A ( ropt_net_140 ) , 
    .X ( chanx_right_out[13] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_731 ( .A ( ropt_net_141 ) , 
    .X ( chany_bottom_out[5] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_732 ( .A ( ropt_net_142 ) , 
    .X ( chany_bottom_out[7] ) ) ;
sky130_fd_sc_hd__conb_1 optlc_110 ( .LO ( SYNOPSYS_UNCONNECTED_1 ) , 
    .HI ( optlc_net_109 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_733 ( .A ( ropt_net_143 ) , 
    .X ( chany_bottom_out[3] ) ) ;
sky130_fd_sc_hd__conb_1 optlc_112 ( .LO ( SYNOPSYS_UNCONNECTED_2 ) , 
    .HI ( optlc_net_110 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_734 ( .A ( ropt_net_144 ) , 
    .X ( chany_bottom_out[15] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_701 ( .A ( ropt_net_111 ) , 
    .X ( ropt_net_146 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_702 ( .A ( chany_bottom_in[3] ) , 
    .X ( ropt_net_156 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_735 ( .A ( ropt_net_145 ) , 
    .X ( chany_bottom_out[10] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_703 ( .A ( chany_bottom_in[9] ) , 
    .X ( ropt_net_154 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_704 ( .A ( ropt_net_114 ) , 
    .X ( ropt_net_143 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_705 ( .A ( chany_bottom_in[5] ) , 
    .X ( ropt_net_140 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_736 ( .A ( ropt_net_146 ) , 
    .X ( chany_bottom_out[16] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_706 ( .A ( ropt_net_116 ) , 
    .X ( chany_bottom_out[11] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_16__15 ( .A ( chanx_right_in[19] ) , 
    .X ( aps_rename_8_ ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_707 ( .A ( chanx_right_in[1] ) , 
    .X ( ropt_net_155 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_708 ( .A ( chanx_right_in[3] ) , 
    .X ( ropt_net_144 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_709 ( .A ( chany_bottom_in[2] ) , 
    .X ( ropt_net_160 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_710 ( .A ( ropt_net_120 ) , 
    .X ( ropt_net_148 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_711 ( .A ( chany_bottom_in[7] ) , 
    .X ( ropt_net_157 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_712 ( 
    .A ( chany_bottom_in[12] ) , .X ( chanx_right_out[6] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_713 ( .A ( chanx_right_in[9] ) , 
    .X ( ropt_net_162 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_714 ( .A ( chanx_right_in[13] ) , 
    .X ( ropt_net_141 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_715 ( .A ( ropt_net_125 ) , 
    .X ( ropt_net_145 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_716 ( .A ( chanx_right_in[12] ) , 
    .X ( ropt_net_158 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_717 ( 
    .A ( chany_bottom_in[15] ) , .X ( ropt_net_161 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_718 ( .A ( chany_bottom_in[0] ) , 
    .X ( ropt_net_153 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_719 ( .A ( ropt_net_129 ) , 
    .X ( ropt_net_142 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_720 ( .A ( chanx_right_in[5] ) , 
    .X ( ropt_net_147 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_721 ( 
    .A ( chany_bottom_in[17] ) , .X ( ropt_net_159 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_722 ( .A ( ropt_net_132 ) , 
    .X ( chanx_right_out[7] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_40 ( .A ( chanx_right_in[0] ) , 
    .X ( BUF_net_40 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_737 ( .A ( ropt_net_147 ) , 
    .X ( chany_bottom_out[13] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_738 ( .A ( ropt_net_148 ) , 
    .X ( chany_bottom_out[8] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_723 ( 
    .A ( chany_bottom_in[19] ) , .X ( chanx_right_out[19] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_44 ( .A ( chanx_right_in[4] ) , 
    .X ( BUF_net_44 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_739 ( .A ( ropt_net_149 ) , 
    .X ( ccff_tail[0] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_740 ( .A ( ropt_net_150 ) , 
    .X ( chanx_right_out[14] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_47 ( .A ( chanx_right_in[8] ) , 
    .X ( ropt_net_125 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_724 ( .A ( ropt_net_134 ) , 
    .X ( ropt_net_151 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_741 ( .A ( ropt_net_151 ) , 
    .X ( chany_bottom_out[1] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_725 ( .A ( ropt_net_135 ) , 
    .X ( ropt_net_150 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_726 ( .A ( ropt_net_136 ) , 
    .X ( chanx_right_out[5] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_727 ( .A ( ropt_net_137 ) , 
    .X ( chanx_right_out[8] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_742 ( .A ( ropt_net_152 ) , 
    .X ( chany_bottom_out[14] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_54 ( .A ( chanx_right_in[17] ) , 
    .X ( ropt_net_134 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_728 ( .A ( ropt_net_138 ) , 
    .X ( ropt_net_149 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_743 ( .A ( ropt_net_153 ) , 
    .X ( chanx_right_out[18] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_57 ( .A ( chany_bottom_in[1] ) , 
    .X ( BUF_net_57 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_744 ( .A ( ropt_net_154 ) , 
    .X ( chanx_right_out[9] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_745 ( .A ( ropt_net_155 ) , 
    .X ( chany_bottom_out[17] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_60 ( .A ( chany_bottom_in[4] ) , 
    .X ( ropt_net_135 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_746 ( .A ( ropt_net_156 ) , 
    .X ( chanx_right_out[15] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_747 ( .A ( ropt_net_157 ) , 
    .X ( chanx_right_out[11] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_729 ( .A ( ropt_net_139 ) , 
    .X ( chanx_right_out[10] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_748 ( .A ( ropt_net_158 ) , 
    .X ( chany_bottom_out[6] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_RR_65 ( .A ( chany_bottom_in[10] ) , 
    .X ( ropt_net_137 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_RR_66 ( .A ( chany_bottom_in[11] ) , 
    .X ( ropt_net_132 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_749 ( .A ( ropt_net_159 ) , 
    .X ( chanx_right_out[1] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_751 ( .A ( ropt_net_160 ) , 
    .X ( chanx_right_out[16] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_753 ( .A ( ropt_net_161 ) , 
    .X ( chanx_right_out[3] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_754 ( .A ( ropt_net_162 ) , 
    .X ( chany_bottom_out[9] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 BUFT_RR_76 ( .A ( chanx_right_in[7] ) , 
    .X ( ropt_net_116 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_79 ( .A ( chanx_right_in[10] ) , 
    .X ( ropt_net_120 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_83 ( .A ( chanx_right_in[15] ) , 
    .X ( ropt_net_114 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 BUFT_P_91 ( .A ( BUF_net_40 ) , 
    .X ( chany_bottom_out[18] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_P_92 ( .A ( chanx_right_in[2] ) , 
    .X ( ropt_net_111 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 BUFT_P_93 ( .A ( BUF_net_44 ) , 
    .X ( ropt_net_152 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 BUFT_P_94 ( .A ( aps_rename_8_ ) , 
    .X ( chany_bottom_out[19] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_P_100 ( .A ( chanx_right_in[11] ) , 
    .X ( ropt_net_129 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 BUFT_P_104 ( .A ( BUF_net_57 ) , 
    .X ( chanx_right_out[17] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_P_106 ( .A ( chany_bottom_in[8] ) , 
    .X ( ropt_net_139 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_P_107 ( .A ( chany_bottom_in[13] ) , 
    .X ( ropt_net_136 ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_11 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_28__58 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_32 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_11 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_32 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
endmodule


module mux_tree_tapbuf_size3_mem_0_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd1_1 FTB_27__57 ( .A ( mem_out[1] ) , 
    .X ( net_net_100 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_100 ( .A ( net_net_100 ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size3_mem_4 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_26__56 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size3_mem_3 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_25__55 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size3_mem_2 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_24__54 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size3_mem_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_23__53 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_26_1 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size3_0_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:2] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_26_1 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( p0 ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_8 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , .X ( out[0] ) ) ;
endmodule


module const1_25_1 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size3_4 ( in , sram , sram_inv , out , p0 ) ;
input  [0:2] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;

const1_25_1 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( p0 ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
endmodule


module const1_24_1 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size3_3 ( in , sram , sram_inv , out , p0 ) ;
input  [0:2] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;

const1_24_1 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( p0 ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
endmodule


module const1_23_1 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size3_2 ( in , sram , sram_inv , out , p0 ) ;
input  [0:2] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;

const1_23_1 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( p0 ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
endmodule


module const1_22_1 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size3_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:2] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;

const1_22_1 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( p0 ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
endmodule


module mux_tree_tapbuf_size7_mem ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_22__52 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size7_mem_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_21__51 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size7_mem_0 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_20__50 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_21_1 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size7 ( in , sram , sram_inv , out , p0 ) ;
input  [0:6] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;

const1_21_1 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_3_ ( .A0 ( p0 ) , .A1 ( in[6] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
endmodule


module const1_20_1 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size7_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:6] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;

const1_20_1 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_3_ ( .A0 ( p0 ) , .A1 ( in[6] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
endmodule


module const1_19_1 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size7_0 ( in , sram , sram_inv , out , p0 ) ;
input  [0:6] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;

const1_19_1 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_3_ ( .A0 ( p0 ) , .A1 ( in[6] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
endmodule


module mux_tree_tapbuf_size4_mem_3 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_19__49 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size4_mem_2 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_18__48 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size4_mem_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_17__47 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size4_mem_0 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_16__46 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size4_mem_4 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_15__45 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size4_mem ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_14__44 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size4_mem_5 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_13__43 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_18_1 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size4_3 ( in , sram , sram_inv , out , p0 ) ;
input  [0:3] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;

const1_18_1 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( in[2] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , .A1 ( in[3] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
endmodule


module const1_17_1 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size4_2 ( in , sram , sram_inv , out , p0 ) ;
input  [0:3] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;

const1_17_1 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( in[2] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , .A1 ( in[3] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
endmodule


module const1_16_2 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size4_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:3] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;

const1_16_2 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( in[2] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , .A1 ( in[3] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
endmodule


module const1_15_2 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size4_0 ( in , sram , sram_inv , out , p0 ) ;
input  [0:3] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;

const1_15_2 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( in[2] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , .A1 ( in[3] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
endmodule


module const1_14_2 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size4_4 ( in , sram , sram_inv , out , p0 ) ;
input  [0:3] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;

const1_14_2 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( in[2] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , .A1 ( in[3] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
endmodule


module const1_13_2 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size4 ( in , sram , sram_inv , out , p0 ) ;
input  [0:3] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;

const1_13_2 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( in[2] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , .A1 ( in[3] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
endmodule


module const1_12_2 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size4_5 ( in , sram , sram_inv , out , p0 ) ;
input  [0:3] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;

const1_12_2 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( in[2] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , .A1 ( in[3] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
endmodule


module mux_tree_tapbuf_size5_mem_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_12__42 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size5_mem_0_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_11__41 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size5_mem_2 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_10__40 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size5_mem_3 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_9__39 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size5_mem_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_8__38 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_11_2 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size5_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:4] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;

const1_11_2 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , .A1 ( in[4] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
endmodule


module const1_10_2 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size5_0_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:4] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;

const1_10_2 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , .A1 ( in[4] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
endmodule


module const1_9_2 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size5_2 ( in , sram , sram_inv , out , p0 ) ;
input  [0:4] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;

const1_9_2 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , .A1 ( in[4] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
endmodule


module const1_8_2 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size5_3 ( in , sram , sram_inv , out , p0 ) ;
input  [0:4] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;

const1_8_2 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , .A1 ( in[4] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
endmodule


module const1_7_2 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size5_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:4] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;

const1_7_2 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , .A1 ( in[4] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
endmodule


module mux_tree_tapbuf_size6_mem_2 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_7__37 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size6_mem_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_6__36 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size6_mem_0_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_5__35 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size6_mem_3 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_4__34 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size6_mem_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_3__33 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size6_mem_5 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_2__32 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size6_mem_4 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_1__31 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_6_2 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size6_2 ( in , sram , sram_inv , out , p0 ) ;
input  [0:5] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;

const1_6_2 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
endmodule


module const1_5_2 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size6_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:5] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;

const1_5_2 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
endmodule


module const1_4_2 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size6_0_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:5] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;

const1_4_2 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_8 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , .X ( out[0] ) ) ;
endmodule


module const1_3_2 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size6_3 ( in , sram , sram_inv , out , p0 ) ;
input  [0:5] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;

const1_3_2 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
endmodule


module const1_2_2 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size6_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:5] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;

const1_2_2 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
endmodule


module const1_1_2 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size6_5 ( in , sram , sram_inv , out , p0 ) ;
input  [0:5] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;

const1_1_2 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
endmodule


module const1_0_2 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size6_4 ( in , sram , sram_inv , out , p0 ) ;
input  [0:5] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;

const1_0_2 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
endmodule


module sb_0__1_ ( prog_clk , chany_top_in , top_left_grid_pin_1_ , 
    chanx_right_in , right_top_grid_pin_42_ , right_top_grid_pin_43_ , 
    right_top_grid_pin_44_ , right_top_grid_pin_45_ , right_top_grid_pin_46_ , 
    right_top_grid_pin_47_ , right_top_grid_pin_48_ , right_top_grid_pin_49_ , 
    chany_bottom_in , bottom_left_grid_pin_1_ , ccff_head , chany_top_out , 
    chanx_right_out , chany_bottom_out , ccff_tail ) ;
input  [0:0] prog_clk ;
input  [0:19] chany_top_in ;
input  [0:0] top_left_grid_pin_1_ ;
input  [0:19] chanx_right_in ;
input  [0:0] right_top_grid_pin_42_ ;
input  [0:0] right_top_grid_pin_43_ ;
input  [0:0] right_top_grid_pin_44_ ;
input  [0:0] right_top_grid_pin_45_ ;
input  [0:0] right_top_grid_pin_46_ ;
input  [0:0] right_top_grid_pin_47_ ;
input  [0:0] right_top_grid_pin_48_ ;
input  [0:0] right_top_grid_pin_49_ ;
input  [0:19] chany_bottom_in ;
input  [0:0] bottom_left_grid_pin_1_ ;
input  [0:0] ccff_head ;
output [0:19] chany_top_out ;
output [0:19] chanx_right_out ;
output [0:19] chany_bottom_out ;
output [0:0] ccff_tail ;

wire [0:1] mux_tree_tapbuf_size2_0_sram ;
wire [0:1] mux_tree_tapbuf_size2_0_sram_inv ;
wire [0:0] mux_tree_tapbuf_size2_mem_0_ccff_tail ;
wire [0:1] mux_tree_tapbuf_size3_0_sram ;
wire [0:1] mux_tree_tapbuf_size3_0_sram_inv ;
wire [0:1] mux_tree_tapbuf_size3_1_sram ;
wire [0:1] mux_tree_tapbuf_size3_1_sram_inv ;
wire [0:1] mux_tree_tapbuf_size3_2_sram ;
wire [0:1] mux_tree_tapbuf_size3_2_sram_inv ;
wire [0:1] mux_tree_tapbuf_size3_3_sram ;
wire [0:1] mux_tree_tapbuf_size3_3_sram_inv ;
wire [0:1] mux_tree_tapbuf_size3_4_sram ;
wire [0:1] mux_tree_tapbuf_size3_4_sram_inv ;
wire [0:0] mux_tree_tapbuf_size3_mem_0_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size3_mem_1_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size3_mem_2_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size3_mem_3_ccff_tail ;
wire [0:2] mux_tree_tapbuf_size4_0_sram ;
wire [0:2] mux_tree_tapbuf_size4_0_sram_inv ;
wire [0:2] mux_tree_tapbuf_size4_1_sram ;
wire [0:2] mux_tree_tapbuf_size4_1_sram_inv ;
wire [0:2] mux_tree_tapbuf_size4_2_sram ;
wire [0:2] mux_tree_tapbuf_size4_2_sram_inv ;
wire [0:2] mux_tree_tapbuf_size4_3_sram ;
wire [0:2] mux_tree_tapbuf_size4_3_sram_inv ;
wire [0:2] mux_tree_tapbuf_size4_4_sram ;
wire [0:2] mux_tree_tapbuf_size4_4_sram_inv ;
wire [0:2] mux_tree_tapbuf_size4_5_sram ;
wire [0:2] mux_tree_tapbuf_size4_5_sram_inv ;
wire [0:2] mux_tree_tapbuf_size4_6_sram ;
wire [0:2] mux_tree_tapbuf_size4_6_sram_inv ;
wire [0:0] mux_tree_tapbuf_size4_mem_0_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size4_mem_1_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size4_mem_2_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size4_mem_3_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size4_mem_4_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size4_mem_5_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size4_mem_6_ccff_tail ;
wire [0:2] mux_tree_tapbuf_size5_0_sram ;
wire [0:2] mux_tree_tapbuf_size5_0_sram_inv ;
wire [0:2] mux_tree_tapbuf_size5_1_sram ;
wire [0:2] mux_tree_tapbuf_size5_1_sram_inv ;
wire [0:2] mux_tree_tapbuf_size5_2_sram ;
wire [0:2] mux_tree_tapbuf_size5_2_sram_inv ;
wire [0:2] mux_tree_tapbuf_size5_3_sram ;
wire [0:2] mux_tree_tapbuf_size5_3_sram_inv ;
wire [0:2] mux_tree_tapbuf_size5_4_sram ;
wire [0:2] mux_tree_tapbuf_size5_4_sram_inv ;
wire [0:0] mux_tree_tapbuf_size5_mem_0_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size5_mem_1_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size5_mem_2_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size5_mem_3_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size5_mem_4_ccff_tail ;
wire [0:2] mux_tree_tapbuf_size6_0_sram ;
wire [0:2] mux_tree_tapbuf_size6_0_sram_inv ;
wire [0:2] mux_tree_tapbuf_size6_1_sram ;
wire [0:2] mux_tree_tapbuf_size6_1_sram_inv ;
wire [0:2] mux_tree_tapbuf_size6_2_sram ;
wire [0:2] mux_tree_tapbuf_size6_2_sram_inv ;
wire [0:2] mux_tree_tapbuf_size6_3_sram ;
wire [0:2] mux_tree_tapbuf_size6_3_sram_inv ;
wire [0:2] mux_tree_tapbuf_size6_4_sram ;
wire [0:2] mux_tree_tapbuf_size6_4_sram_inv ;
wire [0:2] mux_tree_tapbuf_size6_5_sram ;
wire [0:2] mux_tree_tapbuf_size6_5_sram_inv ;
wire [0:2] mux_tree_tapbuf_size6_6_sram ;
wire [0:2] mux_tree_tapbuf_size6_6_sram_inv ;
wire [0:0] mux_tree_tapbuf_size6_mem_0_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size6_mem_1_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size6_mem_2_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size6_mem_3_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size6_mem_4_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size6_mem_5_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size6_mem_6_ccff_tail ;
wire [0:2] mux_tree_tapbuf_size7_0_sram ;
wire [0:2] mux_tree_tapbuf_size7_0_sram_inv ;
wire [0:2] mux_tree_tapbuf_size7_1_sram ;
wire [0:2] mux_tree_tapbuf_size7_1_sram_inv ;
wire [0:2] mux_tree_tapbuf_size7_2_sram ;
wire [0:2] mux_tree_tapbuf_size7_2_sram_inv ;
wire [0:0] mux_tree_tapbuf_size7_mem_0_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size7_mem_1_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size7_mem_2_ccff_tail ;

mux_tree_tapbuf_size6_4 mux_top_track_0 (
    .in ( { top_left_grid_pin_1_[0] , chanx_right_in[1] , chanx_right_in[8] , 
        chanx_right_in[15] , chany_bottom_in[2] , chany_bottom_in[12] } ) ,
    .sram ( mux_tree_tapbuf_size6_0_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size6_0_sram_inv ) , 
    .out ( chany_top_out[0] ) , .p0 ( optlc_net_125 ) ) ;
mux_tree_tapbuf_size6_5 mux_top_track_4 (
    .in ( { top_left_grid_pin_1_[0] , chanx_right_in[3] , chanx_right_in[10] , 
        chanx_right_in[17] , chany_bottom_in[5] , chany_bottom_in[14] } ) ,
    .sram ( mux_tree_tapbuf_size6_1_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size6_1_sram_inv ) , 
    .out ( chany_top_out[2] ) , .p0 ( optlc_net_122 ) ) ;
mux_tree_tapbuf_size6_1 mux_top_track_8 (
    .in ( { top_left_grid_pin_1_[0] , chanx_right_in[4] , chanx_right_in[11] , 
        chanx_right_in[18] , chany_bottom_in[6] , chany_bottom_in[16] } ) ,
    .sram ( mux_tree_tapbuf_size6_2_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size6_2_sram_inv ) , 
    .out ( chany_top_out[4] ) , .p0 ( optlc_net_124 ) ) ;
mux_tree_tapbuf_size6_3 mux_right_track_0 (
    .in ( { chany_top_in[2] , right_top_grid_pin_42_[0] , 
        right_top_grid_pin_44_[0] , right_top_grid_pin_46_[0] , 
        right_top_grid_pin_48_[0] , chany_bottom_in[2] } ) ,
    .sram ( mux_tree_tapbuf_size6_3_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size6_3_sram_inv ) , 
    .out ( chanx_right_out[0] ) , .p0 ( optlc_net_125 ) ) ;
mux_tree_tapbuf_size6_0_1 mux_bottom_track_1 (
    .in ( { chany_top_in[2] , chany_top_in[12] , chanx_right_in[5] , 
        chanx_right_in[12] , chanx_right_in[19] , bottom_left_grid_pin_1_[0] } ) ,
    .sram ( mux_tree_tapbuf_size6_4_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size6_4_sram_inv ) , 
    .out ( chany_bottom_out[0] ) , .p0 ( optlc_net_124 ) ) ;
mux_tree_tapbuf_size6_1 mux_bottom_track_5 (
    .in ( { chany_top_in[5] , chany_top_in[14] , chanx_right_in[3] , 
        chanx_right_in[10] , chanx_right_in[17] , bottom_left_grid_pin_1_[0] } ) ,
    .sram ( mux_tree_tapbuf_size6_5_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size6_5_sram_inv ) , 
    .out ( chany_bottom_out[2] ) , .p0 ( optlc_net_122 ) ) ;
mux_tree_tapbuf_size6_2 mux_bottom_track_9 (
    .in ( { chany_top_in[6] , chany_top_in[16] , chanx_right_in[2] , 
        chanx_right_in[9] , chanx_right_in[16] , bottom_left_grid_pin_1_[0] } ) ,
    .sram ( mux_tree_tapbuf_size6_6_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size6_6_sram_inv ) , 
    .out ( chany_bottom_out[4] ) , .p0 ( optlc_net_122 ) ) ;
mux_tree_tapbuf_size6_mem_4 mem_top_track_0 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( ccff_head ) , 
    .ccff_tail ( mux_tree_tapbuf_size6_mem_0_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size6_0_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size6_0_sram_inv ) ) ;
mux_tree_tapbuf_size6_mem_5 mem_top_track_4 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size5_mem_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size6_mem_1_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size6_1_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size6_1_sram_inv ) ) ;
mux_tree_tapbuf_size6_mem_1 mem_top_track_8 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size6_mem_1_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size6_mem_2_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size6_2_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size6_2_sram_inv ) ) ;
mux_tree_tapbuf_size6_mem_3 mem_right_track_0 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size4_mem_1_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size6_mem_3_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size6_3_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size6_3_sram_inv ) ) ;
mux_tree_tapbuf_size6_mem_0_1 mem_bottom_track_1 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size6_mem_4_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size6_4_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size6_4_sram_inv ) ) ;
mux_tree_tapbuf_size6_mem_1 mem_bottom_track_5 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size5_mem_2_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size6_mem_5_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size6_5_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size6_5_sram_inv ) ) ;
mux_tree_tapbuf_size6_mem_2 mem_bottom_track_9 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size6_mem_5_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size6_mem_6_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size6_6_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size6_6_sram_inv ) ) ;
mux_tree_tapbuf_size5_1 mux_top_track_2 (
    .in ( { chanx_right_in[2] , chanx_right_in[9] , chanx_right_in[16] , 
        chany_bottom_in[4] , chany_bottom_in[13] } ) ,
    .sram ( mux_tree_tapbuf_size5_0_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size5_0_sram_inv ) , 
    .out ( chany_top_out[1] ) , .p0 ( optlc_net_122 ) ) ;
mux_tree_tapbuf_size5_3 mux_top_track_16 (
    .in ( { chanx_right_in[5] , chanx_right_in[12] , chanx_right_in[19] , 
        chany_bottom_in[8] , chany_bottom_in[17] } ) ,
    .sram ( mux_tree_tapbuf_size5_1_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size5_1_sram_inv ) , 
    .out ( chany_top_out[8] ) , .p0 ( optlc_net_124 ) ) ;
mux_tree_tapbuf_size5_2 mux_bottom_track_3 (
    .in ( { chany_top_in[4] , chany_top_in[13] , chanx_right_in[4] , 
        chanx_right_in[11] , chanx_right_in[18] } ) ,
    .sram ( mux_tree_tapbuf_size5_2_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size5_2_sram_inv ) , 
    .out ( chany_bottom_out[1] ) , .p0 ( optlc_net_122 ) ) ;
mux_tree_tapbuf_size5_0_1 mux_bottom_track_17 (
    .in ( { chany_top_in[8] , chany_top_in[17] , chanx_right_in[1] , 
        chanx_right_in[8] , chanx_right_in[15] } ) ,
    .sram ( mux_tree_tapbuf_size5_3_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size5_3_sram_inv ) , 
    .out ( chany_bottom_out[8] ) , .p0 ( optlc_net_122 ) ) ;
mux_tree_tapbuf_size5_1 mux_bottom_track_25 (
    .in ( { chany_top_in[9] , chany_top_in[18] , chanx_right_in[0] , 
        chanx_right_in[7] , chanx_right_in[14] } ) ,
    .sram ( mux_tree_tapbuf_size5_4_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size5_4_sram_inv ) , 
    .out ( chany_bottom_out[12] ) , .p0 ( optlc_net_124 ) ) ;
mux_tree_tapbuf_size5_mem_1 mem_top_track_2 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size6_mem_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size5_mem_0_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size5_0_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size5_0_sram_inv ) ) ;
mux_tree_tapbuf_size5_mem_3 mem_top_track_16 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size6_mem_2_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size5_mem_1_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size5_1_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size5_1_sram_inv ) ) ;
mux_tree_tapbuf_size5_mem_2 mem_bottom_track_3 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size6_mem_4_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size5_mem_2_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size5_2_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size5_2_sram_inv ) ) ;
mux_tree_tapbuf_size5_mem_0_1 mem_bottom_track_17 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size6_mem_6_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size5_mem_3_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size5_3_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size5_3_sram_inv ) ) ;
mux_tree_tapbuf_size5_mem_1 mem_bottom_track_25 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size5_mem_3_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size5_mem_4_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size5_4_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size5_4_sram_inv ) ) ;
mux_tree_tapbuf_size4_5 mux_top_track_24 (
    .in ( { chanx_right_in[6] , chanx_right_in[13] , chany_bottom_in[9] , 
        chany_bottom_in[18] } ) ,
    .sram ( mux_tree_tapbuf_size4_0_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size4_0_sram_inv ) , 
    .out ( chany_top_out[12] ) , .p0 ( optlc_net_123 ) ) ;
mux_tree_tapbuf_size4 mux_top_track_32 (
    .in ( { chanx_right_in[0] , chanx_right_in[7] , chanx_right_in[14] , 
        chany_bottom_in[10] } ) ,
    .sram ( mux_tree_tapbuf_size4_1_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size4_1_sram_inv ) , 
    .out ( chany_top_out[16] ) , .p0 ( optlc_net_123 ) ) ;
mux_tree_tapbuf_size4_4 mux_right_track_8 (
    .in ( { chany_top_in[7] , chany_top_in[8] , right_top_grid_pin_42_[0] , 
        chany_bottom_in[8] } ) ,
    .sram ( mux_tree_tapbuf_size4_2_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size4_2_sram_inv ) , 
    .out ( chanx_right_out[4] ) , .p0 ( optlc_net_123 ) ) ;
mux_tree_tapbuf_size4_0 mux_right_track_10 (
    .in ( { chany_top_in[9] , chany_top_in[11] , right_top_grid_pin_43_[0] , 
        chany_bottom_in[9] } ) ,
    .sram ( mux_tree_tapbuf_size4_3_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size4_3_sram_inv ) , 
    .out ( chanx_right_out[5] ) , .p0 ( optlc_net_123 ) ) ;
mux_tree_tapbuf_size4_1 mux_right_track_12 (
    .in ( { chany_top_in[10] , chany_top_in[15] , right_top_grid_pin_44_[0] , 
        chany_bottom_in[10] } ) ,
    .sram ( mux_tree_tapbuf_size4_4_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size4_4_sram_inv ) , 
    .out ( chanx_right_out[6] ) , .p0 ( optlc_net_123 ) ) ;
mux_tree_tapbuf_size4_2 mux_right_track_14 (
    .in ( { chany_top_in[12] , chany_top_in[19] , right_top_grid_pin_45_[0] , 
        chany_bottom_in[12] } ) ,
    .sram ( mux_tree_tapbuf_size4_5_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size4_5_sram_inv ) , 
    .out ( chanx_right_out[7] ) , .p0 ( optlc_net_125 ) ) ;
mux_tree_tapbuf_size4_3 mux_right_track_24 (
    .in ( { chany_top_in[18] , right_top_grid_pin_42_[0] , 
        chany_bottom_in[18] , chany_bottom_in[19] } ) ,
    .sram ( mux_tree_tapbuf_size4_6_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size4_6_sram_inv ) , 
    .out ( chanx_right_out[12] ) , .p0 ( optlc_net_124 ) ) ;
mux_tree_tapbuf_size4_mem_5 mem_top_track_24 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size5_mem_1_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size4_mem_0_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size4_0_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size4_0_sram_inv ) ) ;
mux_tree_tapbuf_size4_mem mem_top_track_32 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size4_mem_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size4_mem_1_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size4_1_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size4_1_sram_inv ) ) ;
mux_tree_tapbuf_size4_mem_4 mem_right_track_8 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size7_mem_2_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size4_mem_2_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size4_2_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size4_2_sram_inv ) ) ;
mux_tree_tapbuf_size4_mem_0 mem_right_track_10 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size4_mem_2_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size4_mem_3_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size4_3_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size4_3_sram_inv ) ) ;
mux_tree_tapbuf_size4_mem_1 mem_right_track_12 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size4_mem_3_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size4_mem_4_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size4_4_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size4_4_sram_inv ) ) ;
mux_tree_tapbuf_size4_mem_2 mem_right_track_14 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size4_mem_4_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size4_mem_5_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size4_5_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size4_5_sram_inv ) ) ;
mux_tree_tapbuf_size4_mem_3 mem_right_track_24 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size3_mem_3_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size4_mem_6_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size4_6_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size4_6_sram_inv ) ) ;
mux_tree_tapbuf_size7_0 mux_right_track_2 (
    .in ( { chany_top_in[0] , chany_top_in[4] , right_top_grid_pin_43_[0] , 
        right_top_grid_pin_45_[0] , right_top_grid_pin_47_[0] , 
        right_top_grid_pin_49_[0] , chany_bottom_in[4] } ) ,
    .sram ( mux_tree_tapbuf_size7_0_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size7_0_sram_inv ) , 
    .out ( chanx_right_out[1] ) , .p0 ( optlc_net_125 ) ) ;
mux_tree_tapbuf_size7_1 mux_right_track_4 (
    .in ( { chany_top_in[1] , chany_top_in[5] , right_top_grid_pin_42_[0] , 
        right_top_grid_pin_44_[0] , right_top_grid_pin_46_[0] , 
        right_top_grid_pin_48_[0] , chany_bottom_in[5] } ) ,
    .sram ( mux_tree_tapbuf_size7_1_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size7_1_sram_inv ) , 
    .out ( chanx_right_out[2] ) , .p0 ( optlc_net_125 ) ) ;
mux_tree_tapbuf_size7 mux_right_track_6 (
    .in ( { chany_top_in[3] , chany_top_in[6] , right_top_grid_pin_43_[0] , 
        right_top_grid_pin_45_[0] , right_top_grid_pin_47_[0] , 
        right_top_grid_pin_49_[0] , chany_bottom_in[6] } ) ,
    .sram ( mux_tree_tapbuf_size7_2_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size7_2_sram_inv ) , 
    .out ( chanx_right_out[3] ) , .p0 ( optlc_net_125 ) ) ;
mux_tree_tapbuf_size7_mem_0 mem_right_track_2 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size6_mem_3_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size7_mem_0_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size7_0_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size7_0_sram_inv ) ) ;
mux_tree_tapbuf_size7_mem_1 mem_right_track_4 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size7_mem_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size7_mem_1_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size7_1_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size7_1_sram_inv ) ) ;
mux_tree_tapbuf_size7_mem mem_right_track_6 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size7_mem_1_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size7_mem_2_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size7_2_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size7_2_sram_inv ) ) ;
mux_tree_tapbuf_size3_1 mux_right_track_16 (
    .in ( { chany_top_in[13] , right_top_grid_pin_46_[0] , 
        chany_bottom_in[13] } ) ,
    .sram ( mux_tree_tapbuf_size3_0_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size3_0_sram_inv ) , 
    .out ( chanx_right_out[8] ) , .p0 ( optlc_net_125 ) ) ;
mux_tree_tapbuf_size3_2 mux_right_track_18 (
    .in ( { chany_top_in[14] , right_top_grid_pin_47_[0] , 
        chany_bottom_in[14] } ) ,
    .sram ( mux_tree_tapbuf_size3_1_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size3_1_sram_inv ) , 
    .out ( chanx_right_out[9] ) , .p0 ( optlc_net_125 ) ) ;
mux_tree_tapbuf_size3_3 mux_right_track_20 (
    .in ( { chany_top_in[16] , right_top_grid_pin_48_[0] , 
        chany_bottom_in[16] } ) ,
    .sram ( mux_tree_tapbuf_size3_2_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size3_2_sram_inv ) , 
    .out ( chanx_right_out[10] ) , .p0 ( optlc_net_125 ) ) ;
mux_tree_tapbuf_size3_4 mux_right_track_22 (
    .in ( { chany_top_in[17] , right_top_grid_pin_49_[0] , 
        chany_bottom_in[17] } ) ,
    .sram ( mux_tree_tapbuf_size3_3_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size3_3_sram_inv ) , 
    .out ( chanx_right_out[11] ) , .p0 ( optlc_net_123 ) ) ;
mux_tree_tapbuf_size3_0_1 mux_bottom_track_33 (
    .in ( { chany_top_in[10] , chanx_right_in[6] , chanx_right_in[13] } ) ,
    .sram ( mux_tree_tapbuf_size3_4_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size3_4_sram_inv ) , 
    .out ( chany_bottom_out[16] ) , .p0 ( optlc_net_124 ) ) ;
mux_tree_tapbuf_size3_mem_1 mem_right_track_16 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size4_mem_5_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size3_mem_0_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size3_0_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size3_0_sram_inv ) ) ;
mux_tree_tapbuf_size3_mem_2 mem_right_track_18 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size3_mem_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size3_mem_1_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size3_1_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size3_1_sram_inv ) ) ;
mux_tree_tapbuf_size3_mem_3 mem_right_track_20 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size3_mem_1_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size3_mem_2_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size3_2_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size3_2_sram_inv ) ) ;
mux_tree_tapbuf_size3_mem_4 mem_right_track_22 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size3_mem_2_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size3_mem_3_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size3_3_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size3_3_sram_inv ) ) ;
mux_tree_tapbuf_size3_mem_0_1 mem_bottom_track_33 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size5_mem_4_ccff_tail ) ,
    .ccff_tail ( { ropt_net_130 } ) ,
    .mem_out ( mux_tree_tapbuf_size3_4_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size3_4_sram_inv ) ) ;
mux_tree_tapbuf_size2_11 mux_right_track_26 (
    .in ( { right_top_grid_pin_43_[0] , chany_bottom_in[15] } ) ,
    .sram ( mux_tree_tapbuf_size2_0_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_0_sram_inv ) , 
    .out ( chanx_right_out[13] ) , .p0 ( optlc_net_124 ) ) ;
mux_tree_tapbuf_size2_mem_11 mem_right_track_26 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size4_mem_6_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_0_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_0_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_0_sram_inv ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_1__0 ( .A ( chany_top_in[2] ) , 
    .X ( ropt_net_149 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_2__1 ( .A ( chany_top_in[4] ) , 
    .X ( ropt_net_150 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_111 ( .LO ( SYNOPSYS_UNCONNECTED_1 ) , 
    .HI ( optlc_net_122 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_746 ( .A ( ropt_net_153 ) , 
    .X ( chany_top_out[14] ) ) ;
sky130_fd_sc_hd__conb_1 optlc_113 ( .LO ( SYNOPSYS_UNCONNECTED_2 ) , 
    .HI ( optlc_net_123 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_115 ( .LO ( SYNOPSYS_UNCONNECTED_3 ) , 
    .HI ( optlc_net_124 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_7__6 ( .A ( chany_top_in[10] ) , 
    .X ( ropt_net_145 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_8__7 ( .A ( chany_top_in[12] ) , 
    .X ( ropt_net_152 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_748 ( .A ( ropt_net_154 ) , 
    .X ( chany_bottom_out[7] ) ) ;
sky130_fd_sc_hd__conb_1 optlc_117 ( .LO ( SYNOPSYS_UNCONNECTED_4 ) , 
    .HI ( optlc_net_125 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_716 ( .A ( chany_bottom_in[2] ) , 
    .X ( chany_top_out[3] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_749 ( .A ( ropt_net_155 ) , 
    .X ( chany_bottom_out[5] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_717 ( .A ( chany_top_in[14] ) , 
    .X ( chany_bottom_out[15] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_718 ( .A ( chany_top_in[6] ) , 
    .X ( ropt_net_154 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_719 ( .A ( ropt_net_129 ) , 
    .X ( chany_bottom_out[6] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_720 ( .A ( ropt_net_130 ) , 
    .X ( ropt_net_157 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_721 ( .A ( chany_top_in[13] ) , 
    .X ( ropt_net_156 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_722 ( .A ( chany_top_in[17] ) , 
    .X ( ropt_net_160 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_19__18 ( .A ( chany_bottom_in[5] ) , 
    .X ( ropt_net_144 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_723 ( .A ( chany_top_in[16] ) , 
    .X ( ropt_net_169 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_724 ( .A ( ropt_net_134 ) , 
    .X ( chany_top_out[5] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_725 ( .A ( ropt_net_135 ) , 
    .X ( ropt_net_167 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_726 ( .A ( ropt_net_136 ) , 
    .X ( ropt_net_159 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_24__23 ( .A ( chany_bottom_in[10] ) , 
    .X ( chany_top_out[11] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_727 ( .A ( ropt_net_137 ) , 
    .X ( ropt_net_158 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_26__25 ( .A ( chany_bottom_in[12] ) , 
    .X ( ropt_net_148 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_728 ( .A ( ropt_net_138 ) , 
    .X ( ropt_net_168 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_729 ( .A ( ropt_net_139 ) , 
    .X ( ropt_net_153 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_730 ( .A ( ropt_net_140 ) , 
    .X ( chanx_right_out[16] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_731 ( .A ( ropt_net_141 ) , 
    .X ( chany_top_out[18] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_732 ( .A ( ropt_net_142 ) , 
    .X ( chany_top_out[10] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_750 ( .A ( ropt_net_156 ) , 
    .X ( chany_bottom_out[14] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_733 ( .A ( ropt_net_143 ) , 
    .X ( chany_top_out[7] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_70 ( .A ( chany_top_in[9] ) , 
    .X ( ropt_net_137 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_751 ( .A ( ropt_net_157 ) , 
    .X ( ccff_tail[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_72 ( .A ( chany_bottom_in[0] ) , 
    .X ( BUF_net_72 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_RR_73 ( .A ( chany_bottom_in[1] ) , 
    .X ( ropt_net_147 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_752 ( .A ( ropt_net_158 ) , 
    .X ( chany_bottom_out[10] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_RR_75 ( .A ( chany_bottom_in[3] ) , 
    .X ( ropt_net_140 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_RR_76 ( .A ( chany_bottom_in[4] ) , 
    .X ( ropt_net_134 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_RR_77 ( .A ( chany_bottom_in[6] ) , 
    .X ( ropt_net_143 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_78 ( .A ( chany_bottom_in[7] ) , 
    .X ( ropt_net_135 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_RR_79 ( .A ( chany_bottom_in[9] ) , 
    .X ( ropt_net_142 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_80 ( .A ( chany_bottom_in[11] ) , 
    .X ( BUF_net_80 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_81 ( .A ( chany_bottom_in[13] ) , 
    .X ( ropt_net_139 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_82 ( .A ( chany_bottom_in[14] ) , 
    .X ( ropt_net_138 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_RR_83 ( .A ( chany_bottom_in[16] ) , 
    .X ( chany_top_out[17] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_RR_84 ( .A ( chany_bottom_in[17] ) , 
    .X ( ropt_net_141 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_RR_85 ( .A ( chany_bottom_in[18] ) , 
    .X ( chany_top_out[19] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_734 ( .A ( ropt_net_144 ) , 
    .X ( ropt_net_165 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_735 ( .A ( ropt_net_145 ) , 
    .X ( ropt_net_161 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_736 ( .A ( ropt_net_146 ) , 
    .X ( ropt_net_166 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_737 ( .A ( ropt_net_147 ) , 
    .X ( chanx_right_out[17] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_740 ( .A ( ropt_net_148 ) , 
    .X ( ropt_net_162 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_742 ( .A ( ropt_net_149 ) , 
    .X ( ropt_net_164 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_753 ( .A ( ropt_net_159 ) , 
    .X ( chany_bottom_out[9] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_P_98 ( .A ( chany_top_in[18] ) , 
    .X ( ropt_net_146 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_P_99 ( .A ( chany_bottom_in[8] ) , 
    .X ( ropt_net_151 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 BUFT_P_103 ( .A ( chany_top_in[5] ) , 
    .X ( ropt_net_129 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_P_104 ( .A ( chany_top_in[8] ) , 
    .X ( ropt_net_136 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_743 ( .A ( ropt_net_150 ) , 
    .X ( ropt_net_155 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_744 ( .A ( ropt_net_151 ) , 
    .X ( chany_top_out[9] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 BUFT_P_107 ( .A ( BUF_net_72 ) , 
    .X ( chanx_right_out[18] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 BUFT_P_108 ( .A ( BUF_net_80 ) , 
    .X ( chanx_right_out[14] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_745 ( .A ( ropt_net_152 ) , 
    .X ( ropt_net_163 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_755 ( .A ( ropt_net_160 ) , 
    .X ( chany_bottom_out[18] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_757 ( .A ( ropt_net_161 ) , 
    .X ( chany_bottom_out[11] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_758 ( .A ( ropt_net_162 ) , 
    .X ( chany_top_out[13] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_759 ( .A ( ropt_net_163 ) , 
    .X ( chany_bottom_out[13] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_760 ( .A ( ropt_net_164 ) , 
    .X ( chany_bottom_out[3] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_761 ( .A ( ropt_net_165 ) , 
    .X ( chany_top_out[6] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_762 ( .A ( ropt_net_166 ) , 
    .X ( chany_bottom_out[19] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_763 ( .A ( ropt_net_167 ) , 
    .X ( chanx_right_out[15] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_766 ( .A ( ropt_net_168 ) , 
    .X ( chany_top_out[15] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_770 ( .A ( ropt_net_169 ) , 
    .X ( chany_bottom_out[17] ) ) ;
endmodule


module mux_tree_tapbuf_size3_mem_0 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_18__39 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size3_mem ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_17__38 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_31 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size3_0 ( in , sram , sram_inv , out , p0 ) ;
input  [0:2] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;

const1_31 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( p0 ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
endmodule


module const1_16_1 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size3 ( in , sram , sram_inv , out , p0 ) ;
input  [0:2] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;

const1_16_1 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( p0 ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
endmodule


module mux_tree_tapbuf_size5_mem ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_16__37 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size5_mem_0 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_15__36 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_15_1 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size5 ( in , sram , sram_inv , out , p0 ) ;
input  [0:4] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;

const1_15_1 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , .A1 ( in[4] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
endmodule


module const1_14_1 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size5_0 ( in , sram , sram_inv , out , p0 ) ;
input  [0:4] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;

const1_14_1 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , .A1 ( in[4] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
endmodule


module mux_tree_tapbuf_size6_mem ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_14__35 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size6_mem_0 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_13__34 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_13_1 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size6 ( in , sram , sram_inv , out , p0 ) ;
input  [0:5] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;

const1_13_1 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
endmodule


module const1_12_1 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size6_0 ( in , sram , sram_inv , out , p0 ) ;
input  [0:5] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;

const1_12_1 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_7 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_12__33 ( .A ( mem_out[1] ) , 
    .X ( net_aps_33 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_52 ( .A ( net_aps_33 ) , 
    .X ( BUF_net_52 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_P_74 ( .A ( BUF_net_52 ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_6 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_11__32 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_5 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_10__31 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_4 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_9__30 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_3 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_8__29 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_2 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_7__28 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_6__27 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_0 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_5__26 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_9 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_4__25 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_3__24 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_10 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_2__23 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_8 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_1__22 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_11_1 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_7 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_11_1 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
endmodule


module const1_10_1 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_6 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_10_1 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
endmodule


module const1_9_1 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_5 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_9_1 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
endmodule


module const1_8_1 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_4 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_8_1 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
endmodule


module const1_7_1 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_3 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_7_1 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
endmodule


module const1_6_1 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_2 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_6_1 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
endmodule


module const1_5_1 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_5_1 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
endmodule


module const1_4_1 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_0 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_4_1 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
endmodule


module const1_3_1 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_9 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_3_1 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_P_68 ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
endmodule


module const1_2_1 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_2_1 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
endmodule


module const1_1_1 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_10 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_1_1 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
endmodule


module const1_0_1 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_8 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_0_1 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
endmodule


module sb_0__0_ ( prog_clk , chany_top_in , top_left_grid_pin_1_ , 
    chanx_right_in , right_top_grid_pin_42_ , right_top_grid_pin_43_ , 
    right_top_grid_pin_44_ , right_top_grid_pin_45_ , right_top_grid_pin_46_ , 
    right_top_grid_pin_47_ , right_top_grid_pin_48_ , right_top_grid_pin_49_ , 
    right_bottom_grid_pin_1_ , ccff_head , chany_top_out , chanx_right_out , 
    ccff_tail ) ;
input  [0:0] prog_clk ;
input  [0:19] chany_top_in ;
input  [0:0] top_left_grid_pin_1_ ;
input  [0:19] chanx_right_in ;
input  [0:0] right_top_grid_pin_42_ ;
input  [0:0] right_top_grid_pin_43_ ;
input  [0:0] right_top_grid_pin_44_ ;
input  [0:0] right_top_grid_pin_45_ ;
input  [0:0] right_top_grid_pin_46_ ;
input  [0:0] right_top_grid_pin_47_ ;
input  [0:0] right_top_grid_pin_48_ ;
input  [0:0] right_top_grid_pin_49_ ;
input  [0:0] right_bottom_grid_pin_1_ ;
input  [0:0] ccff_head ;
output [0:19] chany_top_out ;
output [0:19] chanx_right_out ;
output [0:0] ccff_tail ;

wire [0:1] mux_tree_tapbuf_size2_0_sram ;
wire [0:1] mux_tree_tapbuf_size2_0_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_10_sram ;
wire [0:1] mux_tree_tapbuf_size2_10_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_11_sram ;
wire [0:1] mux_tree_tapbuf_size2_11_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_1_sram ;
wire [0:1] mux_tree_tapbuf_size2_1_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_2_sram ;
wire [0:1] mux_tree_tapbuf_size2_2_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_3_sram ;
wire [0:1] mux_tree_tapbuf_size2_3_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_4_sram ;
wire [0:1] mux_tree_tapbuf_size2_4_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_5_sram ;
wire [0:1] mux_tree_tapbuf_size2_5_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_6_sram ;
wire [0:1] mux_tree_tapbuf_size2_6_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_7_sram ;
wire [0:1] mux_tree_tapbuf_size2_7_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_8_sram ;
wire [0:1] mux_tree_tapbuf_size2_8_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_9_sram ;
wire [0:1] mux_tree_tapbuf_size2_9_sram_inv ;
wire [0:0] mux_tree_tapbuf_size2_mem_0_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_10_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_1_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_2_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_3_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_4_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_5_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_6_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_7_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_8_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_9_ccff_tail ;
wire [0:1] mux_tree_tapbuf_size3_0_sram ;
wire [0:1] mux_tree_tapbuf_size3_0_sram_inv ;
wire [0:1] mux_tree_tapbuf_size3_1_sram ;
wire [0:1] mux_tree_tapbuf_size3_1_sram_inv ;
wire [0:0] mux_tree_tapbuf_size3_mem_0_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size3_mem_1_ccff_tail ;
wire [0:2] mux_tree_tapbuf_size5_0_sram ;
wire [0:2] mux_tree_tapbuf_size5_0_sram_inv ;
wire [0:2] mux_tree_tapbuf_size5_1_sram ;
wire [0:2] mux_tree_tapbuf_size5_1_sram_inv ;
wire [0:0] mux_tree_tapbuf_size5_mem_0_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size5_mem_1_ccff_tail ;
wire [0:2] mux_tree_tapbuf_size6_0_sram ;
wire [0:2] mux_tree_tapbuf_size6_0_sram_inv ;
wire [0:2] mux_tree_tapbuf_size6_1_sram ;
wire [0:2] mux_tree_tapbuf_size6_1_sram_inv ;
wire [0:0] mux_tree_tapbuf_size6_mem_0_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size6_mem_1_ccff_tail ;

mux_tree_tapbuf_size2_8 mux_top_track_0 (
    .in ( { top_left_grid_pin_1_[0] , chanx_right_in[1] } ) ,
    .sram ( mux_tree_tapbuf_size2_0_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_0_sram_inv ) , 
    .out ( chany_top_out[0] ) , .p0 ( optlc_net_80 ) ) ;
mux_tree_tapbuf_size2_10 mux_top_track_4 (
    .in ( { top_left_grid_pin_1_[0] , chanx_right_in[3] } ) ,
    .sram ( mux_tree_tapbuf_size2_1_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_1_sram_inv ) , 
    .out ( chany_top_out[2] ) , .p0 ( optlc_net_80 ) ) ;
mux_tree_tapbuf_size2 mux_top_track_8 (
    .in ( { top_left_grid_pin_1_[0] , chanx_right_in[5] } ) ,
    .sram ( mux_tree_tapbuf_size2_2_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_2_sram_inv ) , 
    .out ( chany_top_out[4] ) , .p0 ( optlc_net_80 ) ) ;
mux_tree_tapbuf_size2_9 mux_top_track_24 (
    .in ( { top_left_grid_pin_1_[0] , chanx_right_in[13] } ) ,
    .sram ( mux_tree_tapbuf_size2_3_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_3_sram_inv ) ,
    .out ( { ropt_net_91 } ) ,
    .p0 ( optlc_net_81 ) ) ;
mux_tree_tapbuf_size2_0 mux_right_track_10 (
    .in ( { chany_top_in[4] , right_top_grid_pin_43_[0] } ) ,
    .sram ( mux_tree_tapbuf_size2_4_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_4_sram_inv ) , 
    .out ( chanx_right_out[5] ) , .p0 ( optlc_net_81 ) ) ;
mux_tree_tapbuf_size2_1 mux_right_track_12 (
    .in ( { chany_top_in[5] , right_top_grid_pin_44_[0] } ) ,
    .sram ( mux_tree_tapbuf_size2_5_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_5_sram_inv ) , 
    .out ( chanx_right_out[6] ) , .p0 ( optlc_net_80 ) ) ;
mux_tree_tapbuf_size2_2 mux_right_track_14 (
    .in ( { chany_top_in[6] , right_top_grid_pin_45_[0] } ) ,
    .sram ( mux_tree_tapbuf_size2_6_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_6_sram_inv ) , 
    .out ( chanx_right_out[7] ) , .p0 ( optlc_net_79 ) ) ;
mux_tree_tapbuf_size2_3 mux_right_track_16 (
    .in ( { chany_top_in[7] , right_top_grid_pin_46_[0] } ) ,
    .sram ( mux_tree_tapbuf_size2_7_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_7_sram_inv ) , 
    .out ( chanx_right_out[8] ) , .p0 ( optlc_net_82 ) ) ;
mux_tree_tapbuf_size2_4 mux_right_track_18 (
    .in ( { chany_top_in[8] , right_top_grid_pin_47_[0] } ) ,
    .sram ( mux_tree_tapbuf_size2_8_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_8_sram_inv ) , 
    .out ( chanx_right_out[9] ) , .p0 ( optlc_net_82 ) ) ;
mux_tree_tapbuf_size2_5 mux_right_track_20 (
    .in ( { chany_top_in[9] , right_top_grid_pin_48_[0] } ) ,
    .sram ( mux_tree_tapbuf_size2_9_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_9_sram_inv ) , 
    .out ( chanx_right_out[10] ) , .p0 ( optlc_net_82 ) ) ;
mux_tree_tapbuf_size2_6 mux_right_track_22 (
    .in ( { chany_top_in[10] , right_top_grid_pin_49_[0] } ) ,
    .sram ( mux_tree_tapbuf_size2_10_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_10_sram_inv ) , 
    .out ( chanx_right_out[11] ) , .p0 ( optlc_net_82 ) ) ;
mux_tree_tapbuf_size2_7 mux_right_track_26 (
    .in ( { chany_top_in[12] , right_top_grid_pin_43_[0] } ) ,
    .sram ( mux_tree_tapbuf_size2_11_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_11_sram_inv ) , 
    .out ( chanx_right_out[13] ) , .p0 ( optlc_net_79 ) ) ;
mux_tree_tapbuf_size2_mem_8 mem_top_track_0 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( ccff_head ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_0_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_0_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_0_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem_10 mem_top_track_4 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_1_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_1_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_1_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem mem_top_track_8 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_1_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_2_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_2_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_2_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem_9 mem_top_track_24 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_2_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_3_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_3_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_3_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem_0 mem_right_track_10 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size3_mem_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_4_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_4_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_4_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem_1 mem_right_track_12 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_4_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_5_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_5_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_5_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem_2 mem_right_track_14 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_5_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_6_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_6_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_6_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem_3 mem_right_track_16 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_6_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_7_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_7_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_7_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem_4 mem_right_track_18 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_7_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_8_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_8_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_8_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem_5 mem_right_track_20 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_8_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_9_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_9_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_9_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem_6 mem_right_track_22 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_9_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_10_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_10_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_10_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem_7 mem_right_track_26 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size3_mem_1_ccff_tail ) ,
    .ccff_tail ( { ropt_net_83 } ) ,
    .mem_out ( mux_tree_tapbuf_size2_11_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_11_sram_inv ) ) ;
mux_tree_tapbuf_size6_0 mux_right_track_0 (
    .in ( { chany_top_in[19] , right_top_grid_pin_42_[0] , 
        right_top_grid_pin_44_[0] , right_top_grid_pin_46_[0] , 
        right_top_grid_pin_48_[0] , right_bottom_grid_pin_1_[0] } ) ,
    .sram ( mux_tree_tapbuf_size6_0_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size6_0_sram_inv ) , 
    .out ( chanx_right_out[0] ) , .p0 ( optlc_net_81 ) ) ;
mux_tree_tapbuf_size6 mux_right_track_4 (
    .in ( { chany_top_in[1] , right_top_grid_pin_42_[0] , 
        right_top_grid_pin_44_[0] , right_top_grid_pin_46_[0] , 
        right_top_grid_pin_48_[0] , right_bottom_grid_pin_1_[0] } ) ,
    .sram ( mux_tree_tapbuf_size6_1_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size6_1_sram_inv ) , 
    .out ( chanx_right_out[2] ) , .p0 ( optlc_net_79 ) ) ;
mux_tree_tapbuf_size6_mem_0 mem_right_track_0 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_3_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size6_mem_0_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size6_0_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size6_0_sram_inv ) ) ;
mux_tree_tapbuf_size6_mem mem_right_track_4 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size5_mem_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size6_mem_1_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size6_1_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size6_1_sram_inv ) ) ;
mux_tree_tapbuf_size5_0 mux_right_track_2 (
    .in ( { chany_top_in[0] , right_top_grid_pin_43_[0] , 
        right_top_grid_pin_45_[0] , right_top_grid_pin_47_[0] , 
        right_top_grid_pin_49_[0] } ) ,
    .sram ( mux_tree_tapbuf_size5_0_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size5_0_sram_inv ) , 
    .out ( chanx_right_out[1] ) , .p0 ( optlc_net_79 ) ) ;
mux_tree_tapbuf_size5 mux_right_track_6 (
    .in ( { chany_top_in[2] , right_top_grid_pin_43_[0] , 
        right_top_grid_pin_45_[0] , right_top_grid_pin_47_[0] , 
        right_top_grid_pin_49_[0] } ) ,
    .sram ( mux_tree_tapbuf_size5_1_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size5_1_sram_inv ) , 
    .out ( chanx_right_out[3] ) , .p0 ( optlc_net_79 ) ) ;
mux_tree_tapbuf_size5_mem_0 mem_right_track_2 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size6_mem_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size5_mem_0_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size5_0_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size5_0_sram_inv ) ) ;
mux_tree_tapbuf_size5_mem mem_right_track_6 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size6_mem_1_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size5_mem_1_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size5_1_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size5_1_sram_inv ) ) ;
mux_tree_tapbuf_size3 mux_right_track_8 (
    .in ( { chany_top_in[3] , right_top_grid_pin_42_[0] , 
        right_bottom_grid_pin_1_[0] } ) ,
    .sram ( mux_tree_tapbuf_size3_0_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size3_0_sram_inv ) , 
    .out ( chanx_right_out[4] ) , .p0 ( optlc_net_81 ) ) ;
mux_tree_tapbuf_size3_0 mux_right_track_24 (
    .in ( { chany_top_in[11] , right_top_grid_pin_42_[0] , 
        right_bottom_grid_pin_1_[0] } ) ,
    .sram ( mux_tree_tapbuf_size3_1_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size3_1_sram_inv ) , 
    .out ( chanx_right_out[12] ) , .p0 ( optlc_net_81 ) ) ;
mux_tree_tapbuf_size3_mem mem_right_track_8 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size5_mem_1_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size3_mem_0_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size3_0_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size3_0_sram_inv ) ) ;
mux_tree_tapbuf_size3_mem_0 mem_right_track_24 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_10_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size3_mem_1_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size3_1_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size3_1_sram_inv ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_1__0 ( .A ( chany_top_in[13] ) , 
    .X ( ropt_net_98 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_698 ( .A ( ropt_net_102 ) , 
    .X ( chany_top_out[6] ) ) ;
sky130_fd_sc_hd__conb_1 optlc_77 ( .LO ( SYNOPSYS_UNCONNECTED_1 ) , 
    .HI ( optlc_net_79 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_699 ( .A ( ropt_net_103 ) , 
    .X ( chany_top_out[11] ) ) ;
sky130_fd_sc_hd__conb_1 optlc_79 ( .LO ( SYNOPSYS_UNCONNECTED_2 ) , 
    .HI ( optlc_net_80 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_6__5 ( .A ( chany_top_in[18] ) , 
    .X ( ropt_net_101 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_7__6 ( .A ( chanx_right_in[0] ) , 
    .X ( ropt_net_95 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_81 ( .LO ( SYNOPSYS_UNCONNECTED_3 ) , 
    .HI ( optlc_net_81 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_83 ( .LO ( SYNOPSYS_UNCONNECTED_4 ) , 
    .HI ( optlc_net_82 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_10__9 ( .A ( chanx_right_in[6] ) , 
    .X ( ropt_net_97 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_672 ( .A ( ropt_net_83 ) , 
    .X ( ccff_tail[0] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_673 ( .A ( chanx_right_in[17] ) , 
    .X ( ropt_net_108 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_700 ( .A ( ropt_net_104 ) , 
    .X ( chany_top_out[9] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_674 ( .A ( chanx_right_in[2] ) , 
    .X ( ropt_net_110 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_675 ( .A ( chany_top_in[14] ) , 
    .X ( ropt_net_109 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_16__15 ( .A ( chanx_right_in[12] ) , 
    .X ( ropt_net_100 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_676 ( .A ( chany_top_in[17] ) , 
    .X ( ropt_net_112 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_18__17 ( .A ( chanx_right_in[15] ) , 
    .X ( ropt_net_92 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_677 ( .A ( chany_top_in[16] ) , 
    .X ( ropt_net_111 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_701 ( .A ( ropt_net_105 ) , 
    .X ( chanx_right_out[19] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_678 ( .A ( ropt_net_89 ) , 
    .X ( ropt_net_106 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_22__21 ( .A ( chanx_right_in[19] ) , 
    .X ( chany_top_out[18] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_RR_42 ( .A ( chany_top_in[15] ) , 
    .X ( ropt_net_90 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_702 ( .A ( ropt_net_106 ) , 
    .X ( chany_top_out[17] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_RR_44 ( .A ( chanx_right_in[4] ) , 
    .X ( ropt_net_93 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_45 ( .A ( chanx_right_in[7] ) , 
    .X ( ropt_net_94 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_46 ( .A ( chanx_right_in[8] ) , 
    .X ( BUF_net_46 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_47 ( .A ( chanx_right_in[9] ) , 
    .X ( BUF_net_47 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_48 ( .A ( chanx_right_in[10] ) , 
    .X ( ropt_net_99 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_49 ( .A ( chanx_right_in[14] ) , 
    .X ( BUF_net_49 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_679 ( .A ( ropt_net_90 ) , 
    .X ( chanx_right_out[16] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_51 ( .A ( chanx_right_in[18] ) , 
    .X ( ropt_net_89 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_680 ( .A ( ropt_net_91 ) , 
    .X ( chany_top_out[12] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_681 ( .A ( ropt_net_92 ) , 
    .X ( chany_top_out[14] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_682 ( .A ( ropt_net_93 ) , 
    .X ( chany_top_out[3] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_683 ( .A ( ropt_net_94 ) , 
    .X ( ropt_net_102 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_684 ( .A ( ropt_net_95 ) , 
    .X ( chany_top_out[19] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_703 ( .A ( ropt_net_107 ) , 
    .X ( chany_top_out[5] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_P_64 ( .A ( chanx_right_in[11] ) , 
    .X ( ropt_net_96 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_P_65 ( .A ( chanx_right_in[16] ) , 
    .X ( chany_top_out[15] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 BUFT_P_66 ( .A ( BUF_net_47 ) , 
    .X ( chany_top_out[8] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_705 ( .A ( ropt_net_108 ) , 
    .X ( chany_top_out[16] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_706 ( .A ( ropt_net_109 ) , 
    .X ( chanx_right_out[15] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_685 ( .A ( ropt_net_96 ) , 
    .X ( chany_top_out[10] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 BUFT_P_71 ( .A ( BUF_net_46 ) , 
    .X ( chany_top_out[7] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 BUFT_P_72 ( .A ( BUF_net_49 ) , 
    .X ( chany_top_out[13] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_686 ( .A ( ropt_net_97 ) , 
    .X ( ropt_net_107 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_687 ( .A ( ropt_net_98 ) , 
    .X ( chanx_right_out[14] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_688 ( .A ( ropt_net_99 ) , 
    .X ( ropt_net_104 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_689 ( .A ( ropt_net_100 ) , 
    .X ( ropt_net_103 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_690 ( .A ( ropt_net_101 ) , 
    .X ( ropt_net_105 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_707 ( .A ( ropt_net_110 ) , 
    .X ( chany_top_out[1] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_708 ( .A ( ropt_net_111 ) , 
    .X ( chanx_right_out[17] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_709 ( .A ( ropt_net_112 ) , 
    .X ( chanx_right_out[18] ) ) ;
endmodule


module direct_interc_4 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

assign out[0] = in[0] ;
endmodule


module GPIO_sky130_fd_sc_hd__dfxbp_1_mem_3 ( prog_clk , ccff_head , 
    ccff_tail , mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:0] mem_out ;
output [0:0] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( \_gOb0_mem_outb[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_2__2 ( .A ( mem_out[0] ) , 
    .X ( net_aps_2 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_10 ( .A ( net_aps_2 ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module GPIO_3 ( A , IE , OE , Y , in , out , mem_out ) ;
output A ;
output IE ;
output OE ;
output Y ;
input  in ;
output out ;
input  mem_out ;

assign A = in ;
assign out = Y ;

sky130_fd_sc_hd__inv_1 ie_oe_inv ( .A ( BUF_net_7 ) , .Y ( OE ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 FTB_1__1 ( .A ( mem_out ) , .X ( IE ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_7 ( .A ( IE ) , .X ( BUF_net_7 ) ) ;
endmodule


module logical_tile_io_mode_physical__iopad_3 ( prog_clk , gfpga_pad_GPIO_A , 
    gfpga_pad_GPIO_IE , gfpga_pad_GPIO_OE , gfpga_pad_GPIO_Y , iopad_outpad , 
    ccff_head , iopad_inpad , ccff_tail ) ;
input  [0:0] prog_clk ;
output [0:0] gfpga_pad_GPIO_A ;
output [0:0] gfpga_pad_GPIO_IE ;
output [0:0] gfpga_pad_GPIO_OE ;
inout  [0:0] gfpga_pad_GPIO_Y ;
input  [0:0] iopad_outpad ;
input  [0:0] ccff_head ;
output [0:0] iopad_inpad ;
output [0:0] ccff_tail ;

wire [0:0] GPIO_0_en ;

GPIO_3 GPIO_0_ ( .A ( gfpga_pad_GPIO_A[0] ) , .IE ( gfpga_pad_GPIO_IE[0] ) , 
    .OE ( gfpga_pad_GPIO_OE[0] ) , .Y ( gfpga_pad_GPIO_Y[0] ) , 
    .in ( iopad_outpad[0] ) , .out ( iopad_inpad[0] ) , 
    .mem_out ( GPIO_0_en[0] ) ) ;
GPIO_sky130_fd_sc_hd__dfxbp_1_mem_3 GPIO_sky130_fd_sc_hd__dfxbp_1_mem ( 
    .prog_clk ( prog_clk ) , .ccff_head ( ccff_head ) , 
    .ccff_tail ( ccff_tail ) , .mem_out ( GPIO_0_en ) ,
    .mem_outb ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
endmodule


module logical_tile_io_mode_io__3 ( prog_clk , gfpga_pad_GPIO_A , 
    gfpga_pad_GPIO_IE , gfpga_pad_GPIO_OE , gfpga_pad_GPIO_Y , io_outpad , 
    ccff_head , io_inpad , ccff_tail ) ;
input  [0:0] prog_clk ;
output [0:0] gfpga_pad_GPIO_A ;
output [0:0] gfpga_pad_GPIO_IE ;
output [0:0] gfpga_pad_GPIO_OE ;
inout  [0:0] gfpga_pad_GPIO_Y ;
input  [0:0] io_outpad ;
input  [0:0] ccff_head ;
output [0:0] io_inpad ;
output [0:0] ccff_tail ;

logical_tile_io_mode_physical__iopad_3 logical_tile_io_mode_physical__iopad_0 ( 
    .prog_clk ( prog_clk ) , .gfpga_pad_GPIO_A ( gfpga_pad_GPIO_A ) , 
    .gfpga_pad_GPIO_IE ( gfpga_pad_GPIO_IE ) , 
    .gfpga_pad_GPIO_OE ( gfpga_pad_GPIO_OE ) , 
    .gfpga_pad_GPIO_Y ( gfpga_pad_GPIO_Y ) , .iopad_outpad ( io_outpad ) , 
    .ccff_head ( ccff_head ) , .iopad_inpad ( io_inpad ) , 
    .ccff_tail ( ccff_tail ) ) ;
direct_interc_4 direct_interc_0_ (
    .in ( { SYNOPSYS_UNCONNECTED_1 } ) ,
    .out ( io_inpad ) ) ;
direct_interc_4 direct_interc_1_ (
    .in ( { SYNOPSYS_UNCONNECTED_2 } ) ,
    .out ( io_outpad ) ) ;
endmodule


module grid_io_left ( prog_clk , gfpga_pad_GPIO_A , gfpga_pad_GPIO_IE , 
    gfpga_pad_GPIO_OE , gfpga_pad_GPIO_Y , right_width_0_height_0__pin_0_ , 
    ccff_head , right_width_0_height_0__pin_1_upper , 
    right_width_0_height_0__pin_1_lower , ccff_tail ) ;
input  [0:0] prog_clk ;
output [0:0] gfpga_pad_GPIO_A ;
output [0:0] gfpga_pad_GPIO_IE ;
output [0:0] gfpga_pad_GPIO_OE ;
inout  [0:0] gfpga_pad_GPIO_Y ;
input  [0:0] right_width_0_height_0__pin_0_ ;
input  [0:0] ccff_head ;
output [0:0] right_width_0_height_0__pin_1_upper ;
output [0:0] right_width_0_height_0__pin_1_lower ;
output [0:0] ccff_tail ;

logical_tile_io_mode_io__3 logical_tile_io_mode_io__0 ( 
    .prog_clk ( prog_clk ) , .gfpga_pad_GPIO_A ( gfpga_pad_GPIO_A ) ,
    .gfpga_pad_GPIO_IE ( { ropt_net_14 } ) ,
    .gfpga_pad_GPIO_OE ( gfpga_pad_GPIO_OE ) , 
    .gfpga_pad_GPIO_Y ( gfpga_pad_GPIO_Y ) , 
    .io_outpad ( right_width_0_height_0__pin_0_ ) , .ccff_head ( ccff_head ) , 
    .io_inpad ( right_width_0_height_0__pin_1_upper ) ,
    .ccff_tail ( { ropt_net_15 } ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_1__0 ( 
    .A ( right_width_0_height_0__pin_1_upper[0] ) , 
    .X ( right_width_0_height_0__pin_1_lower[0] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_573 ( .A ( ropt_net_14 ) , 
    .X ( gfpga_pad_GPIO_IE[0] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_574 ( .A ( ropt_net_15 ) , 
    .X ( ropt_net_16 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_575 ( .A ( ropt_net_16 ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module direct_interc_3 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

assign out[0] = in[0] ;
endmodule


module GPIO_sky130_fd_sc_hd__dfxbp_1_mem_2 ( prog_clk , ccff_head , 
    ccff_tail , mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:0] mem_out ;
output [0:0] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( \_gOb0_mem_outb[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_2__2 ( .A ( mem_out[0] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module GPIO_2 ( A , IE , OE , Y , in , out , mem_out ) ;
output A ;
output IE ;
output OE ;
output Y ;
input  in ;
output out ;
input  mem_out ;

wire aps_rename_1_ ;

assign A = in ;
assign out = Y ;

sky130_fd_sc_hd__inv_1 ie_oe_inv ( .A ( aps_rename_1_ ) , .Y ( OE ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_1__1 ( .A ( mem_out ) , 
    .X ( aps_rename_1_ ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_5 ( .A ( aps_rename_1_ ) , .X ( IE ) ) ;
endmodule


module logical_tile_io_mode_physical__iopad_2 ( prog_clk , gfpga_pad_GPIO_A , 
    gfpga_pad_GPIO_IE , gfpga_pad_GPIO_OE , gfpga_pad_GPIO_Y , iopad_outpad , 
    ccff_head , iopad_inpad , ccff_tail ) ;
input  [0:0] prog_clk ;
output [0:0] gfpga_pad_GPIO_A ;
output [0:0] gfpga_pad_GPIO_IE ;
output [0:0] gfpga_pad_GPIO_OE ;
inout  [0:0] gfpga_pad_GPIO_Y ;
input  [0:0] iopad_outpad ;
input  [0:0] ccff_head ;
output [0:0] iopad_inpad ;
output [0:0] ccff_tail ;

wire [0:0] GPIO_0_en ;

GPIO_2 GPIO_0_ ( .A ( gfpga_pad_GPIO_A[0] ) , .IE ( gfpga_pad_GPIO_IE[0] ) , 
    .OE ( gfpga_pad_GPIO_OE[0] ) , .Y ( gfpga_pad_GPIO_Y[0] ) , 
    .in ( iopad_outpad[0] ) , .out ( iopad_inpad[0] ) , 
    .mem_out ( GPIO_0_en[0] ) ) ;
GPIO_sky130_fd_sc_hd__dfxbp_1_mem_2 GPIO_sky130_fd_sc_hd__dfxbp_1_mem ( 
    .prog_clk ( prog_clk ) , .ccff_head ( ccff_head ) , 
    .ccff_tail ( ccff_tail ) , .mem_out ( GPIO_0_en ) ,
    .mem_outb ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
endmodule


module logical_tile_io_mode_io__2 ( prog_clk , gfpga_pad_GPIO_A , 
    gfpga_pad_GPIO_IE , gfpga_pad_GPIO_OE , gfpga_pad_GPIO_Y , io_outpad , 
    ccff_head , io_inpad , ccff_tail ) ;
input  [0:0] prog_clk ;
output [0:0] gfpga_pad_GPIO_A ;
output [0:0] gfpga_pad_GPIO_IE ;
output [0:0] gfpga_pad_GPIO_OE ;
inout  [0:0] gfpga_pad_GPIO_Y ;
input  [0:0] io_outpad ;
input  [0:0] ccff_head ;
output [0:0] io_inpad ;
output [0:0] ccff_tail ;

logical_tile_io_mode_physical__iopad_2 logical_tile_io_mode_physical__iopad_0 ( 
    .prog_clk ( prog_clk ) , .gfpga_pad_GPIO_A ( gfpga_pad_GPIO_A ) , 
    .gfpga_pad_GPIO_IE ( gfpga_pad_GPIO_IE ) , 
    .gfpga_pad_GPIO_OE ( gfpga_pad_GPIO_OE ) , 
    .gfpga_pad_GPIO_Y ( gfpga_pad_GPIO_Y ) , .iopad_outpad ( io_outpad ) , 
    .ccff_head ( ccff_head ) , .iopad_inpad ( io_inpad ) , 
    .ccff_tail ( ccff_tail ) ) ;
direct_interc_3 direct_interc_0_ (
    .in ( { SYNOPSYS_UNCONNECTED_1 } ) ,
    .out ( io_inpad ) ) ;
direct_interc_3 direct_interc_1_ (
    .in ( { SYNOPSYS_UNCONNECTED_2 } ) ,
    .out ( io_outpad ) ) ;
endmodule


module grid_io_bottom ( prog_clk , gfpga_pad_GPIO_A , gfpga_pad_GPIO_IE , 
    gfpga_pad_GPIO_OE , gfpga_pad_GPIO_Y , top_width_0_height_0__pin_0_ , 
    ccff_head , top_width_0_height_0__pin_1_upper , 
    top_width_0_height_0__pin_1_lower , ccff_tail ) ;
input  [0:0] prog_clk ;
output [0:0] gfpga_pad_GPIO_A ;
output [0:0] gfpga_pad_GPIO_IE ;
output [0:0] gfpga_pad_GPIO_OE ;
inout  [0:0] gfpga_pad_GPIO_Y ;
input  [0:0] top_width_0_height_0__pin_0_ ;
input  [0:0] ccff_head ;
output [0:0] top_width_0_height_0__pin_1_upper ;
output [0:0] top_width_0_height_0__pin_1_lower ;
output [0:0] ccff_tail ;

logical_tile_io_mode_io__2 logical_tile_io_mode_io__0 ( 
    .prog_clk ( prog_clk ) , .gfpga_pad_GPIO_A ( gfpga_pad_GPIO_A ) ,
    .gfpga_pad_GPIO_IE ( { ropt_net_14 } ) ,
    .gfpga_pad_GPIO_OE ( gfpga_pad_GPIO_OE ) , 
    .gfpga_pad_GPIO_Y ( gfpga_pad_GPIO_Y ) , 
    .io_outpad ( top_width_0_height_0__pin_0_ ) , .ccff_head ( ccff_head ) , 
    .io_inpad ( top_width_0_height_0__pin_1_upper ) ,
    .ccff_tail ( { ropt_net_15 } ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_1__0 ( 
    .A ( top_width_0_height_0__pin_1_upper[0] ) , .X ( aps_rename_2_ ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_573 ( .A ( ropt_net_14 ) , 
    .X ( ropt_net_17 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 BUFT_RR_8 ( .A ( aps_rename_2_ ) , 
    .X ( top_width_0_height_0__pin_1_lower[0] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_574 ( .A ( ropt_net_15 ) , 
    .X ( ccff_tail[0] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_575 ( .A ( ropt_net_17 ) , 
    .X ( gfpga_pad_GPIO_IE[0] ) ) ;
endmodule


module direct_interc_2 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

assign out[0] = in[0] ;
endmodule


module GPIO_sky130_fd_sc_hd__dfxbp_1_mem_1 ( prog_clk , ccff_head , 
    ccff_tail , mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:0] mem_out ;
output [0:0] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( \_gOb0_mem_outb[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_2__2 ( .A ( mem_out[0] ) , 
    .X ( net_net_7 ) ) ;
sky130_fd_sc_hd__dlygate4sd1_1 BUFT_RR_7 ( .A ( net_net_7 ) , 
    .X ( net_net_6 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_RR_9 ( .A ( net_net_6 ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module GPIO_1 ( A , IE , OE , Y , in , out , mem_out ) ;
output A ;
output IE ;
output OE ;
output Y ;
input  in ;
output out ;
input  mem_out ;

wire aps_rename_1_ ;

assign A = in ;
assign out = Y ;

sky130_fd_sc_hd__inv_1 ie_oe_inv ( .A ( IE ) , .Y ( OE ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_1__1 ( .A ( mem_out ) , 
    .X ( aps_rename_1_ ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 BUFT_RR_3 ( .A ( aps_rename_1_ ) , .X ( IE ) ) ;
endmodule


module logical_tile_io_mode_physical__iopad_1 ( prog_clk , gfpga_pad_GPIO_A , 
    gfpga_pad_GPIO_IE , gfpga_pad_GPIO_OE , gfpga_pad_GPIO_Y , iopad_outpad , 
    ccff_head , iopad_inpad , ccff_tail ) ;
input  [0:0] prog_clk ;
output [0:0] gfpga_pad_GPIO_A ;
output [0:0] gfpga_pad_GPIO_IE ;
output [0:0] gfpga_pad_GPIO_OE ;
inout  [0:0] gfpga_pad_GPIO_Y ;
input  [0:0] iopad_outpad ;
input  [0:0] ccff_head ;
output [0:0] iopad_inpad ;
output [0:0] ccff_tail ;

wire [0:0] GPIO_0_en ;

GPIO_1 GPIO_0_ ( .A ( gfpga_pad_GPIO_A[0] ) , .IE ( gfpga_pad_GPIO_IE[0] ) , 
    .OE ( gfpga_pad_GPIO_OE[0] ) , .Y ( gfpga_pad_GPIO_Y[0] ) , 
    .in ( iopad_outpad[0] ) , .out ( iopad_inpad[0] ) , 
    .mem_out ( GPIO_0_en[0] ) ) ;
GPIO_sky130_fd_sc_hd__dfxbp_1_mem_1 GPIO_sky130_fd_sc_hd__dfxbp_1_mem ( 
    .prog_clk ( prog_clk ) , .ccff_head ( ccff_head ) , 
    .ccff_tail ( ccff_tail ) , .mem_out ( GPIO_0_en ) ,
    .mem_outb ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
endmodule


module logical_tile_io_mode_io__1 ( prog_clk , gfpga_pad_GPIO_A , 
    gfpga_pad_GPIO_IE , gfpga_pad_GPIO_OE , gfpga_pad_GPIO_Y , io_outpad , 
    ccff_head , io_inpad , ccff_tail ) ;
input  [0:0] prog_clk ;
output [0:0] gfpga_pad_GPIO_A ;
output [0:0] gfpga_pad_GPIO_IE ;
output [0:0] gfpga_pad_GPIO_OE ;
inout  [0:0] gfpga_pad_GPIO_Y ;
input  [0:0] io_outpad ;
input  [0:0] ccff_head ;
output [0:0] io_inpad ;
output [0:0] ccff_tail ;

logical_tile_io_mode_physical__iopad_1 logical_tile_io_mode_physical__iopad_0 ( 
    .prog_clk ( prog_clk ) , .gfpga_pad_GPIO_A ( gfpga_pad_GPIO_A ) , 
    .gfpga_pad_GPIO_IE ( gfpga_pad_GPIO_IE ) , 
    .gfpga_pad_GPIO_OE ( gfpga_pad_GPIO_OE ) , 
    .gfpga_pad_GPIO_Y ( gfpga_pad_GPIO_Y ) , .iopad_outpad ( io_outpad ) , 
    .ccff_head ( ccff_head ) , .iopad_inpad ( io_inpad ) , 
    .ccff_tail ( ccff_tail ) ) ;
direct_interc_2 direct_interc_0_ (
    .in ( { SYNOPSYS_UNCONNECTED_1 } ) ,
    .out ( io_inpad ) ) ;
direct_interc_2 direct_interc_1_ (
    .in ( { SYNOPSYS_UNCONNECTED_2 } ) ,
    .out ( io_outpad ) ) ;
endmodule


module grid_io_right ( prog_clk , gfpga_pad_GPIO_A , gfpga_pad_GPIO_IE , 
    gfpga_pad_GPIO_OE , gfpga_pad_GPIO_Y , left_width_0_height_0__pin_0_ , 
    ccff_head , left_width_0_height_0__pin_1_upper , 
    left_width_0_height_0__pin_1_lower , ccff_tail ) ;
input  [0:0] prog_clk ;
output [0:0] gfpga_pad_GPIO_A ;
output [0:0] gfpga_pad_GPIO_IE ;
output [0:0] gfpga_pad_GPIO_OE ;
inout  [0:0] gfpga_pad_GPIO_Y ;
input  [0:0] left_width_0_height_0__pin_0_ ;
input  [0:0] ccff_head ;
output [0:0] left_width_0_height_0__pin_1_upper ;
output [0:0] left_width_0_height_0__pin_1_lower ;
output [0:0] ccff_tail ;

logical_tile_io_mode_io__1 logical_tile_io_mode_io__0 ( 
    .prog_clk ( prog_clk ) , .gfpga_pad_GPIO_A ( gfpga_pad_GPIO_A ) , 
    .gfpga_pad_GPIO_IE ( gfpga_pad_GPIO_IE ) , 
    .gfpga_pad_GPIO_OE ( gfpga_pad_GPIO_OE ) , 
    .gfpga_pad_GPIO_Y ( gfpga_pad_GPIO_Y ) , 
    .io_outpad ( left_width_0_height_0__pin_0_ ) , .ccff_head ( ccff_head ) , 
    .io_inpad ( left_width_0_height_0__pin_1_upper ) ,
    .ccff_tail ( { ropt_net_14 } ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_1__0 ( 
    .A ( left_width_0_height_0__pin_1_upper[0] ) , .X ( aps_rename_2_ ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_574 ( .A ( ropt_net_15 ) , 
    .X ( left_width_0_height_0__pin_1_lower[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_P_8 ( .A ( aps_rename_2_ ) , 
    .X ( ropt_net_13 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_572 ( .A ( ropt_net_13 ) , 
    .X ( ropt_net_15 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_573 ( .A ( ropt_net_14 ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module direct_interc_1 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

assign out[0] = in[0] ;
endmodule


module GPIO_sky130_fd_sc_hd__dfxbp_1_mem ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:0] mem_out ;
output [0:0] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( \_gOb0_mem_outb[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_2__2 ( .A ( mem_out[0] ) , 
    .X ( net_net_7 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_RR_9 ( .A ( net_net_7 ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module GPIO ( A , IE , OE , Y , in , out , mem_out ) ;
output A ;
output IE ;
output OE ;
output Y ;
input  in ;
output out ;
input  mem_out ;

wire aps_rename_1_ ;

assign A = in ;
assign out = Y ;

sky130_fd_sc_hd__inv_1 ie_oe_inv ( .A ( aps_rename_1_ ) , .Y ( OE ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_1__1 ( .A ( mem_out ) , 
    .X ( aps_rename_1_ ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_4 ( .A ( aps_rename_1_ ) , .X ( IE ) ) ;
endmodule


module logical_tile_io_mode_physical__iopad ( prog_clk , gfpga_pad_GPIO_A , 
    gfpga_pad_GPIO_IE , gfpga_pad_GPIO_OE , gfpga_pad_GPIO_Y , iopad_outpad , 
    ccff_head , iopad_inpad , ccff_tail ) ;
input  [0:0] prog_clk ;
output [0:0] gfpga_pad_GPIO_A ;
output [0:0] gfpga_pad_GPIO_IE ;
output [0:0] gfpga_pad_GPIO_OE ;
inout  [0:0] gfpga_pad_GPIO_Y ;
input  [0:0] iopad_outpad ;
input  [0:0] ccff_head ;
output [0:0] iopad_inpad ;
output [0:0] ccff_tail ;

wire [0:0] GPIO_0_en ;

GPIO GPIO_0_ ( .A ( gfpga_pad_GPIO_A[0] ) , .IE ( gfpga_pad_GPIO_IE[0] ) , 
    .OE ( gfpga_pad_GPIO_OE[0] ) , .Y ( gfpga_pad_GPIO_Y[0] ) , 
    .in ( iopad_outpad[0] ) , .out ( iopad_inpad[0] ) , 
    .mem_out ( GPIO_0_en[0] ) ) ;
GPIO_sky130_fd_sc_hd__dfxbp_1_mem GPIO_sky130_fd_sc_hd__dfxbp_1_mem ( 
    .prog_clk ( prog_clk ) , .ccff_head ( ccff_head ) , 
    .ccff_tail ( ccff_tail ) , .mem_out ( GPIO_0_en ) ,
    .mem_outb ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
endmodule


module logical_tile_io_mode_io_ ( prog_clk , gfpga_pad_GPIO_A , 
    gfpga_pad_GPIO_IE , gfpga_pad_GPIO_OE , gfpga_pad_GPIO_Y , io_outpad , 
    ccff_head , io_inpad , ccff_tail ) ;
input  [0:0] prog_clk ;
output [0:0] gfpga_pad_GPIO_A ;
output [0:0] gfpga_pad_GPIO_IE ;
output [0:0] gfpga_pad_GPIO_OE ;
inout  [0:0] gfpga_pad_GPIO_Y ;
input  [0:0] io_outpad ;
input  [0:0] ccff_head ;
output [0:0] io_inpad ;
output [0:0] ccff_tail ;

logical_tile_io_mode_physical__iopad logical_tile_io_mode_physical__iopad_0 ( 
    .prog_clk ( prog_clk ) , .gfpga_pad_GPIO_A ( gfpga_pad_GPIO_A ) , 
    .gfpga_pad_GPIO_IE ( gfpga_pad_GPIO_IE ) , 
    .gfpga_pad_GPIO_OE ( gfpga_pad_GPIO_OE ) , 
    .gfpga_pad_GPIO_Y ( gfpga_pad_GPIO_Y ) , .iopad_outpad ( io_outpad ) , 
    .ccff_head ( ccff_head ) , .iopad_inpad ( io_inpad ) , 
    .ccff_tail ( ccff_tail ) ) ;
direct_interc_1 direct_interc_0_ (
    .in ( { SYNOPSYS_UNCONNECTED_1 } ) ,
    .out ( io_inpad ) ) ;
direct_interc_1 direct_interc_1_ (
    .in ( { SYNOPSYS_UNCONNECTED_2 } ) ,
    .out ( io_outpad ) ) ;
endmodule


module grid_io_top ( prog_clk , gfpga_pad_GPIO_A , gfpga_pad_GPIO_IE , 
    gfpga_pad_GPIO_OE , gfpga_pad_GPIO_Y , bottom_width_0_height_0__pin_0_ , 
    ccff_head , bottom_width_0_height_0__pin_1_upper , 
    bottom_width_0_height_0__pin_1_lower , ccff_tail ) ;
input  [0:0] prog_clk ;
output [0:0] gfpga_pad_GPIO_A ;
output [0:0] gfpga_pad_GPIO_IE ;
output [0:0] gfpga_pad_GPIO_OE ;
inout  [0:0] gfpga_pad_GPIO_Y ;
input  [0:0] bottom_width_0_height_0__pin_0_ ;
input  [0:0] ccff_head ;
output [0:0] bottom_width_0_height_0__pin_1_upper ;
output [0:0] bottom_width_0_height_0__pin_1_lower ;
output [0:0] ccff_tail ;

logical_tile_io_mode_io_ logical_tile_io_mode_io__0 ( .prog_clk ( prog_clk ) , 
    .gfpga_pad_GPIO_A ( gfpga_pad_GPIO_A ) ,
    .gfpga_pad_GPIO_IE ( { ropt_net_11 } ) ,
    .gfpga_pad_GPIO_OE ( gfpga_pad_GPIO_OE ) , 
    .gfpga_pad_GPIO_Y ( gfpga_pad_GPIO_Y ) , 
    .io_outpad ( bottom_width_0_height_0__pin_0_ ) , 
    .ccff_head ( ccff_head ) , 
    .io_inpad ( bottom_width_0_height_0__pin_1_upper ) ,
    .ccff_tail ( { ropt_net_13 } ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_1__0 ( 
    .A ( bottom_width_0_height_0__pin_1_upper[0] ) , .X ( aps_rename_2_ ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_571 ( .A ( ropt_net_11 ) , 
    .X ( ropt_net_15 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_8 ( .A ( aps_rename_2_ ) , 
    .X ( ropt_net_12 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_572 ( .A ( ropt_net_12 ) , 
    .X ( ropt_net_14 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_573 ( .A ( ropt_net_13 ) , 
    .X ( ccff_tail[0] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_574 ( .A ( ropt_net_14 ) , 
    .X ( bottom_width_0_height_0__pin_1_lower[0] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_575 ( .A ( ropt_net_15 ) , 
    .X ( gfpga_pad_GPIO_IE[0] ) ) ;
endmodule


module mux_tree_size2_mem_23 ( prog_clk , ccff_head , ccff_tail , mem_out , 
    mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_40__55 ( .A ( mem_out[1] ) , 
    .X ( net_net_88 ) ) ;
sky130_fd_sc_hd__dlygate4sd1_1 BUFT_RR_88 ( .A ( net_net_88 ) , 
    .X ( net_net_87 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 BUFT_RR_118 ( .A ( net_net_87 ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_size2_mem_22 ( prog_clk , ccff_head , ccff_tail , mem_out , 
    mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_39__54 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_size2_mem_21 ( prog_clk , ccff_head , ccff_tail , mem_out , 
    mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_38__53 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_size2_23 ( in , sram , sram_inv , out , p3 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p3 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;

const1 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p3 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , .X ( out[0] ) ) ;
endmodule


module const1_30 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_size2_22 ( in , sram , sram_inv , out , p3 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p3 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;

const1_30 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p3 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , .X ( out[0] ) ) ;
endmodule


module const1_29 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_size2_21 ( in , sram , sram_inv , out , p3 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p3 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;

const1_29 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p3 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , .X ( out[0] ) ) ;
endmodule


module logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff ( 
    Test_en , clk , ff_D , ff_DI , ff_Q , ff_clk , p_abuf1 , p_abuf2 ) ;
input  [0:0] Test_en ;
input  [0:0] clk ;
input  [0:0] ff_D ;
input  [0:0] ff_DI ;
output [0:0] ff_Q ;
input  [0:0] ff_clk ;
output p_abuf1 ;
output p_abuf2 ;

sky130_fd_sc_hd__sdfxbp_1 sky130_fd_sc_hd__sdfxbp_1_0_ ( .D ( ff_D[0] ) , 
    .SCD ( ff_DI[0] ) , .SCE ( Test_en[0] ) , .CLK ( clk[0] ) , 
    .Q ( p_abuf2 ) , .Q_N ( SYNOPSYS_UNCONNECTED_1 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_109 ( .A ( p_abuf2 ) , .X ( ff_Q[0] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 BUFT_RR_112 ( .A ( p_abuf2 ) , 
    .X ( p_abuf1 ) ) ;
endmodule


module logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_14 ( 
    Test_en , clk , ff_D , ff_DI , ff_Q , ff_clk ) ;
input  [0:0] Test_en ;
input  [0:0] clk ;
input  [0:0] ff_D ;
input  [0:0] ff_DI ;
output [0:0] ff_Q ;
input  [0:0] ff_clk ;

sky130_fd_sc_hd__sdfxbp_1 sky130_fd_sc_hd__sdfxbp_1_0_ ( .D ( ff_D[0] ) , 
    .SCD ( ff_DI[0] ) , .SCE ( Test_en[0] ) , .CLK ( clk[0] ) , 
    .Q ( ff_Q[0] ) , .Q_N ( SYNOPSYS_UNCONNECTED_1 ) ) ;
endmodule


module mux_tree_size2_mem ( prog_clk , ccff_head , ccff_tail , mem_out , 
    mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_37__52 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_28 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_size2 ( in , sram , sram_inv , out , p3 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p3 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;

const1_28 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p3 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , .X ( out[0] ) ) ;
endmodule


module frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem ( prog_clk , ccff_head , 
    ccff_tail , mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:16] mem_out ;
output [0:16] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_4_ ( .D ( mem_out[3] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[4] ) , .Q_N ( mem_outb[4] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_5_ ( .D ( mem_out[4] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[5] ) , .Q_N ( mem_outb[5] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_6_ ( .D ( mem_out[5] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[6] ) , .Q_N ( mem_outb[6] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_7_ ( .D ( mem_out[6] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[7] ) , .Q_N ( mem_outb[7] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_8_ ( .D ( mem_out[7] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[8] ) , .Q_N ( mem_outb[8] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_9_ ( .D ( mem_out[8] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[9] ) , .Q_N ( mem_outb[9] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_10_ ( .D ( mem_out[9] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[10] ) , .Q_N ( mem_outb[10] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_11_ ( .D ( mem_out[10] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[11] ) , .Q_N ( mem_outb[11] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_12_ ( .D ( mem_out[11] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[12] ) , .Q_N ( mem_outb[12] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_13_ ( .D ( mem_out[12] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[13] ) , .Q_N ( mem_outb[13] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_14_ ( .D ( mem_out[13] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[14] ) , .Q_N ( mem_outb[14] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_15_ ( .D ( mem_out[14] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[15] ) , .Q_N ( mem_outb[15] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_16_ ( .D ( mem_out[15] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[16] ) , .Q_N ( \_gOb7_mem_outb[16] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_36__51 ( .A ( mem_out[16] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module frac_lut4_mux ( in , sram , sram_inv , lut3_out , lut4_out ) ;
input  [0:15] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:1] lut3_out ;
output [0:0] lut4_out ;

wire [0:0] sky130_fd_sc_hd__buf_2_3_X ;
wire [0:0] sky130_fd_sc_hd__buf_2_4_X ;
wire [0:0] sky130_fd_sc_hd__buf_2_5_X ;
wire [0:0] sky130_fd_sc_hd__buf_2_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_10_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_11_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_12_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_13_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_14_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_12_X[0] ) , .X ( lut3_out[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_1_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_13_X[0] ) , .X ( lut3_out[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_2_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_14_X[0] ) , .X ( lut4_out[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_3_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .X ( sky130_fd_sc_hd__buf_2_3_X[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_4_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , 
    .X ( sky130_fd_sc_hd__buf_2_4_X[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_5_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_10_X[0] ) , 
    .X ( sky130_fd_sc_hd__buf_2_5_X[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_6_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_11_X[0] ) , 
    .X ( sky130_fd_sc_hd__buf_2_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_3_ ( .A0 ( in[7] ) , .A1 ( in[6] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_4_ ( .A0 ( in[9] ) , .A1 ( in[8] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_5_ ( .A0 ( in[11] ) , .A1 ( in[10] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_6_ ( .A0 ( in[13] ) , .A1 ( in[12] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_7_ ( .A0 ( in[15] ) , .A1 ( in[14] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_10_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_11_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( .A0 ( sky130_fd_sc_hd__buf_2_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__buf_2_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_12_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( .A0 ( sky130_fd_sc_hd__buf_2_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__buf_2_5_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_13_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_13_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_12_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_14_X[0] ) ) ;
endmodule


module frac_lut4 ( in , sram , sram_inv , mode , mode_inv , lut3_out , 
    lut4_out ) ;
input  [0:3] in ;
input  [0:15] sram ;
input  [0:15] sram_inv ;
input  [0:0] mode ;
input  [0:0] mode_inv ;
output [0:1] lut3_out ;
output [0:0] lut4_out ;

wire [0:0] sky130_fd_sc_hd__buf_2_0_X ;
wire [0:0] sky130_fd_sc_hd__buf_2_1_X ;
wire [0:0] sky130_fd_sc_hd__buf_2_2_X ;
wire [0:0] sky130_fd_sc_hd__buf_2_3_X ;
wire [0:0] sky130_fd_sc_hd__inv_1_0_Y ;
wire [0:0] sky130_fd_sc_hd__inv_1_1_Y ;
wire [0:0] sky130_fd_sc_hd__inv_1_2_Y ;
wire [0:0] sky130_fd_sc_hd__inv_1_3_Y ;
wire [0:0] sky130_fd_sc_hd__or2_1_0_X ;

sky130_fd_sc_hd__or2_0 sky130_fd_sc_hd__or2_1_0_ ( .A ( mode[0] ) , 
    .B ( in[3] ) , .X ( sky130_fd_sc_hd__or2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__inv_1 sky130_fd_sc_hd__inv_1_0_ ( .A ( in[0] ) , 
    .Y ( sky130_fd_sc_hd__inv_1_0_Y[0] ) ) ;
sky130_fd_sc_hd__inv_1 sky130_fd_sc_hd__inv_1_1_ ( .A ( in[1] ) , 
    .Y ( sky130_fd_sc_hd__inv_1_1_Y[0] ) ) ;
sky130_fd_sc_hd__inv_1 sky130_fd_sc_hd__inv_1_2_ ( .A ( in[2] ) , 
    .Y ( sky130_fd_sc_hd__inv_1_2_Y[0] ) ) ;
sky130_fd_sc_hd__inv_1 sky130_fd_sc_hd__inv_1_3_ ( 
    .A ( sky130_fd_sc_hd__or2_1_0_X[0] ) , 
    .Y ( sky130_fd_sc_hd__inv_1_3_Y[0] ) ) ;
sky130_fd_sc_hd__buf_2 sky130_fd_sc_hd__buf_2_0_ ( .A ( in[0] ) , 
    .X ( sky130_fd_sc_hd__buf_2_0_X[0] ) ) ;
sky130_fd_sc_hd__buf_2 sky130_fd_sc_hd__buf_2_1_ ( .A ( in[1] ) , 
    .X ( sky130_fd_sc_hd__buf_2_1_X[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_2_ ( .A ( in[2] ) , 
    .X ( sky130_fd_sc_hd__buf_2_2_X[0] ) ) ;
sky130_fd_sc_hd__buf_2 sky130_fd_sc_hd__buf_2_3_ ( 
    .A ( sky130_fd_sc_hd__or2_1_0_X[0] ) , 
    .X ( sky130_fd_sc_hd__buf_2_3_X[0] ) ) ;
frac_lut4_mux frac_lut4_mux_0_ ( .in ( sram ) ,
    .sram ( { sky130_fd_sc_hd__buf_2_0_X[0] , sky130_fd_sc_hd__buf_2_1_X[0] , 
        sky130_fd_sc_hd__buf_2_2_X[0] , sky130_fd_sc_hd__buf_2_3_X[0] } ) ,
    .sram_inv ( { sky130_fd_sc_hd__inv_1_0_Y[0] , 
        sky130_fd_sc_hd__inv_1_1_Y[0] , sky130_fd_sc_hd__inv_1_2_Y[0] , 
        sky130_fd_sc_hd__inv_1_3_Y[0] } ) ,
    .lut3_out ( lut3_out ) , .lut4_out ( lut4_out ) ) ;
endmodule


module logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4 ( 
    prog_clk , frac_lut4_in , ccff_head , frac_lut4_lut3_out , 
    frac_lut4_lut4_out , ccff_tail ) ;
input  [0:0] prog_clk ;
input  [0:3] frac_lut4_in ;
input  [0:0] ccff_head ;
output [0:1] frac_lut4_lut3_out ;
output [0:0] frac_lut4_lut4_out ;
output [0:0] ccff_tail ;

wire [0:0] frac_lut4_0_mode ;
wire [0:15] frac_lut4_0_sram ;
wire [0:15] frac_lut4_0_sram_inv ;

frac_lut4 frac_lut4_0_ ( .in ( frac_lut4_in ) , .sram ( frac_lut4_0_sram ) , 
    .sram_inv ( frac_lut4_0_sram_inv ) , .mode ( frac_lut4_0_mode ) ,
    .mode_inv ( { SYNOPSYS_UNCONNECTED_1 } ) ,
    .lut3_out ( frac_lut4_lut3_out ) , .lut4_out ( frac_lut4_lut4_out ) ) ;
frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem ( 
    .prog_clk ( prog_clk ) , .ccff_head ( ccff_head ) , 
    .ccff_tail ( ccff_tail ) ,
    .mem_out ( { frac_lut4_0_sram[0] , frac_lut4_0_sram[1] , 
        frac_lut4_0_sram[2] , frac_lut4_0_sram[3] , frac_lut4_0_sram[4] , 
        frac_lut4_0_sram[5] , frac_lut4_0_sram[6] , frac_lut4_0_sram[7] , 
        frac_lut4_0_sram[8] , frac_lut4_0_sram[9] , frac_lut4_0_sram[10] , 
        frac_lut4_0_sram[11] , frac_lut4_0_sram[12] , frac_lut4_0_sram[13] , 
        frac_lut4_0_sram[14] , frac_lut4_0_sram[15] , frac_lut4_0_mode[0] } ) ,
    .mem_outb ( { frac_lut4_0_sram_inv[0] , frac_lut4_0_sram_inv[1] , 
        frac_lut4_0_sram_inv[2] , frac_lut4_0_sram_inv[3] , 
        frac_lut4_0_sram_inv[4] , frac_lut4_0_sram_inv[5] , 
        frac_lut4_0_sram_inv[6] , frac_lut4_0_sram_inv[7] , 
        frac_lut4_0_sram_inv[8] , frac_lut4_0_sram_inv[9] , 
        frac_lut4_0_sram_inv[10] , frac_lut4_0_sram_inv[11] , 
        frac_lut4_0_sram_inv[12] , frac_lut4_0_sram_inv[13] , 
        frac_lut4_0_sram_inv[14] , frac_lut4_0_sram_inv[15] , 
        SYNOPSYS_UNCONNECTED_2 } ) ) ;
endmodule


module logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic ( 
    prog_clk , frac_logic_in , ccff_head , frac_logic_out , ccff_tail , p3 ) ;
input  [0:0] prog_clk ;
input  [0:3] frac_logic_in ;
input  [0:0] ccff_head ;
output [0:1] frac_logic_out ;
output [0:0] ccff_tail ;
input  p3 ;

wire [0:0] logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_ccff_tail ;
wire [0:0] logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_frac_lut4_lut3_out ;
wire [0:0] logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_frac_lut4_lut4_out ;
wire [0:1] mux_tree_size2_0_sram ;
wire [0:1] mux_tree_size2_0_sram_inv ;

logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4 logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0 ( 
    .prog_clk ( prog_clk ) , .frac_lut4_in ( frac_logic_in ) , 
    .ccff_head ( ccff_head ) ,
    .frac_lut4_lut3_out ( { 
        logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_frac_lut4_lut3_out[0] , 
        frac_logic_out[1] } ) ,
    
    .frac_lut4_lut4_out ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_frac_lut4_lut4_out ) , 
    .ccff_tail ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_ccff_tail ) ) ;
mux_tree_size2 mux_frac_logic_out_0 (
    .in ( { 
        logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_frac_lut4_lut4_out[0] , 
        logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_frac_lut4_lut3_out[0]
         } ) ,
    .sram ( mux_tree_size2_0_sram ) , 
    .sram_inv ( mux_tree_size2_0_sram_inv ) , .out ( frac_logic_out[0] ) , 
    .p3 ( p3 ) ) ;
mux_tree_size2_mem mem_frac_logic_out_0 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_ccff_tail ) , 
    .ccff_tail ( ccff_tail ) , .mem_out ( mux_tree_size2_0_sram ) , 
    .mem_outb ( mux_tree_size2_0_sram_inv ) ) ;
direct_interc direct_interc_0_ (
    .in ( { SYNOPSYS_UNCONNECTED_1 } ) ,
    .out ( frac_logic_out[1] ) ) ;
direct_interc direct_interc_1_ (
    .in ( { SYNOPSYS_UNCONNECTED_2 } ) ,
    .out ( frac_logic_in[0] ) ) ;
direct_interc direct_interc_2_ (
    .in ( { SYNOPSYS_UNCONNECTED_3 } ) ,
    .out ( frac_logic_in[1] ) ) ;
direct_interc direct_interc_3_ (
    .in ( { SYNOPSYS_UNCONNECTED_4 } ) ,
    .out ( frac_logic_in[2] ) ) ;
direct_interc direct_interc_4_ (
    .in ( { SYNOPSYS_UNCONNECTED_5 } ) ,
    .out ( frac_logic_in[3] ) ) ;
endmodule


module logical_tile_clb_mode_default__fle_mode_physical__fabric ( prog_clk , 
    Test_en , clk , fabric_in , fabric_regin , fabric_scin , fabric_clk , 
    ccff_head , fabric_out , fabric_regout , fabric_scout , ccff_tail , 
    p_abuf1 , p_abuf2 , p3 ) ;
input  [0:0] prog_clk ;
input  [0:0] Test_en ;
input  [0:0] clk ;
input  [0:3] fabric_in ;
input  [0:0] fabric_regin ;
input  [0:0] fabric_scin ;
input  [0:0] fabric_clk ;
input  [0:0] ccff_head ;
output [0:1] fabric_out ;
output [0:0] fabric_regout ;
output [0:0] fabric_scout ;
output [0:0] ccff_tail ;
output p_abuf1 ;
output p_abuf2 ;
input  p3 ;

wire [0:0] logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1_ff_Q ;
wire [0:0] logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0_ff_Q ;
wire [0:0] logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_ccff_tail ;
wire [0:1] logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_frac_logic_out ;
wire [0:1] mux_tree_size2_0_sram ;
wire [0:1] mux_tree_size2_0_sram_inv ;
wire [0:1] mux_tree_size2_1_sram ;
wire [0:1] mux_tree_size2_1_sram_inv ;
wire [0:0] mux_tree_size2_2_out ;
wire [0:1] mux_tree_size2_2_sram ;
wire [0:1] mux_tree_size2_2_sram_inv ;
wire [0:0] mux_tree_size2_mem_0_ccff_tail ;
wire [0:0] mux_tree_size2_mem_1_ccff_tail ;

assign p_abuf1 = p_abuf2 ;

logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0 ( 
    .prog_clk ( prog_clk ) , .frac_logic_in ( fabric_in ) , 
    .ccff_head ( ccff_head ) , 
    .frac_logic_out ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_frac_logic_out ) , 
    .ccff_tail ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_ccff_tail ) , 
    .p3 ( p3 ) ) ;
logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_14 logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0 ( 
    .Test_en ( Test_en ) , .clk ( clk ) , .ff_D ( mux_tree_size2_2_out ) , 
    .ff_DI ( fabric_scin ) , 
    .ff_Q ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0_ff_Q ) ,
    .ff_clk ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1 ( 
    .Test_en ( Test_en ) , .clk ( clk ) , 
    .ff_D ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_frac_logic_out[1] ) , 
    .ff_DI ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0_ff_Q ) , 
    .ff_Q ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1_ff_Q ) ,
    .ff_clk ( { SYNOPSYS_UNCONNECTED_2 } ) ,
    .p_abuf1 ( fabric_scout[0] ) , .p_abuf2 ( p_abuf2 ) ) ;
mux_tree_size2_21 mux_fabric_out_0 (
    .in ( { 
        logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0_ff_Q[0] , 
        logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_frac_logic_out[0]
         } ) ,
    .sram ( mux_tree_size2_0_sram ) , 
    .sram_inv ( mux_tree_size2_0_sram_inv ) , .out ( fabric_out[0] ) , 
    .p3 ( p3 ) ) ;
mux_tree_size2_22 mux_fabric_out_1 (
    .in ( { 
        logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1_ff_Q[0] , 
        logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_frac_logic_out[1]
         } ) ,
    .sram ( mux_tree_size2_1_sram ) , 
    .sram_inv ( mux_tree_size2_1_sram_inv ) , .out ( fabric_out[1] ) , 
    .p3 ( p3 ) ) ;
mux_tree_size2_23 mux_ff_0_D_0 (
    .in ( { 
        logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_frac_logic_out[0] , 
        fabric_regin[0] } ) ,
    .sram ( mux_tree_size2_2_sram ) , 
    .sram_inv ( mux_tree_size2_2_sram_inv ) , .out ( mux_tree_size2_2_out ) , 
    .p3 ( p3 ) ) ;
mux_tree_size2_mem_21 mem_fabric_out_0 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_size2_mem_0_ccff_tail ) , 
    .mem_out ( mux_tree_size2_0_sram ) , 
    .mem_outb ( mux_tree_size2_0_sram_inv ) ) ;
mux_tree_size2_mem_22 mem_fabric_out_1 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_size2_mem_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_size2_mem_1_ccff_tail ) , 
    .mem_out ( mux_tree_size2_1_sram ) , 
    .mem_outb ( mux_tree_size2_1_sram_inv ) ) ;
mux_tree_size2_mem_23 mem_ff_0_D_0 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_size2_mem_1_ccff_tail ) , .ccff_tail ( ccff_tail ) , 
    .mem_out ( mux_tree_size2_2_sram ) , 
    .mem_outb ( mux_tree_size2_2_sram_inv ) ) ;
direct_interc direct_interc_0_ (
    .in ( { SYNOPSYS_UNCONNECTED_3 } ) ,
    .out ( { p_abuf2 } ) ) ;
direct_interc direct_interc_1_ (
    .in ( { SYNOPSYS_UNCONNECTED_4 } ) ,
    .out ( { p_abuf2 } ) ) ;
direct_interc direct_interc_2_ (
    .in ( { SYNOPSYS_UNCONNECTED_5 } ) ,
    .out ( fabric_in[0] ) ) ;
direct_interc direct_interc_3_ (
    .in ( { SYNOPSYS_UNCONNECTED_6 } ) ,
    .out ( fabric_in[1] ) ) ;
direct_interc direct_interc_4_ (
    .in ( { SYNOPSYS_UNCONNECTED_7 } ) ,
    .out ( fabric_in[2] ) ) ;
direct_interc direct_interc_5_ (
    .in ( { SYNOPSYS_UNCONNECTED_8 } ) ,
    .out ( fabric_in[3] ) ) ;
direct_interc direct_interc_6_ (
    .in ( { SYNOPSYS_UNCONNECTED_9 } ) ,
    .out ( fabric_scin ) ) ;
direct_interc direct_interc_7_ (
    .in ( { SYNOPSYS_UNCONNECTED_10 } ) ,
    .out ( fabric_clk ) ) ;
direct_interc direct_interc_8_ (
    .in ( { SYNOPSYS_UNCONNECTED_11 } ) ,
    
    .out ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_frac_logic_out[1] ) ) ;
direct_interc direct_interc_9_ (
    .in ( { SYNOPSYS_UNCONNECTED_12 } ) ,
    
    .out ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0_ff_Q ) ) ;
direct_interc direct_interc_10_ (
    .in ( { SYNOPSYS_UNCONNECTED_13 } ) ,
    .out ( fabric_clk ) ) ;
sky130_fd_sc_hd__dlygate4sd1_1 FTB_1__263 ( .A ( fabric_scout[0] ) , 
    .X ( fabric_regout[0] ) ) ;
endmodule


module logical_tile_clb_mode_default__fle ( prog_clk , Test_en , clk , 
    fle_in , fle_regin , fle_scin , fle_clk , ccff_head , fle_out , 
    fle_regout , fle_scout , ccff_tail , p_abuf0 , p_abuf1 , p3 ) ;
input  [0:0] prog_clk ;
input  [0:0] Test_en ;
input  [0:0] clk ;
input  [0:3] fle_in ;
input  [0:0] fle_regin ;
input  [0:0] fle_scin ;
input  [0:0] fle_clk ;
input  [0:0] ccff_head ;
output [0:1] fle_out ;
output [0:0] fle_regout ;
output [0:0] fle_scout ;
output [0:0] ccff_tail ;
output p_abuf0 ;
output p_abuf1 ;
input  p3 ;

logical_tile_clb_mode_default__fle_mode_physical__fabric logical_tile_clb_mode_default__fle_mode_physical__fabric_0 ( 
    .prog_clk ( prog_clk ) , .Test_en ( Test_en ) , .clk ( clk ) , 
    .fabric_in ( fle_in ) , .fabric_regin ( fle_regin ) , 
    .fabric_scin ( fle_scin ) , .fabric_clk ( fle_clk ) , 
    .ccff_head ( ccff_head ) , .fabric_out ( fle_out ) , 
    .fabric_regout ( fle_regout ) , .fabric_scout ( fle_scout ) , 
    .ccff_tail ( ccff_tail ) , .p_abuf1 ( p_abuf0 ) , .p_abuf2 ( p_abuf1 ) , 
    .p3 ( p3 ) ) ;
direct_interc direct_interc_0_ (
    .in ( { SYNOPSYS_UNCONNECTED_1 } ) ,
    .out ( fle_out[0] ) ) ;
direct_interc direct_interc_1_ (
    .in ( { SYNOPSYS_UNCONNECTED_2 } ) ,
    .out ( fle_out[1] ) ) ;
direct_interc direct_interc_2_ (
    .in ( { SYNOPSYS_UNCONNECTED_3 } ) ,
    .out ( { p_abuf1 } ) ) ;
direct_interc direct_interc_3_ (
    .in ( { SYNOPSYS_UNCONNECTED_4 } ) ,
    .out ( { p_abuf0 } ) ) ;
direct_interc direct_interc_4_ (
    .in ( { SYNOPSYS_UNCONNECTED_5 } ) ,
    .out ( fle_in[0] ) ) ;
direct_interc direct_interc_5_ (
    .in ( { SYNOPSYS_UNCONNECTED_6 } ) ,
    .out ( fle_in[1] ) ) ;
direct_interc direct_interc_6_ (
    .in ( { SYNOPSYS_UNCONNECTED_7 } ) ,
    .out ( fle_in[2] ) ) ;
direct_interc direct_interc_7_ (
    .in ( { SYNOPSYS_UNCONNECTED_8 } ) ,
    .out ( fle_in[3] ) ) ;
direct_interc direct_interc_8_ (
    .in ( { SYNOPSYS_UNCONNECTED_9 } ) ,
    .out ( fle_regin ) ) ;
direct_interc direct_interc_9_ (
    .in ( { SYNOPSYS_UNCONNECTED_10 } ) ,
    .out ( fle_scin ) ) ;
direct_interc direct_interc_10_ (
    .in ( { SYNOPSYS_UNCONNECTED_11 } ) ,
    .out ( fle_clk ) ) ;
endmodule


module mux_tree_size2_mem_20 ( prog_clk , ccff_head , ccff_tail , mem_out , 
    mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_35__50 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_size2_mem_19 ( prog_clk , ccff_head , ccff_tail , mem_out , 
    mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_34__49 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_size2_mem_18 ( prog_clk , ccff_head , ccff_tail , mem_out , 
    mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_33__48 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_27 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_size2_20 ( in , sram , sram_inv , out , p3 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p3 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;

const1_27 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p3 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , .X ( out[0] ) ) ;
endmodule


module const1_26 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_size2_19 ( in , sram , sram_inv , out , p3 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p3 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;

const1_26 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p3 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , .X ( out[0] ) ) ;
endmodule


module const1_25 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_size2_18 ( in , sram , sram_inv , out , p3 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p3 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;

const1_25 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p3 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , .X ( out[0] ) ) ;
endmodule


module logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_13 ( 
    Test_en , clk , ff_D , ff_DI , ff_Q , ff_clk ) ;
input  [0:0] Test_en ;
input  [0:0] clk ;
input  [0:0] ff_D ;
input  [0:0] ff_DI ;
output [0:0] ff_Q ;
input  [0:0] ff_clk ;

sky130_fd_sc_hd__sdfxbp_1 sky130_fd_sc_hd__sdfxbp_1_0_ ( .D ( ff_D[0] ) , 
    .SCD ( ff_DI[0] ) , .SCE ( Test_en[0] ) , .CLK ( clk[0] ) , 
    .Q ( ff_Q[0] ) , .Q_N ( SYNOPSYS_UNCONNECTED_1 ) ) ;
endmodule


module logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_12 ( 
    Test_en , clk , ff_D , ff_DI , ff_Q , ff_clk ) ;
input  [0:0] Test_en ;
input  [0:0] clk ;
input  [0:0] ff_D ;
input  [0:0] ff_DI ;
output [0:0] ff_Q ;
input  [0:0] ff_clk ;

sky130_fd_sc_hd__sdfxbp_1 sky130_fd_sc_hd__sdfxbp_1_0_ ( .D ( ff_D[0] ) , 
    .SCD ( ff_DI[0] ) , .SCE ( Test_en[0] ) , .CLK ( clk[0] ) , 
    .Q ( ff_Q[0] ) , .Q_N ( SYNOPSYS_UNCONNECTED_1 ) ) ;
endmodule


module mux_tree_size2_mem_30 ( prog_clk , ccff_head , ccff_tail , mem_out , 
    mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_32__47 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_24 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_size2_30 ( in , sram , sram_inv , out , p2 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p2 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;

const1_24 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p2 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , .X ( out[0] ) ) ;
endmodule


module frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem_6 ( prog_clk , ccff_head , 
    ccff_tail , mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:16] mem_out ;
output [0:16] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_4_ ( .D ( mem_out[3] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[4] ) , .Q_N ( mem_outb[4] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_5_ ( .D ( mem_out[4] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[5] ) , .Q_N ( mem_outb[5] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_6_ ( .D ( mem_out[5] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[6] ) , .Q_N ( mem_outb[6] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_7_ ( .D ( mem_out[6] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[7] ) , .Q_N ( mem_outb[7] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_8_ ( .D ( mem_out[7] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[8] ) , .Q_N ( mem_outb[8] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_9_ ( .D ( mem_out[8] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[9] ) , .Q_N ( mem_outb[9] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_10_ ( .D ( mem_out[9] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[10] ) , .Q_N ( mem_outb[10] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_11_ ( .D ( mem_out[10] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[11] ) , .Q_N ( mem_outb[11] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_12_ ( .D ( mem_out[11] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[12] ) , .Q_N ( mem_outb[12] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_13_ ( .D ( mem_out[12] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[13] ) , .Q_N ( mem_outb[13] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_14_ ( .D ( mem_out[13] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[14] ) , .Q_N ( mem_outb[14] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_15_ ( .D ( mem_out[14] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[15] ) , .Q_N ( mem_outb[15] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_16_ ( .D ( mem_out[15] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[16] ) , .Q_N ( \_gOb6_mem_outb[16] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_31__46 ( .A ( mem_out[16] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module frac_lut4_mux_6 ( in , sram , sram_inv , lut3_out , lut4_out ) ;
input  [0:15] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:1] lut3_out ;
output [0:0] lut4_out ;

wire [0:0] sky130_fd_sc_hd__buf_2_3_X ;
wire [0:0] sky130_fd_sc_hd__buf_2_4_X ;
wire [0:0] sky130_fd_sc_hd__buf_2_5_X ;
wire [0:0] sky130_fd_sc_hd__buf_2_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_10_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_11_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_12_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_13_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_14_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_12_X[0] ) , .X ( lut3_out[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_1_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_13_X[0] ) , .X ( lut3_out[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_2_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_14_X[0] ) , .X ( lut4_out[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_3_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .X ( sky130_fd_sc_hd__buf_2_3_X[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_4_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , 
    .X ( sky130_fd_sc_hd__buf_2_4_X[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_5_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_10_X[0] ) , 
    .X ( sky130_fd_sc_hd__buf_2_5_X[0] ) ) ;
sky130_fd_sc_hd__buf_2 sky130_fd_sc_hd__buf_2_6_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_11_X[0] ) , 
    .X ( sky130_fd_sc_hd__buf_2_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_3_ ( .A0 ( in[7] ) , .A1 ( in[6] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_4_ ( .A0 ( in[9] ) , .A1 ( in[8] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_5_ ( .A0 ( in[11] ) , .A1 ( in[10] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_6_ ( .A0 ( in[13] ) , .A1 ( in[12] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_7_ ( .A0 ( in[15] ) , .A1 ( in[14] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_10_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_11_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( .A0 ( sky130_fd_sc_hd__buf_2_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__buf_2_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_12_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( .A0 ( sky130_fd_sc_hd__buf_2_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__buf_2_5_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_13_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_13_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_12_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_14_X[0] ) ) ;
endmodule


module frac_lut4_6 ( in , sram , sram_inv , mode , mode_inv , lut3_out , 
    lut4_out ) ;
input  [0:3] in ;
input  [0:15] sram ;
input  [0:15] sram_inv ;
input  [0:0] mode ;
input  [0:0] mode_inv ;
output [0:1] lut3_out ;
output [0:0] lut4_out ;

wire [0:0] sky130_fd_sc_hd__buf_2_0_X ;
wire [0:0] sky130_fd_sc_hd__buf_2_1_X ;
wire [0:0] sky130_fd_sc_hd__buf_2_2_X ;
wire [0:0] sky130_fd_sc_hd__buf_2_3_X ;
wire [0:0] sky130_fd_sc_hd__inv_1_0_Y ;
wire [0:0] sky130_fd_sc_hd__inv_1_1_Y ;
wire [0:0] sky130_fd_sc_hd__inv_1_2_Y ;
wire [0:0] sky130_fd_sc_hd__inv_1_3_Y ;
wire [0:0] sky130_fd_sc_hd__or2_1_0_X ;

sky130_fd_sc_hd__or2_0 sky130_fd_sc_hd__or2_1_0_ ( .A ( mode[0] ) , 
    .B ( in[3] ) , .X ( sky130_fd_sc_hd__or2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__inv_1 sky130_fd_sc_hd__inv_1_0_ ( .A ( in[0] ) , 
    .Y ( sky130_fd_sc_hd__inv_1_0_Y[0] ) ) ;
sky130_fd_sc_hd__inv_1 sky130_fd_sc_hd__inv_1_1_ ( .A ( in[1] ) , 
    .Y ( sky130_fd_sc_hd__inv_1_1_Y[0] ) ) ;
sky130_fd_sc_hd__inv_1 sky130_fd_sc_hd__inv_1_2_ ( .A ( in[2] ) , 
    .Y ( sky130_fd_sc_hd__inv_1_2_Y[0] ) ) ;
sky130_fd_sc_hd__inv_1 sky130_fd_sc_hd__inv_1_3_ ( 
    .A ( sky130_fd_sc_hd__or2_1_0_X[0] ) , 
    .Y ( sky130_fd_sc_hd__inv_1_3_Y[0] ) ) ;
sky130_fd_sc_hd__buf_2 sky130_fd_sc_hd__buf_2_0_ ( .A ( in[0] ) , 
    .X ( sky130_fd_sc_hd__buf_2_0_X[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_1_ ( .A ( in[1] ) , 
    .X ( sky130_fd_sc_hd__buf_2_1_X[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_2_ ( .A ( in[2] ) , 
    .X ( sky130_fd_sc_hd__buf_2_2_X[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_3_ ( 
    .A ( sky130_fd_sc_hd__or2_1_0_X[0] ) , 
    .X ( sky130_fd_sc_hd__buf_2_3_X[0] ) ) ;
frac_lut4_mux_6 frac_lut4_mux_0_ ( .in ( sram ) ,
    .sram ( { sky130_fd_sc_hd__buf_2_0_X[0] , sky130_fd_sc_hd__buf_2_1_X[0] , 
        sky130_fd_sc_hd__buf_2_2_X[0] , sky130_fd_sc_hd__buf_2_3_X[0] } ) ,
    .sram_inv ( { sky130_fd_sc_hd__inv_1_0_Y[0] , 
        sky130_fd_sc_hd__inv_1_1_Y[0] , sky130_fd_sc_hd__inv_1_2_Y[0] , 
        sky130_fd_sc_hd__inv_1_3_Y[0] } ) ,
    .lut3_out ( lut3_out ) , .lut4_out ( lut4_out ) ) ;
endmodule


module logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_6 ( 
    prog_clk , frac_lut4_in , ccff_head , frac_lut4_lut3_out , 
    frac_lut4_lut4_out , ccff_tail ) ;
input  [0:0] prog_clk ;
input  [0:3] frac_lut4_in ;
input  [0:0] ccff_head ;
output [0:1] frac_lut4_lut3_out ;
output [0:0] frac_lut4_lut4_out ;
output [0:0] ccff_tail ;

wire [0:0] frac_lut4_0_mode ;
wire [0:15] frac_lut4_0_sram ;
wire [0:15] frac_lut4_0_sram_inv ;

frac_lut4_6 frac_lut4_0_ ( .in ( frac_lut4_in ) , .sram ( frac_lut4_0_sram ) , 
    .sram_inv ( frac_lut4_0_sram_inv ) , .mode ( frac_lut4_0_mode ) ,
    .mode_inv ( { SYNOPSYS_UNCONNECTED_1 } ) ,
    .lut3_out ( frac_lut4_lut3_out ) , .lut4_out ( frac_lut4_lut4_out ) ) ;
frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem_6 frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem ( 
    .prog_clk ( prog_clk ) , .ccff_head ( ccff_head ) , 
    .ccff_tail ( ccff_tail ) ,
    .mem_out ( { frac_lut4_0_sram[0] , frac_lut4_0_sram[1] , 
        frac_lut4_0_sram[2] , frac_lut4_0_sram[3] , frac_lut4_0_sram[4] , 
        frac_lut4_0_sram[5] , frac_lut4_0_sram[6] , frac_lut4_0_sram[7] , 
        frac_lut4_0_sram[8] , frac_lut4_0_sram[9] , frac_lut4_0_sram[10] , 
        frac_lut4_0_sram[11] , frac_lut4_0_sram[12] , frac_lut4_0_sram[13] , 
        frac_lut4_0_sram[14] , frac_lut4_0_sram[15] , frac_lut4_0_mode[0] } ) ,
    .mem_outb ( { frac_lut4_0_sram_inv[0] , frac_lut4_0_sram_inv[1] , 
        frac_lut4_0_sram_inv[2] , frac_lut4_0_sram_inv[3] , 
        frac_lut4_0_sram_inv[4] , frac_lut4_0_sram_inv[5] , 
        frac_lut4_0_sram_inv[6] , frac_lut4_0_sram_inv[7] , 
        frac_lut4_0_sram_inv[8] , frac_lut4_0_sram_inv[9] , 
        frac_lut4_0_sram_inv[10] , frac_lut4_0_sram_inv[11] , 
        frac_lut4_0_sram_inv[12] , frac_lut4_0_sram_inv[13] , 
        frac_lut4_0_sram_inv[14] , frac_lut4_0_sram_inv[15] , 
        SYNOPSYS_UNCONNECTED_2 } ) ) ;
endmodule


module logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_6 ( 
    prog_clk , frac_logic_in , ccff_head , frac_logic_out , ccff_tail , p2 ) ;
input  [0:0] prog_clk ;
input  [0:3] frac_logic_in ;
input  [0:0] ccff_head ;
output [0:1] frac_logic_out ;
output [0:0] ccff_tail ;
input  p2 ;

wire [0:0] logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_ccff_tail ;
wire [0:0] logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_frac_lut4_lut3_out ;
wire [0:0] logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_frac_lut4_lut4_out ;
wire [0:1] mux_tree_size2_0_sram ;
wire [0:1] mux_tree_size2_0_sram_inv ;

logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_6 logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0 ( 
    .prog_clk ( prog_clk ) , .frac_lut4_in ( frac_logic_in ) , 
    .ccff_head ( ccff_head ) ,
    .frac_lut4_lut3_out ( { 
        logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_frac_lut4_lut3_out[0] , 
        frac_logic_out[1] } ) ,
    
    .frac_lut4_lut4_out ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_frac_lut4_lut4_out ) , 
    .ccff_tail ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_ccff_tail ) ) ;
mux_tree_size2_30 mux_frac_logic_out_0 (
    .in ( { 
        logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_frac_lut4_lut4_out[0] , 
        logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_frac_lut4_lut3_out[0]
         } ) ,
    .sram ( mux_tree_size2_0_sram ) , 
    .sram_inv ( mux_tree_size2_0_sram_inv ) , .out ( frac_logic_out[0] ) , 
    .p2 ( p2 ) ) ;
mux_tree_size2_mem_30 mem_frac_logic_out_0 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_ccff_tail ) , 
    .ccff_tail ( ccff_tail ) , .mem_out ( mux_tree_size2_0_sram ) , 
    .mem_outb ( mux_tree_size2_0_sram_inv ) ) ;
direct_interc direct_interc_0_ (
    .in ( { SYNOPSYS_UNCONNECTED_1 } ) ,
    .out ( frac_logic_out[1] ) ) ;
direct_interc direct_interc_1_ (
    .in ( { SYNOPSYS_UNCONNECTED_2 } ) ,
    .out ( frac_logic_in[0] ) ) ;
direct_interc direct_interc_2_ (
    .in ( { SYNOPSYS_UNCONNECTED_3 } ) ,
    .out ( frac_logic_in[1] ) ) ;
direct_interc direct_interc_3_ (
    .in ( { SYNOPSYS_UNCONNECTED_4 } ) ,
    .out ( frac_logic_in[2] ) ) ;
direct_interc direct_interc_4_ (
    .in ( { SYNOPSYS_UNCONNECTED_5 } ) ,
    .out ( frac_logic_in[3] ) ) ;
endmodule


module logical_tile_clb_mode_default__fle_mode_physical__fabric_6 ( prog_clk , 
    Test_en , clk , fabric_in , fabric_regin , fabric_scin , fabric_clk , 
    ccff_head , fabric_out , fabric_regout , fabric_scout , ccff_tail , p2 , 
    p3 ) ;
input  [0:0] prog_clk ;
input  [0:0] Test_en ;
input  [0:0] clk ;
input  [0:3] fabric_in ;
input  [0:0] fabric_regin ;
input  [0:0] fabric_scin ;
input  [0:0] fabric_clk ;
input  [0:0] ccff_head ;
output [0:1] fabric_out ;
output [0:0] fabric_regout ;
output [0:0] fabric_scout ;
output [0:0] ccff_tail ;
input  p2 ;
input  p3 ;

wire [0:0] logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0_ff_Q ;
wire [0:0] logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_ccff_tail ;
wire [0:1] logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_frac_logic_out ;
wire [0:1] mux_tree_size2_0_sram ;
wire [0:1] mux_tree_size2_0_sram_inv ;
wire [0:1] mux_tree_size2_1_sram ;
wire [0:1] mux_tree_size2_1_sram_inv ;
wire [0:0] mux_tree_size2_2_out ;
wire [0:1] mux_tree_size2_2_sram ;
wire [0:1] mux_tree_size2_2_sram_inv ;
wire [0:0] mux_tree_size2_mem_0_ccff_tail ;
wire [0:0] mux_tree_size2_mem_1_ccff_tail ;

assign fabric_regout[0] = fabric_scout[0] ;

logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_6 logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0 ( 
    .prog_clk ( prog_clk ) , .frac_logic_in ( fabric_in ) , 
    .ccff_head ( ccff_head ) , 
    .frac_logic_out ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_frac_logic_out ) , 
    .ccff_tail ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_ccff_tail ) , 
    .p2 ( p2 ) ) ;
logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_12 logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0 ( 
    .Test_en ( Test_en ) , .clk ( clk ) , .ff_D ( mux_tree_size2_2_out ) , 
    .ff_DI ( fabric_scin ) , 
    .ff_Q ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0_ff_Q ) ,
    .ff_clk ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_13 logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1 ( 
    .Test_en ( Test_en ) , .clk ( clk ) , 
    .ff_D ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_frac_logic_out[1] ) , 
    .ff_DI ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0_ff_Q ) , 
    .ff_Q ( fabric_scout ) ,
    .ff_clk ( { SYNOPSYS_UNCONNECTED_2 } ) ) ;
mux_tree_size2_18 mux_fabric_out_0 (
    .in ( { 
        logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0_ff_Q[0] , 
        logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_frac_logic_out[0]
         } ) ,
    .sram ( mux_tree_size2_0_sram ) , 
    .sram_inv ( mux_tree_size2_0_sram_inv ) , .out ( fabric_out[0] ) , 
    .p3 ( p3 ) ) ;
mux_tree_size2_19 mux_fabric_out_1 (
    .in ( { fabric_scout[0] , 
        logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_frac_logic_out[1]
         } ) ,
    .sram ( mux_tree_size2_1_sram ) , 
    .sram_inv ( mux_tree_size2_1_sram_inv ) , .out ( fabric_out[1] ) , 
    .p3 ( p3 ) ) ;
mux_tree_size2_20 mux_ff_0_D_0 (
    .in ( { 
        logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_frac_logic_out[0] , 
        fabric_regin[0] } ) ,
    .sram ( mux_tree_size2_2_sram ) , 
    .sram_inv ( mux_tree_size2_2_sram_inv ) , .out ( mux_tree_size2_2_out ) , 
    .p3 ( p3 ) ) ;
mux_tree_size2_mem_18 mem_fabric_out_0 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_size2_mem_0_ccff_tail ) , 
    .mem_out ( mux_tree_size2_0_sram ) , 
    .mem_outb ( mux_tree_size2_0_sram_inv ) ) ;
mux_tree_size2_mem_19 mem_fabric_out_1 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_size2_mem_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_size2_mem_1_ccff_tail ) , 
    .mem_out ( mux_tree_size2_1_sram ) , 
    .mem_outb ( mux_tree_size2_1_sram_inv ) ) ;
mux_tree_size2_mem_20 mem_ff_0_D_0 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_size2_mem_1_ccff_tail ) , .ccff_tail ( ccff_tail ) , 
    .mem_out ( mux_tree_size2_2_sram ) , 
    .mem_outb ( mux_tree_size2_2_sram_inv ) ) ;
direct_interc direct_interc_0_ (
    .in ( { SYNOPSYS_UNCONNECTED_3 } ) ,
    .out ( fabric_scout ) ) ;
direct_interc direct_interc_1_ (
    .in ( { SYNOPSYS_UNCONNECTED_4 } ) ,
    .out ( fabric_scout ) ) ;
direct_interc direct_interc_2_ (
    .in ( { SYNOPSYS_UNCONNECTED_5 } ) ,
    .out ( fabric_in[0] ) ) ;
direct_interc direct_interc_3_ (
    .in ( { SYNOPSYS_UNCONNECTED_6 } ) ,
    .out ( fabric_in[1] ) ) ;
direct_interc direct_interc_4_ (
    .in ( { SYNOPSYS_UNCONNECTED_7 } ) ,
    .out ( fabric_in[2] ) ) ;
direct_interc direct_interc_5_ (
    .in ( { SYNOPSYS_UNCONNECTED_8 } ) ,
    .out ( fabric_in[3] ) ) ;
direct_interc direct_interc_6_ (
    .in ( { SYNOPSYS_UNCONNECTED_9 } ) ,
    .out ( fabric_scin ) ) ;
direct_interc direct_interc_7_ (
    .in ( { SYNOPSYS_UNCONNECTED_10 } ) ,
    .out ( fabric_clk ) ) ;
direct_interc direct_interc_8_ (
    .in ( { SYNOPSYS_UNCONNECTED_11 } ) ,
    
    .out ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_frac_logic_out[1] ) ) ;
direct_interc direct_interc_9_ (
    .in ( { SYNOPSYS_UNCONNECTED_12 } ) ,
    
    .out ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0_ff_Q ) ) ;
direct_interc direct_interc_10_ (
    .in ( { SYNOPSYS_UNCONNECTED_13 } ) ,
    .out ( fabric_clk ) ) ;
endmodule


module logical_tile_clb_mode_default__fle_6 ( prog_clk , Test_en , clk , 
    fle_in , fle_regin , fle_scin , fle_clk , ccff_head , fle_out , 
    fle_regout , fle_scout , ccff_tail , p2 , p3 ) ;
input  [0:0] prog_clk ;
input  [0:0] Test_en ;
input  [0:0] clk ;
input  [0:3] fle_in ;
input  [0:0] fle_regin ;
input  [0:0] fle_scin ;
input  [0:0] fle_clk ;
input  [0:0] ccff_head ;
output [0:1] fle_out ;
output [0:0] fle_regout ;
output [0:0] fle_scout ;
output [0:0] ccff_tail ;
input  p2 ;
input  p3 ;

logical_tile_clb_mode_default__fle_mode_physical__fabric_6 logical_tile_clb_mode_default__fle_mode_physical__fabric_0 ( 
    .prog_clk ( prog_clk ) , .Test_en ( Test_en ) , .clk ( clk ) , 
    .fabric_in ( fle_in ) , .fabric_regin ( fle_regin ) , 
    .fabric_scin ( fle_scin ) , .fabric_clk ( fle_clk ) , 
    .ccff_head ( ccff_head ) , .fabric_out ( fle_out ) , 
    .fabric_regout ( fle_regout ) , .fabric_scout ( fle_scout ) , 
    .ccff_tail ( ccff_tail ) , .p2 ( p2 ) , .p3 ( p3 ) ) ;
direct_interc direct_interc_0_ (
    .in ( { SYNOPSYS_UNCONNECTED_1 } ) ,
    .out ( fle_out[0] ) ) ;
direct_interc direct_interc_1_ (
    .in ( { SYNOPSYS_UNCONNECTED_2 } ) ,
    .out ( fle_out[1] ) ) ;
direct_interc direct_interc_2_ (
    .in ( { SYNOPSYS_UNCONNECTED_3 } ) ,
    .out ( fle_regout ) ) ;
direct_interc direct_interc_3_ (
    .in ( { SYNOPSYS_UNCONNECTED_4 } ) ,
    .out ( fle_scout ) ) ;
direct_interc direct_interc_4_ (
    .in ( { SYNOPSYS_UNCONNECTED_5 } ) ,
    .out ( fle_in[0] ) ) ;
direct_interc direct_interc_5_ (
    .in ( { SYNOPSYS_UNCONNECTED_6 } ) ,
    .out ( fle_in[1] ) ) ;
direct_interc direct_interc_6_ (
    .in ( { SYNOPSYS_UNCONNECTED_7 } ) ,
    .out ( fle_in[2] ) ) ;
direct_interc direct_interc_7_ (
    .in ( { SYNOPSYS_UNCONNECTED_8 } ) ,
    .out ( fle_in[3] ) ) ;
direct_interc direct_interc_8_ (
    .in ( { SYNOPSYS_UNCONNECTED_9 } ) ,
    .out ( fle_regin ) ) ;
direct_interc direct_interc_9_ (
    .in ( { SYNOPSYS_UNCONNECTED_10 } ) ,
    .out ( fle_scin ) ) ;
direct_interc direct_interc_10_ (
    .in ( { SYNOPSYS_UNCONNECTED_11 } ) ,
    .out ( fle_clk ) ) ;
endmodule


module mux_tree_size2_mem_17 ( prog_clk , ccff_head , ccff_tail , mem_out , 
    mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_30__45 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_size2_mem_16 ( prog_clk , ccff_head , ccff_tail , mem_out , 
    mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_29__44 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_size2_mem_15 ( prog_clk , ccff_head , ccff_tail , mem_out , 
    mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_28__43 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_23 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_size2_17 ( in , sram , sram_inv , out , p2 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p2 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;

const1_23 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p2 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , .X ( out[0] ) ) ;
endmodule


module const1_22 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_size2_16 ( in , sram , sram_inv , out , p2 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p2 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;

const1_22 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p2 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , .X ( out[0] ) ) ;
endmodule


module const1_21 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_size2_15 ( in , sram , sram_inv , out , p2 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p2 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;

const1_21 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p2 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , .X ( out[0] ) ) ;
endmodule


module logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_11 ( 
    Test_en , clk , ff_D , ff_DI , ff_Q , ff_clk ) ;
input  [0:0] Test_en ;
input  [0:0] clk ;
input  [0:0] ff_D ;
input  [0:0] ff_DI ;
output [0:0] ff_Q ;
input  [0:0] ff_clk ;

sky130_fd_sc_hd__sdfxbp_1 sky130_fd_sc_hd__sdfxbp_1_0_ ( .D ( ff_D[0] ) , 
    .SCD ( ff_DI[0] ) , .SCE ( Test_en[0] ) , .CLK ( clk[0] ) , 
    .Q ( ff_Q[0] ) , .Q_N ( SYNOPSYS_UNCONNECTED_1 ) ) ;
endmodule


module logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_10 ( 
    Test_en , clk , ff_D , ff_DI , ff_Q , ff_clk ) ;
input  [0:0] Test_en ;
input  [0:0] clk ;
input  [0:0] ff_D ;
input  [0:0] ff_DI ;
output [0:0] ff_Q ;
input  [0:0] ff_clk ;

sky130_fd_sc_hd__sdfxbp_1 sky130_fd_sc_hd__sdfxbp_1_0_ ( .D ( ff_D[0] ) , 
    .SCD ( ff_DI[0] ) , .SCE ( Test_en[0] ) , .CLK ( clk[0] ) , 
    .Q ( ff_Q[0] ) , .Q_N ( SYNOPSYS_UNCONNECTED_1 ) ) ;
endmodule


module mux_tree_size2_mem_29 ( prog_clk , ccff_head , ccff_tail , mem_out , 
    mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_27__42 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_20 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_size2_29 ( in , sram , sram_inv , out , p2 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p2 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;

const1_20 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p2 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , .X ( out[0] ) ) ;
endmodule


module frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem_5 ( prog_clk , ccff_head , 
    ccff_tail , mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:16] mem_out ;
output [0:16] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_4_ ( .D ( mem_out[3] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[4] ) , .Q_N ( mem_outb[4] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_5_ ( .D ( mem_out[4] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[5] ) , .Q_N ( mem_outb[5] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_6_ ( .D ( mem_out[5] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[6] ) , .Q_N ( mem_outb[6] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_7_ ( .D ( mem_out[6] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[7] ) , .Q_N ( mem_outb[7] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_8_ ( .D ( mem_out[7] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[8] ) , .Q_N ( mem_outb[8] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_9_ ( .D ( mem_out[8] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[9] ) , .Q_N ( mem_outb[9] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_10_ ( .D ( mem_out[9] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[10] ) , .Q_N ( mem_outb[10] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_11_ ( .D ( mem_out[10] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[11] ) , .Q_N ( mem_outb[11] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_12_ ( .D ( mem_out[11] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[12] ) , .Q_N ( mem_outb[12] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_13_ ( .D ( mem_out[12] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[13] ) , .Q_N ( mem_outb[13] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_14_ ( .D ( mem_out[13] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[14] ) , .Q_N ( mem_outb[14] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_15_ ( .D ( mem_out[14] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[15] ) , .Q_N ( mem_outb[15] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_16_ ( .D ( mem_out[15] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[16] ) , .Q_N ( \_gOb5_mem_outb[16] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_26__41 ( .A ( mem_out[16] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module frac_lut4_mux_5 ( in , sram , sram_inv , lut3_out , lut4_out ) ;
input  [0:15] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:1] lut3_out ;
output [0:0] lut4_out ;

wire [0:0] sky130_fd_sc_hd__buf_2_3_X ;
wire [0:0] sky130_fd_sc_hd__buf_2_4_X ;
wire [0:0] sky130_fd_sc_hd__buf_2_5_X ;
wire [0:0] sky130_fd_sc_hd__buf_2_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_10_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_11_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_12_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_13_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_14_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_12_X[0] ) , .X ( lut3_out[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_1_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_13_X[0] ) , .X ( lut3_out[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_2_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_14_X[0] ) , .X ( lut4_out[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_3_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .X ( sky130_fd_sc_hd__buf_2_3_X[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_4_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , 
    .X ( sky130_fd_sc_hd__buf_2_4_X[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_5_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_10_X[0] ) , 
    .X ( sky130_fd_sc_hd__buf_2_5_X[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_6_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_11_X[0] ) , 
    .X ( sky130_fd_sc_hd__buf_2_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_3_ ( .A0 ( in[7] ) , .A1 ( in[6] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_4_ ( .A0 ( in[9] ) , .A1 ( in[8] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_5_ ( .A0 ( in[11] ) , .A1 ( in[10] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_6_ ( .A0 ( in[13] ) , .A1 ( in[12] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_7_ ( .A0 ( in[15] ) , .A1 ( in[14] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_10_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_11_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( .A0 ( sky130_fd_sc_hd__buf_2_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__buf_2_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_12_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( .A0 ( sky130_fd_sc_hd__buf_2_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__buf_2_5_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_13_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_13_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_12_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_14_X[0] ) ) ;
endmodule


module frac_lut4_5 ( in , sram , sram_inv , mode , mode_inv , lut3_out , 
    lut4_out ) ;
input  [0:3] in ;
input  [0:15] sram ;
input  [0:15] sram_inv ;
input  [0:0] mode ;
input  [0:0] mode_inv ;
output [0:1] lut3_out ;
output [0:0] lut4_out ;

wire [0:0] sky130_fd_sc_hd__buf_2_0_X ;
wire [0:0] sky130_fd_sc_hd__buf_2_1_X ;
wire [0:0] sky130_fd_sc_hd__buf_2_2_X ;
wire [0:0] sky130_fd_sc_hd__buf_2_3_X ;
wire [0:0] sky130_fd_sc_hd__inv_1_0_Y ;
wire [0:0] sky130_fd_sc_hd__inv_1_1_Y ;
wire [0:0] sky130_fd_sc_hd__inv_1_2_Y ;
wire [0:0] sky130_fd_sc_hd__inv_1_3_Y ;
wire [0:0] sky130_fd_sc_hd__or2_1_0_X ;

sky130_fd_sc_hd__or2_0 sky130_fd_sc_hd__or2_1_0_ ( .A ( mode[0] ) , 
    .B ( in[3] ) , .X ( sky130_fd_sc_hd__or2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__inv_1 sky130_fd_sc_hd__inv_1_0_ ( .A ( in[0] ) , 
    .Y ( sky130_fd_sc_hd__inv_1_0_Y[0] ) ) ;
sky130_fd_sc_hd__inv_1 sky130_fd_sc_hd__inv_1_1_ ( .A ( in[1] ) , 
    .Y ( sky130_fd_sc_hd__inv_1_1_Y[0] ) ) ;
sky130_fd_sc_hd__inv_1 sky130_fd_sc_hd__inv_1_2_ ( .A ( in[2] ) , 
    .Y ( sky130_fd_sc_hd__inv_1_2_Y[0] ) ) ;
sky130_fd_sc_hd__inv_1 sky130_fd_sc_hd__inv_1_3_ ( 
    .A ( sky130_fd_sc_hd__or2_1_0_X[0] ) , 
    .Y ( sky130_fd_sc_hd__inv_1_3_Y[0] ) ) ;
sky130_fd_sc_hd__buf_2 sky130_fd_sc_hd__buf_2_0_ ( .A ( in[0] ) , 
    .X ( sky130_fd_sc_hd__buf_2_0_X[0] ) ) ;
sky130_fd_sc_hd__buf_2 sky130_fd_sc_hd__buf_2_1_ ( .A ( in[1] ) , 
    .X ( sky130_fd_sc_hd__buf_2_1_X[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_2_ ( .A ( in[2] ) , 
    .X ( sky130_fd_sc_hd__buf_2_2_X[0] ) ) ;
sky130_fd_sc_hd__buf_2 sky130_fd_sc_hd__buf_2_3_ ( 
    .A ( sky130_fd_sc_hd__or2_1_0_X[0] ) , 
    .X ( sky130_fd_sc_hd__buf_2_3_X[0] ) ) ;
frac_lut4_mux_5 frac_lut4_mux_0_ ( .in ( sram ) ,
    .sram ( { sky130_fd_sc_hd__buf_2_0_X[0] , sky130_fd_sc_hd__buf_2_1_X[0] , 
        sky130_fd_sc_hd__buf_2_2_X[0] , sky130_fd_sc_hd__buf_2_3_X[0] } ) ,
    .sram_inv ( { sky130_fd_sc_hd__inv_1_0_Y[0] , 
        sky130_fd_sc_hd__inv_1_1_Y[0] , sky130_fd_sc_hd__inv_1_2_Y[0] , 
        sky130_fd_sc_hd__inv_1_3_Y[0] } ) ,
    .lut3_out ( lut3_out ) , .lut4_out ( lut4_out ) ) ;
endmodule


module logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_5 ( 
    prog_clk , frac_lut4_in , ccff_head , frac_lut4_lut3_out , 
    frac_lut4_lut4_out , ccff_tail ) ;
input  [0:0] prog_clk ;
input  [0:3] frac_lut4_in ;
input  [0:0] ccff_head ;
output [0:1] frac_lut4_lut3_out ;
output [0:0] frac_lut4_lut4_out ;
output [0:0] ccff_tail ;

wire [0:0] frac_lut4_0_mode ;
wire [0:15] frac_lut4_0_sram ;
wire [0:15] frac_lut4_0_sram_inv ;

frac_lut4_5 frac_lut4_0_ ( .in ( frac_lut4_in ) , .sram ( frac_lut4_0_sram ) , 
    .sram_inv ( frac_lut4_0_sram_inv ) , .mode ( frac_lut4_0_mode ) ,
    .mode_inv ( { SYNOPSYS_UNCONNECTED_1 } ) ,
    .lut3_out ( frac_lut4_lut3_out ) , .lut4_out ( frac_lut4_lut4_out ) ) ;
frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem_5 frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem ( 
    .prog_clk ( prog_clk ) , .ccff_head ( ccff_head ) , 
    .ccff_tail ( ccff_tail ) ,
    .mem_out ( { frac_lut4_0_sram[0] , frac_lut4_0_sram[1] , 
        frac_lut4_0_sram[2] , frac_lut4_0_sram[3] , frac_lut4_0_sram[4] , 
        frac_lut4_0_sram[5] , frac_lut4_0_sram[6] , frac_lut4_0_sram[7] , 
        frac_lut4_0_sram[8] , frac_lut4_0_sram[9] , frac_lut4_0_sram[10] , 
        frac_lut4_0_sram[11] , frac_lut4_0_sram[12] , frac_lut4_0_sram[13] , 
        frac_lut4_0_sram[14] , frac_lut4_0_sram[15] , frac_lut4_0_mode[0] } ) ,
    .mem_outb ( { frac_lut4_0_sram_inv[0] , frac_lut4_0_sram_inv[1] , 
        frac_lut4_0_sram_inv[2] , frac_lut4_0_sram_inv[3] , 
        frac_lut4_0_sram_inv[4] , frac_lut4_0_sram_inv[5] , 
        frac_lut4_0_sram_inv[6] , frac_lut4_0_sram_inv[7] , 
        frac_lut4_0_sram_inv[8] , frac_lut4_0_sram_inv[9] , 
        frac_lut4_0_sram_inv[10] , frac_lut4_0_sram_inv[11] , 
        frac_lut4_0_sram_inv[12] , frac_lut4_0_sram_inv[13] , 
        frac_lut4_0_sram_inv[14] , frac_lut4_0_sram_inv[15] , 
        SYNOPSYS_UNCONNECTED_2 } ) ) ;
endmodule


module logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_5 ( 
    prog_clk , frac_logic_in , ccff_head , frac_logic_out , ccff_tail , p2 ) ;
input  [0:0] prog_clk ;
input  [0:3] frac_logic_in ;
input  [0:0] ccff_head ;
output [0:1] frac_logic_out ;
output [0:0] ccff_tail ;
input  p2 ;

wire [0:0] logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_ccff_tail ;
wire [0:0] logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_frac_lut4_lut3_out ;
wire [0:0] logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_frac_lut4_lut4_out ;
wire [0:1] mux_tree_size2_0_sram ;
wire [0:1] mux_tree_size2_0_sram_inv ;

logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_5 logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0 ( 
    .prog_clk ( prog_clk ) , .frac_lut4_in ( frac_logic_in ) , 
    .ccff_head ( ccff_head ) ,
    .frac_lut4_lut3_out ( { 
        logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_frac_lut4_lut3_out[0] , 
        frac_logic_out[1] } ) ,
    
    .frac_lut4_lut4_out ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_frac_lut4_lut4_out ) , 
    .ccff_tail ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_ccff_tail ) ) ;
mux_tree_size2_29 mux_frac_logic_out_0 (
    .in ( { 
        logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_frac_lut4_lut4_out[0] , 
        logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_frac_lut4_lut3_out[0]
         } ) ,
    .sram ( mux_tree_size2_0_sram ) , 
    .sram_inv ( mux_tree_size2_0_sram_inv ) , .out ( frac_logic_out[0] ) , 
    .p2 ( p2 ) ) ;
mux_tree_size2_mem_29 mem_frac_logic_out_0 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_ccff_tail ) , 
    .ccff_tail ( ccff_tail ) , .mem_out ( mux_tree_size2_0_sram ) , 
    .mem_outb ( mux_tree_size2_0_sram_inv ) ) ;
direct_interc direct_interc_0_ (
    .in ( { SYNOPSYS_UNCONNECTED_1 } ) ,
    .out ( frac_logic_out[1] ) ) ;
direct_interc direct_interc_1_ (
    .in ( { SYNOPSYS_UNCONNECTED_2 } ) ,
    .out ( frac_logic_in[0] ) ) ;
direct_interc direct_interc_2_ (
    .in ( { SYNOPSYS_UNCONNECTED_3 } ) ,
    .out ( frac_logic_in[1] ) ) ;
direct_interc direct_interc_3_ (
    .in ( { SYNOPSYS_UNCONNECTED_4 } ) ,
    .out ( frac_logic_in[2] ) ) ;
direct_interc direct_interc_4_ (
    .in ( { SYNOPSYS_UNCONNECTED_5 } ) ,
    .out ( frac_logic_in[3] ) ) ;
endmodule


module logical_tile_clb_mode_default__fle_mode_physical__fabric_5 ( prog_clk , 
    Test_en , clk , fabric_in , fabric_regin , fabric_scin , fabric_clk , 
    ccff_head , fabric_out , fabric_regout , fabric_scout , ccff_tail , p2 ) ;
input  [0:0] prog_clk ;
input  [0:0] Test_en ;
input  [0:0] clk ;
input  [0:3] fabric_in ;
input  [0:0] fabric_regin ;
input  [0:0] fabric_scin ;
input  [0:0] fabric_clk ;
input  [0:0] ccff_head ;
output [0:1] fabric_out ;
output [0:0] fabric_regout ;
output [0:0] fabric_scout ;
output [0:0] ccff_tail ;
input  p2 ;

wire [0:0] logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0_ff_Q ;
wire [0:0] logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_ccff_tail ;
wire [0:1] logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_frac_logic_out ;
wire [0:1] mux_tree_size2_0_sram ;
wire [0:1] mux_tree_size2_0_sram_inv ;
wire [0:1] mux_tree_size2_1_sram ;
wire [0:1] mux_tree_size2_1_sram_inv ;
wire [0:0] mux_tree_size2_2_out ;
wire [0:1] mux_tree_size2_2_sram ;
wire [0:1] mux_tree_size2_2_sram_inv ;
wire [0:0] mux_tree_size2_mem_0_ccff_tail ;
wire [0:0] mux_tree_size2_mem_1_ccff_tail ;

assign fabric_regout[0] = fabric_scout[0] ;

logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_5 logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0 ( 
    .prog_clk ( prog_clk ) , .frac_logic_in ( fabric_in ) , 
    .ccff_head ( ccff_head ) , 
    .frac_logic_out ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_frac_logic_out ) , 
    .ccff_tail ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_ccff_tail ) , 
    .p2 ( p2 ) ) ;
logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_10 logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0 ( 
    .Test_en ( Test_en ) , .clk ( clk ) , .ff_D ( mux_tree_size2_2_out ) , 
    .ff_DI ( fabric_scin ) , 
    .ff_Q ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0_ff_Q ) ,
    .ff_clk ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_11 logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1 ( 
    .Test_en ( Test_en ) , .clk ( clk ) , 
    .ff_D ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_frac_logic_out[1] ) , 
    .ff_DI ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0_ff_Q ) , 
    .ff_Q ( fabric_scout ) ,
    .ff_clk ( { SYNOPSYS_UNCONNECTED_2 } ) ) ;
mux_tree_size2_15 mux_fabric_out_0 (
    .in ( { 
        logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0_ff_Q[0] , 
        logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_frac_logic_out[0]
         } ) ,
    .sram ( mux_tree_size2_0_sram ) , 
    .sram_inv ( mux_tree_size2_0_sram_inv ) , .out ( fabric_out[0] ) , 
    .p2 ( p2 ) ) ;
mux_tree_size2_16 mux_fabric_out_1 (
    .in ( { fabric_scout[0] , 
        logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_frac_logic_out[1]
         } ) ,
    .sram ( mux_tree_size2_1_sram ) , 
    .sram_inv ( mux_tree_size2_1_sram_inv ) , .out ( fabric_out[1] ) , 
    .p2 ( p2 ) ) ;
mux_tree_size2_17 mux_ff_0_D_0 (
    .in ( { 
        logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_frac_logic_out[0] , 
        fabric_regin[0] } ) ,
    .sram ( mux_tree_size2_2_sram ) , 
    .sram_inv ( mux_tree_size2_2_sram_inv ) , .out ( mux_tree_size2_2_out ) , 
    .p2 ( p2 ) ) ;
mux_tree_size2_mem_15 mem_fabric_out_0 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_size2_mem_0_ccff_tail ) , 
    .mem_out ( mux_tree_size2_0_sram ) , 
    .mem_outb ( mux_tree_size2_0_sram_inv ) ) ;
mux_tree_size2_mem_16 mem_fabric_out_1 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_size2_mem_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_size2_mem_1_ccff_tail ) , 
    .mem_out ( mux_tree_size2_1_sram ) , 
    .mem_outb ( mux_tree_size2_1_sram_inv ) ) ;
mux_tree_size2_mem_17 mem_ff_0_D_0 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_size2_mem_1_ccff_tail ) , .ccff_tail ( ccff_tail ) , 
    .mem_out ( mux_tree_size2_2_sram ) , 
    .mem_outb ( mux_tree_size2_2_sram_inv ) ) ;
direct_interc direct_interc_0_ (
    .in ( { SYNOPSYS_UNCONNECTED_3 } ) ,
    .out ( fabric_scout ) ) ;
direct_interc direct_interc_1_ (
    .in ( { SYNOPSYS_UNCONNECTED_4 } ) ,
    .out ( fabric_scout ) ) ;
direct_interc direct_interc_2_ (
    .in ( { SYNOPSYS_UNCONNECTED_5 } ) ,
    .out ( fabric_in[0] ) ) ;
direct_interc direct_interc_3_ (
    .in ( { SYNOPSYS_UNCONNECTED_6 } ) ,
    .out ( fabric_in[1] ) ) ;
direct_interc direct_interc_4_ (
    .in ( { SYNOPSYS_UNCONNECTED_7 } ) ,
    .out ( fabric_in[2] ) ) ;
direct_interc direct_interc_5_ (
    .in ( { SYNOPSYS_UNCONNECTED_8 } ) ,
    .out ( fabric_in[3] ) ) ;
direct_interc direct_interc_6_ (
    .in ( { SYNOPSYS_UNCONNECTED_9 } ) ,
    .out ( fabric_scin ) ) ;
direct_interc direct_interc_7_ (
    .in ( { SYNOPSYS_UNCONNECTED_10 } ) ,
    .out ( fabric_clk ) ) ;
direct_interc direct_interc_8_ (
    .in ( { SYNOPSYS_UNCONNECTED_11 } ) ,
    
    .out ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_frac_logic_out[1] ) ) ;
direct_interc direct_interc_9_ (
    .in ( { SYNOPSYS_UNCONNECTED_12 } ) ,
    
    .out ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0_ff_Q ) ) ;
direct_interc direct_interc_10_ (
    .in ( { SYNOPSYS_UNCONNECTED_13 } ) ,
    .out ( fabric_clk ) ) ;
endmodule


module logical_tile_clb_mode_default__fle_5 ( prog_clk , Test_en , clk , 
    fle_in , fle_regin , fle_scin , fle_clk , ccff_head , fle_out , 
    fle_regout , fle_scout , ccff_tail , p2 ) ;
input  [0:0] prog_clk ;
input  [0:0] Test_en ;
input  [0:0] clk ;
input  [0:3] fle_in ;
input  [0:0] fle_regin ;
input  [0:0] fle_scin ;
input  [0:0] fle_clk ;
input  [0:0] ccff_head ;
output [0:1] fle_out ;
output [0:0] fle_regout ;
output [0:0] fle_scout ;
output [0:0] ccff_tail ;
input  p2 ;

logical_tile_clb_mode_default__fle_mode_physical__fabric_5 logical_tile_clb_mode_default__fle_mode_physical__fabric_0 ( 
    .prog_clk ( prog_clk ) , .Test_en ( Test_en ) , .clk ( clk ) , 
    .fabric_in ( fle_in ) , .fabric_regin ( fle_regin ) , 
    .fabric_scin ( fle_scin ) , .fabric_clk ( fle_clk ) , 
    .ccff_head ( ccff_head ) , .fabric_out ( fle_out ) , 
    .fabric_regout ( fle_regout ) , .fabric_scout ( fle_scout ) , 
    .ccff_tail ( ccff_tail ) , .p2 ( p2 ) ) ;
direct_interc direct_interc_0_ (
    .in ( { SYNOPSYS_UNCONNECTED_1 } ) ,
    .out ( fle_out[0] ) ) ;
direct_interc direct_interc_1_ (
    .in ( { SYNOPSYS_UNCONNECTED_2 } ) ,
    .out ( fle_out[1] ) ) ;
direct_interc direct_interc_2_ (
    .in ( { SYNOPSYS_UNCONNECTED_3 } ) ,
    .out ( fle_regout ) ) ;
direct_interc direct_interc_3_ (
    .in ( { SYNOPSYS_UNCONNECTED_4 } ) ,
    .out ( fle_scout ) ) ;
direct_interc direct_interc_4_ (
    .in ( { SYNOPSYS_UNCONNECTED_5 } ) ,
    .out ( fle_in[0] ) ) ;
direct_interc direct_interc_5_ (
    .in ( { SYNOPSYS_UNCONNECTED_6 } ) ,
    .out ( fle_in[1] ) ) ;
direct_interc direct_interc_6_ (
    .in ( { SYNOPSYS_UNCONNECTED_7 } ) ,
    .out ( fle_in[2] ) ) ;
direct_interc direct_interc_7_ (
    .in ( { SYNOPSYS_UNCONNECTED_8 } ) ,
    .out ( fle_in[3] ) ) ;
direct_interc direct_interc_8_ (
    .in ( { SYNOPSYS_UNCONNECTED_9 } ) ,
    .out ( fle_regin ) ) ;
direct_interc direct_interc_9_ (
    .in ( { SYNOPSYS_UNCONNECTED_10 } ) ,
    .out ( fle_scin ) ) ;
direct_interc direct_interc_10_ (
    .in ( { SYNOPSYS_UNCONNECTED_11 } ) ,
    .out ( fle_clk ) ) ;
endmodule


module mux_tree_size2_mem_14 ( prog_clk , ccff_head , ccff_tail , mem_out , 
    mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_25__40 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_size2_mem_13 ( prog_clk , ccff_head , ccff_tail , mem_out , 
    mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_24__39 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_size2_mem_12 ( prog_clk , ccff_head , ccff_tail , mem_out , 
    mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_23__38 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_19 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_size2_14 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;

const1_19 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , .X ( out[0] ) ) ;
endmodule


module const1_18 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_size2_13 ( in , sram , sram_inv , out , p2 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p2 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;

const1_18 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p2 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , .X ( out[0] ) ) ;
endmodule


module const1_17 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_size2_12 ( in , sram , sram_inv , out , p2 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p2 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;

const1_17 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p2 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , .X ( out[0] ) ) ;
endmodule


module logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_9 ( 
    Test_en , clk , ff_D , ff_DI , ff_Q , ff_clk ) ;
input  [0:0] Test_en ;
input  [0:0] clk ;
input  [0:0] ff_D ;
input  [0:0] ff_DI ;
output [0:0] ff_Q ;
input  [0:0] ff_clk ;

sky130_fd_sc_hd__sdfxbp_1 sky130_fd_sc_hd__sdfxbp_1_0_ ( .D ( ff_D[0] ) , 
    .SCD ( ff_DI[0] ) , .SCE ( Test_en[0] ) , .CLK ( clk[0] ) , 
    .Q ( ff_Q[0] ) , .Q_N ( SYNOPSYS_UNCONNECTED_1 ) ) ;
endmodule


module logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_8 ( 
    Test_en , clk , ff_D , ff_DI , ff_Q , ff_clk ) ;
input  [0:0] Test_en ;
input  [0:0] clk ;
input  [0:0] ff_D ;
input  [0:0] ff_DI ;
output [0:0] ff_Q ;
input  [0:0] ff_clk ;

sky130_fd_sc_hd__sdfxbp_1 sky130_fd_sc_hd__sdfxbp_1_0_ ( .D ( ff_D[0] ) , 
    .SCD ( ff_DI[0] ) , .SCE ( Test_en[0] ) , .CLK ( clk[0] ) , 
    .Q ( ff_Q[0] ) , .Q_N ( SYNOPSYS_UNCONNECTED_1 ) ) ;
endmodule


module mux_tree_size2_mem_28 ( prog_clk , ccff_head , ccff_tail , mem_out , 
    mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_22__37 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_16 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_size2_28 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;

const1_16 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , .X ( out[0] ) ) ;
endmodule


module frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem_4 ( prog_clk , ccff_head , 
    ccff_tail , mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:16] mem_out ;
output [0:16] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_4_ ( .D ( mem_out[3] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[4] ) , .Q_N ( mem_outb[4] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_5_ ( .D ( mem_out[4] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[5] ) , .Q_N ( mem_outb[5] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_6_ ( .D ( mem_out[5] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[6] ) , .Q_N ( mem_outb[6] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_7_ ( .D ( mem_out[6] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[7] ) , .Q_N ( mem_outb[7] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_8_ ( .D ( mem_out[7] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[8] ) , .Q_N ( mem_outb[8] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_9_ ( .D ( mem_out[8] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[9] ) , .Q_N ( mem_outb[9] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_10_ ( .D ( mem_out[9] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[10] ) , .Q_N ( mem_outb[10] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_11_ ( .D ( mem_out[10] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[11] ) , .Q_N ( mem_outb[11] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_12_ ( .D ( mem_out[11] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[12] ) , .Q_N ( mem_outb[12] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_13_ ( .D ( mem_out[12] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[13] ) , .Q_N ( mem_outb[13] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_14_ ( .D ( mem_out[13] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[14] ) , .Q_N ( mem_outb[14] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_15_ ( .D ( mem_out[14] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[15] ) , .Q_N ( mem_outb[15] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_16_ ( .D ( mem_out[15] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[16] ) , .Q_N ( \_gOb4_mem_outb[16] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_21__36 ( .A ( mem_out[16] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module frac_lut4_mux_4 ( in , sram , sram_inv , lut3_out , lut4_out ) ;
input  [0:15] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:1] lut3_out ;
output [0:0] lut4_out ;

wire [0:0] sky130_fd_sc_hd__buf_2_3_X ;
wire [0:0] sky130_fd_sc_hd__buf_2_4_X ;
wire [0:0] sky130_fd_sc_hd__buf_2_5_X ;
wire [0:0] sky130_fd_sc_hd__buf_2_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_10_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_11_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_12_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_13_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_14_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_12_X[0] ) , .X ( lut3_out[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_1_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_13_X[0] ) , .X ( lut3_out[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_2_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_14_X[0] ) , .X ( lut4_out[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_3_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .X ( sky130_fd_sc_hd__buf_2_3_X[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_4_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , 
    .X ( sky130_fd_sc_hd__buf_2_4_X[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_5_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_10_X[0] ) , 
    .X ( sky130_fd_sc_hd__buf_2_5_X[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_6_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_11_X[0] ) , 
    .X ( sky130_fd_sc_hd__buf_2_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_3_ ( .A0 ( in[7] ) , .A1 ( in[6] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_4_ ( .A0 ( in[9] ) , .A1 ( in[8] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_5_ ( .A0 ( in[11] ) , .A1 ( in[10] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_6_ ( .A0 ( in[13] ) , .A1 ( in[12] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_7_ ( .A0 ( in[15] ) , .A1 ( in[14] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_10_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_11_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( .A0 ( sky130_fd_sc_hd__buf_2_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__buf_2_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_12_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( .A0 ( sky130_fd_sc_hd__buf_2_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__buf_2_5_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_13_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_13_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_12_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_14_X[0] ) ) ;
endmodule


module frac_lut4_4 ( in , sram , sram_inv , mode , mode_inv , lut3_out , 
    lut4_out ) ;
input  [0:3] in ;
input  [0:15] sram ;
input  [0:15] sram_inv ;
input  [0:0] mode ;
input  [0:0] mode_inv ;
output [0:1] lut3_out ;
output [0:0] lut4_out ;

wire [0:0] sky130_fd_sc_hd__buf_2_0_X ;
wire [0:0] sky130_fd_sc_hd__buf_2_1_X ;
wire [0:0] sky130_fd_sc_hd__buf_2_2_X ;
wire [0:0] sky130_fd_sc_hd__buf_2_3_X ;
wire [0:0] sky130_fd_sc_hd__inv_1_0_Y ;
wire [0:0] sky130_fd_sc_hd__inv_1_1_Y ;
wire [0:0] sky130_fd_sc_hd__inv_1_2_Y ;
wire [0:0] sky130_fd_sc_hd__inv_1_3_Y ;
wire [0:0] sky130_fd_sc_hd__or2_1_0_X ;

sky130_fd_sc_hd__or2_0 sky130_fd_sc_hd__or2_1_0_ ( .A ( mode[0] ) , 
    .B ( in[3] ) , .X ( sky130_fd_sc_hd__or2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__inv_1 sky130_fd_sc_hd__inv_1_0_ ( .A ( in[0] ) , 
    .Y ( sky130_fd_sc_hd__inv_1_0_Y[0] ) ) ;
sky130_fd_sc_hd__inv_1 sky130_fd_sc_hd__inv_1_1_ ( .A ( in[1] ) , 
    .Y ( sky130_fd_sc_hd__inv_1_1_Y[0] ) ) ;
sky130_fd_sc_hd__inv_1 sky130_fd_sc_hd__inv_1_2_ ( .A ( in[2] ) , 
    .Y ( sky130_fd_sc_hd__inv_1_2_Y[0] ) ) ;
sky130_fd_sc_hd__inv_1 sky130_fd_sc_hd__inv_1_3_ ( 
    .A ( sky130_fd_sc_hd__or2_1_0_X[0] ) , 
    .Y ( sky130_fd_sc_hd__inv_1_3_Y[0] ) ) ;
sky130_fd_sc_hd__buf_2 sky130_fd_sc_hd__buf_2_0_ ( .A ( in[0] ) , 
    .X ( sky130_fd_sc_hd__buf_2_0_X[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_1_ ( .A ( in[1] ) , 
    .X ( sky130_fd_sc_hd__buf_2_1_X[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_2_ ( .A ( in[2] ) , 
    .X ( sky130_fd_sc_hd__buf_2_2_X[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_3_ ( 
    .A ( sky130_fd_sc_hd__or2_1_0_X[0] ) , 
    .X ( sky130_fd_sc_hd__buf_2_3_X[0] ) ) ;
frac_lut4_mux_4 frac_lut4_mux_0_ ( .in ( sram ) ,
    .sram ( { sky130_fd_sc_hd__buf_2_0_X[0] , sky130_fd_sc_hd__buf_2_1_X[0] , 
        sky130_fd_sc_hd__buf_2_2_X[0] , sky130_fd_sc_hd__buf_2_3_X[0] } ) ,
    .sram_inv ( { sky130_fd_sc_hd__inv_1_0_Y[0] , 
        sky130_fd_sc_hd__inv_1_1_Y[0] , sky130_fd_sc_hd__inv_1_2_Y[0] , 
        sky130_fd_sc_hd__inv_1_3_Y[0] } ) ,
    .lut3_out ( lut3_out ) , .lut4_out ( lut4_out ) ) ;
endmodule


module logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_4 ( 
    prog_clk , frac_lut4_in , ccff_head , frac_lut4_lut3_out , 
    frac_lut4_lut4_out , ccff_tail ) ;
input  [0:0] prog_clk ;
input  [0:3] frac_lut4_in ;
input  [0:0] ccff_head ;
output [0:1] frac_lut4_lut3_out ;
output [0:0] frac_lut4_lut4_out ;
output [0:0] ccff_tail ;

wire [0:0] frac_lut4_0_mode ;
wire [0:15] frac_lut4_0_sram ;
wire [0:15] frac_lut4_0_sram_inv ;

frac_lut4_4 frac_lut4_0_ ( .in ( frac_lut4_in ) , .sram ( frac_lut4_0_sram ) , 
    .sram_inv ( frac_lut4_0_sram_inv ) , .mode ( frac_lut4_0_mode ) ,
    .mode_inv ( { SYNOPSYS_UNCONNECTED_1 } ) ,
    .lut3_out ( frac_lut4_lut3_out ) , .lut4_out ( frac_lut4_lut4_out ) ) ;
frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem_4 frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem ( 
    .prog_clk ( prog_clk ) , .ccff_head ( ccff_head ) , 
    .ccff_tail ( ccff_tail ) ,
    .mem_out ( { frac_lut4_0_sram[0] , frac_lut4_0_sram[1] , 
        frac_lut4_0_sram[2] , frac_lut4_0_sram[3] , frac_lut4_0_sram[4] , 
        frac_lut4_0_sram[5] , frac_lut4_0_sram[6] , frac_lut4_0_sram[7] , 
        frac_lut4_0_sram[8] , frac_lut4_0_sram[9] , frac_lut4_0_sram[10] , 
        frac_lut4_0_sram[11] , frac_lut4_0_sram[12] , frac_lut4_0_sram[13] , 
        frac_lut4_0_sram[14] , frac_lut4_0_sram[15] , frac_lut4_0_mode[0] } ) ,
    .mem_outb ( { frac_lut4_0_sram_inv[0] , frac_lut4_0_sram_inv[1] , 
        frac_lut4_0_sram_inv[2] , frac_lut4_0_sram_inv[3] , 
        frac_lut4_0_sram_inv[4] , frac_lut4_0_sram_inv[5] , 
        frac_lut4_0_sram_inv[6] , frac_lut4_0_sram_inv[7] , 
        frac_lut4_0_sram_inv[8] , frac_lut4_0_sram_inv[9] , 
        frac_lut4_0_sram_inv[10] , frac_lut4_0_sram_inv[11] , 
        frac_lut4_0_sram_inv[12] , frac_lut4_0_sram_inv[13] , 
        frac_lut4_0_sram_inv[14] , frac_lut4_0_sram_inv[15] , 
        SYNOPSYS_UNCONNECTED_2 } ) ) ;
endmodule


module logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_4 ( 
    prog_clk , frac_logic_in , ccff_head , frac_logic_out , ccff_tail , p0 ) ;
input  [0:0] prog_clk ;
input  [0:3] frac_logic_in ;
input  [0:0] ccff_head ;
output [0:1] frac_logic_out ;
output [0:0] ccff_tail ;
input  p0 ;

wire [0:0] logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_ccff_tail ;
wire [0:0] logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_frac_lut4_lut3_out ;
wire [0:0] logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_frac_lut4_lut4_out ;
wire [0:1] mux_tree_size2_0_sram ;
wire [0:1] mux_tree_size2_0_sram_inv ;

logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_4 logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0 ( 
    .prog_clk ( prog_clk ) , .frac_lut4_in ( frac_logic_in ) , 
    .ccff_head ( ccff_head ) ,
    .frac_lut4_lut3_out ( { 
        logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_frac_lut4_lut3_out[0] , 
        frac_logic_out[1] } ) ,
    
    .frac_lut4_lut4_out ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_frac_lut4_lut4_out ) , 
    .ccff_tail ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_ccff_tail ) ) ;
mux_tree_size2_28 mux_frac_logic_out_0 (
    .in ( { 
        logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_frac_lut4_lut4_out[0] , 
        logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_frac_lut4_lut3_out[0]
         } ) ,
    .sram ( mux_tree_size2_0_sram ) , 
    .sram_inv ( mux_tree_size2_0_sram_inv ) , .out ( frac_logic_out[0] ) , 
    .p0 ( p0 ) ) ;
mux_tree_size2_mem_28 mem_frac_logic_out_0 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_ccff_tail ) , 
    .ccff_tail ( ccff_tail ) , .mem_out ( mux_tree_size2_0_sram ) , 
    .mem_outb ( mux_tree_size2_0_sram_inv ) ) ;
direct_interc direct_interc_0_ (
    .in ( { SYNOPSYS_UNCONNECTED_1 } ) ,
    .out ( frac_logic_out[1] ) ) ;
direct_interc direct_interc_1_ (
    .in ( { SYNOPSYS_UNCONNECTED_2 } ) ,
    .out ( frac_logic_in[0] ) ) ;
direct_interc direct_interc_2_ (
    .in ( { SYNOPSYS_UNCONNECTED_3 } ) ,
    .out ( frac_logic_in[1] ) ) ;
direct_interc direct_interc_3_ (
    .in ( { SYNOPSYS_UNCONNECTED_4 } ) ,
    .out ( frac_logic_in[2] ) ) ;
direct_interc direct_interc_4_ (
    .in ( { SYNOPSYS_UNCONNECTED_5 } ) ,
    .out ( frac_logic_in[3] ) ) ;
endmodule


module logical_tile_clb_mode_default__fle_mode_physical__fabric_4 ( prog_clk , 
    Test_en , clk , fabric_in , fabric_regin , fabric_scin , fabric_clk , 
    ccff_head , fabric_out , fabric_regout , fabric_scout , ccff_tail , p0 , 
    p2 ) ;
input  [0:0] prog_clk ;
input  [0:0] Test_en ;
input  [0:0] clk ;
input  [0:3] fabric_in ;
input  [0:0] fabric_regin ;
input  [0:0] fabric_scin ;
input  [0:0] fabric_clk ;
input  [0:0] ccff_head ;
output [0:1] fabric_out ;
output [0:0] fabric_regout ;
output [0:0] fabric_scout ;
output [0:0] ccff_tail ;
input  p0 ;
input  p2 ;

wire [0:0] logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0_ff_Q ;
wire [0:0] logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_ccff_tail ;
wire [0:1] logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_frac_logic_out ;
wire [0:1] mux_tree_size2_0_sram ;
wire [0:1] mux_tree_size2_0_sram_inv ;
wire [0:1] mux_tree_size2_1_sram ;
wire [0:1] mux_tree_size2_1_sram_inv ;
wire [0:0] mux_tree_size2_2_out ;
wire [0:1] mux_tree_size2_2_sram ;
wire [0:1] mux_tree_size2_2_sram_inv ;
wire [0:0] mux_tree_size2_mem_0_ccff_tail ;
wire [0:0] mux_tree_size2_mem_1_ccff_tail ;

assign fabric_regout[0] = fabric_scout[0] ;

logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_4 logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0 ( 
    .prog_clk ( prog_clk ) , .frac_logic_in ( fabric_in ) , 
    .ccff_head ( ccff_head ) , 
    .frac_logic_out ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_frac_logic_out ) , 
    .ccff_tail ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_ccff_tail ) , 
    .p0 ( p0 ) ) ;
logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_8 logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0 ( 
    .Test_en ( Test_en ) , .clk ( clk ) , .ff_D ( mux_tree_size2_2_out ) , 
    .ff_DI ( fabric_scin ) , 
    .ff_Q ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0_ff_Q ) ,
    .ff_clk ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_9 logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1 ( 
    .Test_en ( Test_en ) , .clk ( clk ) , 
    .ff_D ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_frac_logic_out[1] ) , 
    .ff_DI ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0_ff_Q ) , 
    .ff_Q ( fabric_scout ) ,
    .ff_clk ( { SYNOPSYS_UNCONNECTED_2 } ) ) ;
mux_tree_size2_12 mux_fabric_out_0 (
    .in ( { 
        logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0_ff_Q[0] , 
        logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_frac_logic_out[0]
         } ) ,
    .sram ( mux_tree_size2_0_sram ) , 
    .sram_inv ( mux_tree_size2_0_sram_inv ) , .out ( fabric_out[0] ) , 
    .p2 ( p2 ) ) ;
mux_tree_size2_13 mux_fabric_out_1 (
    .in ( { fabric_scout[0] , 
        logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_frac_logic_out[1]
         } ) ,
    .sram ( mux_tree_size2_1_sram ) , 
    .sram_inv ( mux_tree_size2_1_sram_inv ) , .out ( fabric_out[1] ) , 
    .p2 ( p2 ) ) ;
mux_tree_size2_14 mux_ff_0_D_0 (
    .in ( { 
        logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_frac_logic_out[0] , 
        fabric_regin[0] } ) ,
    .sram ( mux_tree_size2_2_sram ) , 
    .sram_inv ( mux_tree_size2_2_sram_inv ) , .out ( mux_tree_size2_2_out ) , 
    .p0 ( p0 ) ) ;
mux_tree_size2_mem_12 mem_fabric_out_0 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_size2_mem_0_ccff_tail ) , 
    .mem_out ( mux_tree_size2_0_sram ) , 
    .mem_outb ( mux_tree_size2_0_sram_inv ) ) ;
mux_tree_size2_mem_13 mem_fabric_out_1 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_size2_mem_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_size2_mem_1_ccff_tail ) , 
    .mem_out ( mux_tree_size2_1_sram ) , 
    .mem_outb ( mux_tree_size2_1_sram_inv ) ) ;
mux_tree_size2_mem_14 mem_ff_0_D_0 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_size2_mem_1_ccff_tail ) , .ccff_tail ( ccff_tail ) , 
    .mem_out ( mux_tree_size2_2_sram ) , 
    .mem_outb ( mux_tree_size2_2_sram_inv ) ) ;
direct_interc direct_interc_0_ (
    .in ( { SYNOPSYS_UNCONNECTED_3 } ) ,
    .out ( fabric_scout ) ) ;
direct_interc direct_interc_1_ (
    .in ( { SYNOPSYS_UNCONNECTED_4 } ) ,
    .out ( fabric_scout ) ) ;
direct_interc direct_interc_2_ (
    .in ( { SYNOPSYS_UNCONNECTED_5 } ) ,
    .out ( fabric_in[0] ) ) ;
direct_interc direct_interc_3_ (
    .in ( { SYNOPSYS_UNCONNECTED_6 } ) ,
    .out ( fabric_in[1] ) ) ;
direct_interc direct_interc_4_ (
    .in ( { SYNOPSYS_UNCONNECTED_7 } ) ,
    .out ( fabric_in[2] ) ) ;
direct_interc direct_interc_5_ (
    .in ( { SYNOPSYS_UNCONNECTED_8 } ) ,
    .out ( fabric_in[3] ) ) ;
direct_interc direct_interc_6_ (
    .in ( { SYNOPSYS_UNCONNECTED_9 } ) ,
    .out ( fabric_scin ) ) ;
direct_interc direct_interc_7_ (
    .in ( { SYNOPSYS_UNCONNECTED_10 } ) ,
    .out ( fabric_clk ) ) ;
direct_interc direct_interc_8_ (
    .in ( { SYNOPSYS_UNCONNECTED_11 } ) ,
    
    .out ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_frac_logic_out[1] ) ) ;
direct_interc direct_interc_9_ (
    .in ( { SYNOPSYS_UNCONNECTED_12 } ) ,
    
    .out ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0_ff_Q ) ) ;
direct_interc direct_interc_10_ (
    .in ( { SYNOPSYS_UNCONNECTED_13 } ) ,
    .out ( fabric_clk ) ) ;
endmodule


module logical_tile_clb_mode_default__fle_4 ( prog_clk , Test_en , clk , 
    fle_in , fle_regin , fle_scin , fle_clk , ccff_head , fle_out , 
    fle_regout , fle_scout , ccff_tail , p0 , p2 ) ;
input  [0:0] prog_clk ;
input  [0:0] Test_en ;
input  [0:0] clk ;
input  [0:3] fle_in ;
input  [0:0] fle_regin ;
input  [0:0] fle_scin ;
input  [0:0] fle_clk ;
input  [0:0] ccff_head ;
output [0:1] fle_out ;
output [0:0] fle_regout ;
output [0:0] fle_scout ;
output [0:0] ccff_tail ;
input  p0 ;
input  p2 ;

logical_tile_clb_mode_default__fle_mode_physical__fabric_4 logical_tile_clb_mode_default__fle_mode_physical__fabric_0 ( 
    .prog_clk ( prog_clk ) , .Test_en ( Test_en ) , .clk ( clk ) , 
    .fabric_in ( fle_in ) , .fabric_regin ( fle_regin ) , 
    .fabric_scin ( fle_scin ) , .fabric_clk ( fle_clk ) , 
    .ccff_head ( ccff_head ) , .fabric_out ( fle_out ) , 
    .fabric_regout ( fle_regout ) , .fabric_scout ( fle_scout ) , 
    .ccff_tail ( ccff_tail ) , .p0 ( p0 ) , .p2 ( p2 ) ) ;
direct_interc direct_interc_0_ (
    .in ( { SYNOPSYS_UNCONNECTED_1 } ) ,
    .out ( fle_out[0] ) ) ;
direct_interc direct_interc_1_ (
    .in ( { SYNOPSYS_UNCONNECTED_2 } ) ,
    .out ( fle_out[1] ) ) ;
direct_interc direct_interc_2_ (
    .in ( { SYNOPSYS_UNCONNECTED_3 } ) ,
    .out ( fle_regout ) ) ;
direct_interc direct_interc_3_ (
    .in ( { SYNOPSYS_UNCONNECTED_4 } ) ,
    .out ( fle_scout ) ) ;
direct_interc direct_interc_4_ (
    .in ( { SYNOPSYS_UNCONNECTED_5 } ) ,
    .out ( fle_in[0] ) ) ;
direct_interc direct_interc_5_ (
    .in ( { SYNOPSYS_UNCONNECTED_6 } ) ,
    .out ( fle_in[1] ) ) ;
direct_interc direct_interc_6_ (
    .in ( { SYNOPSYS_UNCONNECTED_7 } ) ,
    .out ( fle_in[2] ) ) ;
direct_interc direct_interc_7_ (
    .in ( { SYNOPSYS_UNCONNECTED_8 } ) ,
    .out ( fle_in[3] ) ) ;
direct_interc direct_interc_8_ (
    .in ( { SYNOPSYS_UNCONNECTED_9 } ) ,
    .out ( fle_regin ) ) ;
direct_interc direct_interc_9_ (
    .in ( { SYNOPSYS_UNCONNECTED_10 } ) ,
    .out ( fle_scin ) ) ;
direct_interc direct_interc_10_ (
    .in ( { SYNOPSYS_UNCONNECTED_11 } ) ,
    .out ( fle_clk ) ) ;
endmodule


module mux_tree_size2_mem_11 ( prog_clk , ccff_head , ccff_tail , mem_out , 
    mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_20__35 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_size2_mem_10 ( prog_clk , ccff_head , ccff_tail , mem_out , 
    mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_19__34 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_size2_mem_9 ( prog_clk , ccff_head , ccff_tail , mem_out , 
    mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_18__33 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_15 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_size2_11 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;

const1_15 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , .X ( out[0] ) ) ;
endmodule


module const1_14 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_size2_10 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;

const1_14 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , .X ( out[0] ) ) ;
endmodule


module const1_13 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_size2_9 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;

const1_13 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , .X ( out[0] ) ) ;
endmodule


module logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_7 ( 
    Test_en , clk , ff_D , ff_DI , ff_Q , ff_clk ) ;
input  [0:0] Test_en ;
input  [0:0] clk ;
input  [0:0] ff_D ;
input  [0:0] ff_DI ;
output [0:0] ff_Q ;
input  [0:0] ff_clk ;

sky130_fd_sc_hd__sdfxbp_1 sky130_fd_sc_hd__sdfxbp_1_0_ ( .D ( ff_D[0] ) , 
    .SCD ( ff_DI[0] ) , .SCE ( Test_en[0] ) , .CLK ( clk[0] ) , 
    .Q ( ff_Q[0] ) , .Q_N ( SYNOPSYS_UNCONNECTED_1 ) ) ;
endmodule


module logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_6 ( 
    Test_en , clk , ff_D , ff_DI , ff_Q , ff_clk ) ;
input  [0:0] Test_en ;
input  [0:0] clk ;
input  [0:0] ff_D ;
input  [0:0] ff_DI ;
output [0:0] ff_Q ;
input  [0:0] ff_clk ;

sky130_fd_sc_hd__sdfxbp_1 sky130_fd_sc_hd__sdfxbp_1_0_ ( .D ( ff_D[0] ) , 
    .SCD ( ff_DI[0] ) , .SCE ( Test_en[0] ) , .CLK ( clk[0] ) , 
    .Q ( ff_Q[0] ) , .Q_N ( SYNOPSYS_UNCONNECTED_1 ) ) ;
endmodule


module mux_tree_size2_mem_27 ( prog_clk , ccff_head , ccff_tail , mem_out , 
    mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_17__32 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_12 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_size2_27 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;

const1_12 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , .X ( out[0] ) ) ;
endmodule


module frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem_3 ( prog_clk , ccff_head , 
    ccff_tail , mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:16] mem_out ;
output [0:16] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_4_ ( .D ( mem_out[3] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[4] ) , .Q_N ( mem_outb[4] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_5_ ( .D ( mem_out[4] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[5] ) , .Q_N ( mem_outb[5] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_6_ ( .D ( mem_out[5] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[6] ) , .Q_N ( mem_outb[6] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_7_ ( .D ( mem_out[6] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[7] ) , .Q_N ( mem_outb[7] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_8_ ( .D ( mem_out[7] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[8] ) , .Q_N ( mem_outb[8] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_9_ ( .D ( mem_out[8] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[9] ) , .Q_N ( mem_outb[9] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_10_ ( .D ( mem_out[9] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[10] ) , .Q_N ( mem_outb[10] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_11_ ( .D ( mem_out[10] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[11] ) , .Q_N ( mem_outb[11] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_12_ ( .D ( mem_out[11] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[12] ) , .Q_N ( mem_outb[12] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_13_ ( .D ( mem_out[12] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[13] ) , .Q_N ( mem_outb[13] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_14_ ( .D ( mem_out[13] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[14] ) , .Q_N ( mem_outb[14] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_15_ ( .D ( mem_out[14] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[15] ) , .Q_N ( mem_outb[15] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_16_ ( .D ( mem_out[15] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[16] ) , .Q_N ( \_gOb3_mem_outb[16] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_16__31 ( .A ( mem_out[16] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module frac_lut4_mux_3 ( in , sram , sram_inv , lut3_out , lut4_out ) ;
input  [0:15] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:1] lut3_out ;
output [0:0] lut4_out ;

wire [0:0] sky130_fd_sc_hd__buf_2_3_X ;
wire [0:0] sky130_fd_sc_hd__buf_2_4_X ;
wire [0:0] sky130_fd_sc_hd__buf_2_5_X ;
wire [0:0] sky130_fd_sc_hd__buf_2_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_10_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_11_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_12_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_13_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_14_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_12_X[0] ) , .X ( lut3_out[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_1_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_13_X[0] ) , .X ( lut3_out[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_2_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_14_X[0] ) , .X ( lut4_out[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_3_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .X ( sky130_fd_sc_hd__buf_2_3_X[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_4_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , 
    .X ( sky130_fd_sc_hd__buf_2_4_X[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_5_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_10_X[0] ) , 
    .X ( sky130_fd_sc_hd__buf_2_5_X[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_6_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_11_X[0] ) , 
    .X ( sky130_fd_sc_hd__buf_2_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_3_ ( .A0 ( in[7] ) , .A1 ( in[6] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_4_ ( .A0 ( in[9] ) , .A1 ( in[8] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_5_ ( .A0 ( in[11] ) , .A1 ( in[10] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_6_ ( .A0 ( in[13] ) , .A1 ( in[12] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_7_ ( .A0 ( in[15] ) , .A1 ( in[14] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_10_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_11_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( .A0 ( sky130_fd_sc_hd__buf_2_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__buf_2_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_12_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( .A0 ( sky130_fd_sc_hd__buf_2_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__buf_2_5_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_13_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_13_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_12_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_14_X[0] ) ) ;
endmodule


module frac_lut4_3 ( in , sram , sram_inv , mode , mode_inv , lut3_out , 
    lut4_out ) ;
input  [0:3] in ;
input  [0:15] sram ;
input  [0:15] sram_inv ;
input  [0:0] mode ;
input  [0:0] mode_inv ;
output [0:1] lut3_out ;
output [0:0] lut4_out ;

wire [0:0] sky130_fd_sc_hd__buf_2_0_X ;
wire [0:0] sky130_fd_sc_hd__buf_2_1_X ;
wire [0:0] sky130_fd_sc_hd__buf_2_2_X ;
wire [0:0] sky130_fd_sc_hd__buf_2_3_X ;
wire [0:0] sky130_fd_sc_hd__inv_1_0_Y ;
wire [0:0] sky130_fd_sc_hd__inv_1_1_Y ;
wire [0:0] sky130_fd_sc_hd__inv_1_2_Y ;
wire [0:0] sky130_fd_sc_hd__inv_1_3_Y ;
wire [0:0] sky130_fd_sc_hd__or2_1_0_X ;

sky130_fd_sc_hd__or2_0 sky130_fd_sc_hd__or2_1_0_ ( .A ( mode[0] ) , 
    .B ( in[3] ) , .X ( sky130_fd_sc_hd__or2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__inv_1 sky130_fd_sc_hd__inv_1_0_ ( .A ( in[0] ) , 
    .Y ( sky130_fd_sc_hd__inv_1_0_Y[0] ) ) ;
sky130_fd_sc_hd__inv_1 sky130_fd_sc_hd__inv_1_1_ ( .A ( in[1] ) , 
    .Y ( sky130_fd_sc_hd__inv_1_1_Y[0] ) ) ;
sky130_fd_sc_hd__inv_1 sky130_fd_sc_hd__inv_1_2_ ( .A ( in[2] ) , 
    .Y ( sky130_fd_sc_hd__inv_1_2_Y[0] ) ) ;
sky130_fd_sc_hd__inv_1 sky130_fd_sc_hd__inv_1_3_ ( 
    .A ( sky130_fd_sc_hd__or2_1_0_X[0] ) , 
    .Y ( sky130_fd_sc_hd__inv_1_3_Y[0] ) ) ;
sky130_fd_sc_hd__buf_2 sky130_fd_sc_hd__buf_2_0_ ( .A ( in[0] ) , 
    .X ( sky130_fd_sc_hd__buf_2_0_X[0] ) ) ;
sky130_fd_sc_hd__buf_2 sky130_fd_sc_hd__buf_2_1_ ( .A ( in[1] ) , 
    .X ( sky130_fd_sc_hd__buf_2_1_X[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_2_ ( .A ( in[2] ) , 
    .X ( sky130_fd_sc_hd__buf_2_2_X[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_3_ ( 
    .A ( sky130_fd_sc_hd__or2_1_0_X[0] ) , 
    .X ( sky130_fd_sc_hd__buf_2_3_X[0] ) ) ;
frac_lut4_mux_3 frac_lut4_mux_0_ ( .in ( sram ) ,
    .sram ( { sky130_fd_sc_hd__buf_2_0_X[0] , sky130_fd_sc_hd__buf_2_1_X[0] , 
        sky130_fd_sc_hd__buf_2_2_X[0] , sky130_fd_sc_hd__buf_2_3_X[0] } ) ,
    .sram_inv ( { sky130_fd_sc_hd__inv_1_0_Y[0] , 
        sky130_fd_sc_hd__inv_1_1_Y[0] , sky130_fd_sc_hd__inv_1_2_Y[0] , 
        sky130_fd_sc_hd__inv_1_3_Y[0] } ) ,
    .lut3_out ( lut3_out ) , .lut4_out ( lut4_out ) ) ;
endmodule


module logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_3 ( 
    prog_clk , frac_lut4_in , ccff_head , frac_lut4_lut3_out , 
    frac_lut4_lut4_out , ccff_tail ) ;
input  [0:0] prog_clk ;
input  [0:3] frac_lut4_in ;
input  [0:0] ccff_head ;
output [0:1] frac_lut4_lut3_out ;
output [0:0] frac_lut4_lut4_out ;
output [0:0] ccff_tail ;

wire [0:0] frac_lut4_0_mode ;
wire [0:15] frac_lut4_0_sram ;
wire [0:15] frac_lut4_0_sram_inv ;

frac_lut4_3 frac_lut4_0_ ( .in ( frac_lut4_in ) , .sram ( frac_lut4_0_sram ) , 
    .sram_inv ( frac_lut4_0_sram_inv ) , .mode ( frac_lut4_0_mode ) ,
    .mode_inv ( { SYNOPSYS_UNCONNECTED_1 } ) ,
    .lut3_out ( frac_lut4_lut3_out ) , .lut4_out ( frac_lut4_lut4_out ) ) ;
frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem_3 frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem ( 
    .prog_clk ( prog_clk ) , .ccff_head ( ccff_head ) , 
    .ccff_tail ( ccff_tail ) ,
    .mem_out ( { frac_lut4_0_sram[0] , frac_lut4_0_sram[1] , 
        frac_lut4_0_sram[2] , frac_lut4_0_sram[3] , frac_lut4_0_sram[4] , 
        frac_lut4_0_sram[5] , frac_lut4_0_sram[6] , frac_lut4_0_sram[7] , 
        frac_lut4_0_sram[8] , frac_lut4_0_sram[9] , frac_lut4_0_sram[10] , 
        frac_lut4_0_sram[11] , frac_lut4_0_sram[12] , frac_lut4_0_sram[13] , 
        frac_lut4_0_sram[14] , frac_lut4_0_sram[15] , frac_lut4_0_mode[0] } ) ,
    .mem_outb ( { frac_lut4_0_sram_inv[0] , frac_lut4_0_sram_inv[1] , 
        frac_lut4_0_sram_inv[2] , frac_lut4_0_sram_inv[3] , 
        frac_lut4_0_sram_inv[4] , frac_lut4_0_sram_inv[5] , 
        frac_lut4_0_sram_inv[6] , frac_lut4_0_sram_inv[7] , 
        frac_lut4_0_sram_inv[8] , frac_lut4_0_sram_inv[9] , 
        frac_lut4_0_sram_inv[10] , frac_lut4_0_sram_inv[11] , 
        frac_lut4_0_sram_inv[12] , frac_lut4_0_sram_inv[13] , 
        frac_lut4_0_sram_inv[14] , frac_lut4_0_sram_inv[15] , 
        SYNOPSYS_UNCONNECTED_2 } ) ) ;
endmodule


module logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_3 ( 
    prog_clk , frac_logic_in , ccff_head , frac_logic_out , ccff_tail , p0 ) ;
input  [0:0] prog_clk ;
input  [0:3] frac_logic_in ;
input  [0:0] ccff_head ;
output [0:1] frac_logic_out ;
output [0:0] ccff_tail ;
input  p0 ;

wire [0:0] logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_ccff_tail ;
wire [0:0] logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_frac_lut4_lut3_out ;
wire [0:0] logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_frac_lut4_lut4_out ;
wire [0:1] mux_tree_size2_0_sram ;
wire [0:1] mux_tree_size2_0_sram_inv ;

logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_3 logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0 ( 
    .prog_clk ( prog_clk ) , .frac_lut4_in ( frac_logic_in ) , 
    .ccff_head ( ccff_head ) ,
    .frac_lut4_lut3_out ( { 
        logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_frac_lut4_lut3_out[0] , 
        frac_logic_out[1] } ) ,
    
    .frac_lut4_lut4_out ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_frac_lut4_lut4_out ) , 
    .ccff_tail ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_ccff_tail ) ) ;
mux_tree_size2_27 mux_frac_logic_out_0 (
    .in ( { 
        logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_frac_lut4_lut4_out[0] , 
        logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_frac_lut4_lut3_out[0]
         } ) ,
    .sram ( mux_tree_size2_0_sram ) , 
    .sram_inv ( mux_tree_size2_0_sram_inv ) , .out ( frac_logic_out[0] ) , 
    .p0 ( p0 ) ) ;
mux_tree_size2_mem_27 mem_frac_logic_out_0 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_ccff_tail ) , 
    .ccff_tail ( ccff_tail ) , .mem_out ( mux_tree_size2_0_sram ) , 
    .mem_outb ( mux_tree_size2_0_sram_inv ) ) ;
direct_interc direct_interc_0_ (
    .in ( { SYNOPSYS_UNCONNECTED_1 } ) ,
    .out ( frac_logic_out[1] ) ) ;
direct_interc direct_interc_1_ (
    .in ( { SYNOPSYS_UNCONNECTED_2 } ) ,
    .out ( frac_logic_in[0] ) ) ;
direct_interc direct_interc_2_ (
    .in ( { SYNOPSYS_UNCONNECTED_3 } ) ,
    .out ( frac_logic_in[1] ) ) ;
direct_interc direct_interc_3_ (
    .in ( { SYNOPSYS_UNCONNECTED_4 } ) ,
    .out ( frac_logic_in[2] ) ) ;
direct_interc direct_interc_4_ (
    .in ( { SYNOPSYS_UNCONNECTED_5 } ) ,
    .out ( frac_logic_in[3] ) ) ;
endmodule


module logical_tile_clb_mode_default__fle_mode_physical__fabric_3 ( prog_clk , 
    Test_en , clk , fabric_in , fabric_regin , fabric_scin , fabric_clk , 
    ccff_head , fabric_out , fabric_regout , fabric_scout , ccff_tail , p0 ) ;
input  [0:0] prog_clk ;
input  [0:0] Test_en ;
input  [0:0] clk ;
input  [0:3] fabric_in ;
input  [0:0] fabric_regin ;
input  [0:0] fabric_scin ;
input  [0:0] fabric_clk ;
input  [0:0] ccff_head ;
output [0:1] fabric_out ;
output [0:0] fabric_regout ;
output [0:0] fabric_scout ;
output [0:0] ccff_tail ;
input  p0 ;

wire [0:0] logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0_ff_Q ;
wire [0:0] logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_ccff_tail ;
wire [0:1] logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_frac_logic_out ;
wire [0:1] mux_tree_size2_0_sram ;
wire [0:1] mux_tree_size2_0_sram_inv ;
wire [0:1] mux_tree_size2_1_sram ;
wire [0:1] mux_tree_size2_1_sram_inv ;
wire [0:0] mux_tree_size2_2_out ;
wire [0:1] mux_tree_size2_2_sram ;
wire [0:1] mux_tree_size2_2_sram_inv ;
wire [0:0] mux_tree_size2_mem_0_ccff_tail ;
wire [0:0] mux_tree_size2_mem_1_ccff_tail ;

assign fabric_regout[0] = fabric_scout[0] ;

logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_3 logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0 ( 
    .prog_clk ( prog_clk ) , .frac_logic_in ( fabric_in ) , 
    .ccff_head ( ccff_head ) , 
    .frac_logic_out ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_frac_logic_out ) , 
    .ccff_tail ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_ccff_tail ) , 
    .p0 ( p0 ) ) ;
logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_6 logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0 ( 
    .Test_en ( Test_en ) , .clk ( clk ) , .ff_D ( mux_tree_size2_2_out ) , 
    .ff_DI ( fabric_scin ) , 
    .ff_Q ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0_ff_Q ) ,
    .ff_clk ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_7 logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1 ( 
    .Test_en ( Test_en ) , .clk ( clk ) , 
    .ff_D ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_frac_logic_out[1] ) , 
    .ff_DI ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0_ff_Q ) , 
    .ff_Q ( fabric_scout ) ,
    .ff_clk ( { SYNOPSYS_UNCONNECTED_2 } ) ) ;
mux_tree_size2_9 mux_fabric_out_0 (
    .in ( { 
        logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0_ff_Q[0] , 
        logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_frac_logic_out[0]
         } ) ,
    .sram ( mux_tree_size2_0_sram ) , 
    .sram_inv ( mux_tree_size2_0_sram_inv ) , .out ( fabric_out[0] ) , 
    .p0 ( p0 ) ) ;
mux_tree_size2_10 mux_fabric_out_1 (
    .in ( { fabric_scout[0] , 
        logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_frac_logic_out[1]
         } ) ,
    .sram ( mux_tree_size2_1_sram ) , 
    .sram_inv ( mux_tree_size2_1_sram_inv ) , .out ( fabric_out[1] ) , 
    .p0 ( p0 ) ) ;
mux_tree_size2_11 mux_ff_0_D_0 (
    .in ( { 
        logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_frac_logic_out[0] , 
        fabric_regin[0] } ) ,
    .sram ( mux_tree_size2_2_sram ) , 
    .sram_inv ( mux_tree_size2_2_sram_inv ) , .out ( mux_tree_size2_2_out ) , 
    .p0 ( p0 ) ) ;
mux_tree_size2_mem_9 mem_fabric_out_0 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_size2_mem_0_ccff_tail ) , 
    .mem_out ( mux_tree_size2_0_sram ) , 
    .mem_outb ( mux_tree_size2_0_sram_inv ) ) ;
mux_tree_size2_mem_10 mem_fabric_out_1 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_size2_mem_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_size2_mem_1_ccff_tail ) , 
    .mem_out ( mux_tree_size2_1_sram ) , 
    .mem_outb ( mux_tree_size2_1_sram_inv ) ) ;
mux_tree_size2_mem_11 mem_ff_0_D_0 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_size2_mem_1_ccff_tail ) , .ccff_tail ( ccff_tail ) , 
    .mem_out ( mux_tree_size2_2_sram ) , 
    .mem_outb ( mux_tree_size2_2_sram_inv ) ) ;
direct_interc direct_interc_0_ (
    .in ( { SYNOPSYS_UNCONNECTED_3 } ) ,
    .out ( fabric_scout ) ) ;
direct_interc direct_interc_1_ (
    .in ( { SYNOPSYS_UNCONNECTED_4 } ) ,
    .out ( fabric_scout ) ) ;
direct_interc direct_interc_2_ (
    .in ( { SYNOPSYS_UNCONNECTED_5 } ) ,
    .out ( fabric_in[0] ) ) ;
direct_interc direct_interc_3_ (
    .in ( { SYNOPSYS_UNCONNECTED_6 } ) ,
    .out ( fabric_in[1] ) ) ;
direct_interc direct_interc_4_ (
    .in ( { SYNOPSYS_UNCONNECTED_7 } ) ,
    .out ( fabric_in[2] ) ) ;
direct_interc direct_interc_5_ (
    .in ( { SYNOPSYS_UNCONNECTED_8 } ) ,
    .out ( fabric_in[3] ) ) ;
direct_interc direct_interc_6_ (
    .in ( { SYNOPSYS_UNCONNECTED_9 } ) ,
    .out ( fabric_scin ) ) ;
direct_interc direct_interc_7_ (
    .in ( { SYNOPSYS_UNCONNECTED_10 } ) ,
    .out ( fabric_clk ) ) ;
direct_interc direct_interc_8_ (
    .in ( { SYNOPSYS_UNCONNECTED_11 } ) ,
    
    .out ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_frac_logic_out[1] ) ) ;
direct_interc direct_interc_9_ (
    .in ( { SYNOPSYS_UNCONNECTED_12 } ) ,
    
    .out ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0_ff_Q ) ) ;
direct_interc direct_interc_10_ (
    .in ( { SYNOPSYS_UNCONNECTED_13 } ) ,
    .out ( fabric_clk ) ) ;
endmodule


module logical_tile_clb_mode_default__fle_3 ( prog_clk , Test_en , clk , 
    fle_in , fle_regin , fle_scin , fle_clk , ccff_head , fle_out , 
    fle_regout , fle_scout , ccff_tail , p0 ) ;
input  [0:0] prog_clk ;
input  [0:0] Test_en ;
input  [0:0] clk ;
input  [0:3] fle_in ;
input  [0:0] fle_regin ;
input  [0:0] fle_scin ;
input  [0:0] fle_clk ;
input  [0:0] ccff_head ;
output [0:1] fle_out ;
output [0:0] fle_regout ;
output [0:0] fle_scout ;
output [0:0] ccff_tail ;
input  p0 ;

logical_tile_clb_mode_default__fle_mode_physical__fabric_3 logical_tile_clb_mode_default__fle_mode_physical__fabric_0 ( 
    .prog_clk ( prog_clk ) , .Test_en ( Test_en ) , .clk ( clk ) , 
    .fabric_in ( fle_in ) , .fabric_regin ( fle_regin ) , 
    .fabric_scin ( fle_scin ) , .fabric_clk ( fle_clk ) , 
    .ccff_head ( ccff_head ) , .fabric_out ( fle_out ) , 
    .fabric_regout ( fle_regout ) , .fabric_scout ( fle_scout ) , 
    .ccff_tail ( ccff_tail ) , .p0 ( p0 ) ) ;
direct_interc direct_interc_0_ (
    .in ( { SYNOPSYS_UNCONNECTED_1 } ) ,
    .out ( fle_out[0] ) ) ;
direct_interc direct_interc_1_ (
    .in ( { SYNOPSYS_UNCONNECTED_2 } ) ,
    .out ( fle_out[1] ) ) ;
direct_interc direct_interc_2_ (
    .in ( { SYNOPSYS_UNCONNECTED_3 } ) ,
    .out ( fle_regout ) ) ;
direct_interc direct_interc_3_ (
    .in ( { SYNOPSYS_UNCONNECTED_4 } ) ,
    .out ( fle_scout ) ) ;
direct_interc direct_interc_4_ (
    .in ( { SYNOPSYS_UNCONNECTED_5 } ) ,
    .out ( fle_in[0] ) ) ;
direct_interc direct_interc_5_ (
    .in ( { SYNOPSYS_UNCONNECTED_6 } ) ,
    .out ( fle_in[1] ) ) ;
direct_interc direct_interc_6_ (
    .in ( { SYNOPSYS_UNCONNECTED_7 } ) ,
    .out ( fle_in[2] ) ) ;
direct_interc direct_interc_7_ (
    .in ( { SYNOPSYS_UNCONNECTED_8 } ) ,
    .out ( fle_in[3] ) ) ;
direct_interc direct_interc_8_ (
    .in ( { SYNOPSYS_UNCONNECTED_9 } ) ,
    .out ( fle_regin ) ) ;
direct_interc direct_interc_9_ (
    .in ( { SYNOPSYS_UNCONNECTED_10 } ) ,
    .out ( fle_scin ) ) ;
direct_interc direct_interc_10_ (
    .in ( { SYNOPSYS_UNCONNECTED_11 } ) ,
    .out ( fle_clk ) ) ;
endmodule


module mux_tree_size2_mem_8 ( prog_clk , ccff_head , ccff_tail , mem_out , 
    mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_15__30 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_size2_mem_7 ( prog_clk , ccff_head , ccff_tail , mem_out , 
    mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_14__29 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_size2_mem_6 ( prog_clk , ccff_head , ccff_tail , mem_out , 
    mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_13__28 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_11 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_size2_8 ( in , sram , sram_inv , out , p1 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p1 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;

const1_11 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p1 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , .X ( out[0] ) ) ;
endmodule


module const1_10 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_size2_7 ( in , sram , sram_inv , out , p1 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p1 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;

const1_10 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p1 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , .X ( out[0] ) ) ;
endmodule


module const1_9 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_size2_6 ( in , sram , sram_inv , out , p1 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p1 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;

const1_9 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p1 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , .X ( out[0] ) ) ;
endmodule


module logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_5 ( 
    Test_en , clk , ff_D , ff_DI , ff_Q , ff_clk ) ;
input  [0:0] Test_en ;
input  [0:0] clk ;
input  [0:0] ff_D ;
input  [0:0] ff_DI ;
output [0:0] ff_Q ;
input  [0:0] ff_clk ;

sky130_fd_sc_hd__sdfxbp_1 sky130_fd_sc_hd__sdfxbp_1_0_ ( .D ( ff_D[0] ) , 
    .SCD ( ff_DI[0] ) , .SCE ( Test_en[0] ) , .CLK ( clk[0] ) , 
    .Q ( ff_Q[0] ) , .Q_N ( SYNOPSYS_UNCONNECTED_1 ) ) ;
endmodule


module logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_4 ( 
    Test_en , clk , ff_D , ff_DI , ff_Q , ff_clk ) ;
input  [0:0] Test_en ;
input  [0:0] clk ;
input  [0:0] ff_D ;
input  [0:0] ff_DI ;
output [0:0] ff_Q ;
input  [0:0] ff_clk ;

sky130_fd_sc_hd__sdfxbp_1 sky130_fd_sc_hd__sdfxbp_1_0_ ( .D ( ff_D[0] ) , 
    .SCD ( ff_DI[0] ) , .SCE ( Test_en[0] ) , .CLK ( clk[0] ) , 
    .Q ( ff_Q[0] ) , .Q_N ( SYNOPSYS_UNCONNECTED_1 ) ) ;
endmodule


module mux_tree_size2_mem_26 ( prog_clk , ccff_head , ccff_tail , mem_out , 
    mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_12__27 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_8 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_size2_26 ( in , sram , sram_inv , out , p1 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p1 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;

const1_8 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p1 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , .X ( out[0] ) ) ;
endmodule


module frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem_2 ( prog_clk , ccff_head , 
    ccff_tail , mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:16] mem_out ;
output [0:16] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_4_ ( .D ( mem_out[3] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[4] ) , .Q_N ( mem_outb[4] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_5_ ( .D ( mem_out[4] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[5] ) , .Q_N ( mem_outb[5] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_6_ ( .D ( mem_out[5] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[6] ) , .Q_N ( mem_outb[6] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_7_ ( .D ( mem_out[6] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[7] ) , .Q_N ( mem_outb[7] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_8_ ( .D ( mem_out[7] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[8] ) , .Q_N ( mem_outb[8] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_9_ ( .D ( mem_out[8] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[9] ) , .Q_N ( mem_outb[9] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_10_ ( .D ( mem_out[9] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[10] ) , .Q_N ( mem_outb[10] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_11_ ( .D ( mem_out[10] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[11] ) , .Q_N ( mem_outb[11] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_12_ ( .D ( mem_out[11] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[12] ) , .Q_N ( mem_outb[12] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_13_ ( .D ( mem_out[12] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[13] ) , .Q_N ( mem_outb[13] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_14_ ( .D ( mem_out[13] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[14] ) , .Q_N ( mem_outb[14] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_15_ ( .D ( mem_out[14] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[15] ) , .Q_N ( mem_outb[15] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_16_ ( .D ( mem_out[15] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[16] ) , .Q_N ( \_gOb2_mem_outb[16] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_11__26 ( .A ( mem_out[16] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module frac_lut4_mux_2 ( in , sram , sram_inv , lut3_out , lut4_out ) ;
input  [0:15] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:1] lut3_out ;
output [0:0] lut4_out ;

wire [0:0] sky130_fd_sc_hd__buf_2_3_X ;
wire [0:0] sky130_fd_sc_hd__buf_2_4_X ;
wire [0:0] sky130_fd_sc_hd__buf_2_5_X ;
wire [0:0] sky130_fd_sc_hd__buf_2_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_10_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_11_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_12_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_13_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_14_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_12_X[0] ) , .X ( lut3_out[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_1_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_13_X[0] ) , .X ( lut3_out[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_2_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_14_X[0] ) , .X ( lut4_out[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_3_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .X ( sky130_fd_sc_hd__buf_2_3_X[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_4_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , 
    .X ( sky130_fd_sc_hd__buf_2_4_X[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_5_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_10_X[0] ) , 
    .X ( sky130_fd_sc_hd__buf_2_5_X[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_6_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_11_X[0] ) , 
    .X ( sky130_fd_sc_hd__buf_2_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_3_ ( .A0 ( in[7] ) , .A1 ( in[6] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_4_ ( .A0 ( in[9] ) , .A1 ( in[8] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_5_ ( .A0 ( in[11] ) , .A1 ( in[10] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_6_ ( .A0 ( in[13] ) , .A1 ( in[12] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_7_ ( .A0 ( in[15] ) , .A1 ( in[14] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_10_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_11_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( .A0 ( sky130_fd_sc_hd__buf_2_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__buf_2_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_12_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( .A0 ( sky130_fd_sc_hd__buf_2_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__buf_2_5_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_13_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_13_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_12_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_14_X[0] ) ) ;
endmodule


module frac_lut4_2 ( in , sram , sram_inv , mode , mode_inv , lut3_out , 
    lut4_out ) ;
input  [0:3] in ;
input  [0:15] sram ;
input  [0:15] sram_inv ;
input  [0:0] mode ;
input  [0:0] mode_inv ;
output [0:1] lut3_out ;
output [0:0] lut4_out ;

wire [0:0] sky130_fd_sc_hd__buf_2_0_X ;
wire [0:0] sky130_fd_sc_hd__buf_2_1_X ;
wire [0:0] sky130_fd_sc_hd__buf_2_2_X ;
wire [0:0] sky130_fd_sc_hd__buf_2_3_X ;
wire [0:0] sky130_fd_sc_hd__inv_1_0_Y ;
wire [0:0] sky130_fd_sc_hd__inv_1_1_Y ;
wire [0:0] sky130_fd_sc_hd__inv_1_2_Y ;
wire [0:0] sky130_fd_sc_hd__inv_1_3_Y ;
wire [0:0] sky130_fd_sc_hd__or2_1_0_X ;

sky130_fd_sc_hd__or2_0 sky130_fd_sc_hd__or2_1_0_ ( .A ( mode[0] ) , 
    .B ( in[3] ) , .X ( sky130_fd_sc_hd__or2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__inv_1 sky130_fd_sc_hd__inv_1_0_ ( .A ( in[0] ) , 
    .Y ( sky130_fd_sc_hd__inv_1_0_Y[0] ) ) ;
sky130_fd_sc_hd__inv_1 sky130_fd_sc_hd__inv_1_1_ ( .A ( in[1] ) , 
    .Y ( sky130_fd_sc_hd__inv_1_1_Y[0] ) ) ;
sky130_fd_sc_hd__inv_1 sky130_fd_sc_hd__inv_1_2_ ( .A ( in[2] ) , 
    .Y ( sky130_fd_sc_hd__inv_1_2_Y[0] ) ) ;
sky130_fd_sc_hd__inv_1 sky130_fd_sc_hd__inv_1_3_ ( 
    .A ( sky130_fd_sc_hd__or2_1_0_X[0] ) , 
    .Y ( sky130_fd_sc_hd__inv_1_3_Y[0] ) ) ;
sky130_fd_sc_hd__buf_2 sky130_fd_sc_hd__buf_2_0_ ( .A ( in[0] ) , 
    .X ( sky130_fd_sc_hd__buf_2_0_X[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_1_ ( .A ( in[1] ) , 
    .X ( sky130_fd_sc_hd__buf_2_1_X[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_2_ ( .A ( in[2] ) , 
    .X ( sky130_fd_sc_hd__buf_2_2_X[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_3_ ( 
    .A ( sky130_fd_sc_hd__or2_1_0_X[0] ) , 
    .X ( sky130_fd_sc_hd__buf_2_3_X[0] ) ) ;
frac_lut4_mux_2 frac_lut4_mux_0_ ( .in ( sram ) ,
    .sram ( { sky130_fd_sc_hd__buf_2_0_X[0] , sky130_fd_sc_hd__buf_2_1_X[0] , 
        sky130_fd_sc_hd__buf_2_2_X[0] , sky130_fd_sc_hd__buf_2_3_X[0] } ) ,
    .sram_inv ( { sky130_fd_sc_hd__inv_1_0_Y[0] , 
        sky130_fd_sc_hd__inv_1_1_Y[0] , sky130_fd_sc_hd__inv_1_2_Y[0] , 
        sky130_fd_sc_hd__inv_1_3_Y[0] } ) ,
    .lut3_out ( lut3_out ) , .lut4_out ( lut4_out ) ) ;
endmodule


module logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_2 ( 
    prog_clk , frac_lut4_in , ccff_head , frac_lut4_lut3_out , 
    frac_lut4_lut4_out , ccff_tail ) ;
input  [0:0] prog_clk ;
input  [0:3] frac_lut4_in ;
input  [0:0] ccff_head ;
output [0:1] frac_lut4_lut3_out ;
output [0:0] frac_lut4_lut4_out ;
output [0:0] ccff_tail ;

wire [0:0] frac_lut4_0_mode ;
wire [0:15] frac_lut4_0_sram ;
wire [0:15] frac_lut4_0_sram_inv ;

frac_lut4_2 frac_lut4_0_ ( .in ( frac_lut4_in ) , .sram ( frac_lut4_0_sram ) , 
    .sram_inv ( frac_lut4_0_sram_inv ) , .mode ( frac_lut4_0_mode ) ,
    .mode_inv ( { SYNOPSYS_UNCONNECTED_1 } ) ,
    .lut3_out ( frac_lut4_lut3_out ) , .lut4_out ( frac_lut4_lut4_out ) ) ;
frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem_2 frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem ( 
    .prog_clk ( prog_clk ) , .ccff_head ( ccff_head ) , 
    .ccff_tail ( ccff_tail ) ,
    .mem_out ( { frac_lut4_0_sram[0] , frac_lut4_0_sram[1] , 
        frac_lut4_0_sram[2] , frac_lut4_0_sram[3] , frac_lut4_0_sram[4] , 
        frac_lut4_0_sram[5] , frac_lut4_0_sram[6] , frac_lut4_0_sram[7] , 
        frac_lut4_0_sram[8] , frac_lut4_0_sram[9] , frac_lut4_0_sram[10] , 
        frac_lut4_0_sram[11] , frac_lut4_0_sram[12] , frac_lut4_0_sram[13] , 
        frac_lut4_0_sram[14] , frac_lut4_0_sram[15] , frac_lut4_0_mode[0] } ) ,
    .mem_outb ( { frac_lut4_0_sram_inv[0] , frac_lut4_0_sram_inv[1] , 
        frac_lut4_0_sram_inv[2] , frac_lut4_0_sram_inv[3] , 
        frac_lut4_0_sram_inv[4] , frac_lut4_0_sram_inv[5] , 
        frac_lut4_0_sram_inv[6] , frac_lut4_0_sram_inv[7] , 
        frac_lut4_0_sram_inv[8] , frac_lut4_0_sram_inv[9] , 
        frac_lut4_0_sram_inv[10] , frac_lut4_0_sram_inv[11] , 
        frac_lut4_0_sram_inv[12] , frac_lut4_0_sram_inv[13] , 
        frac_lut4_0_sram_inv[14] , frac_lut4_0_sram_inv[15] , 
        SYNOPSYS_UNCONNECTED_2 } ) ) ;
endmodule


module logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_2 ( 
    prog_clk , frac_logic_in , ccff_head , frac_logic_out , ccff_tail , p1 ) ;
input  [0:0] prog_clk ;
input  [0:3] frac_logic_in ;
input  [0:0] ccff_head ;
output [0:1] frac_logic_out ;
output [0:0] ccff_tail ;
input  p1 ;

wire [0:0] logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_ccff_tail ;
wire [0:0] logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_frac_lut4_lut3_out ;
wire [0:0] logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_frac_lut4_lut4_out ;
wire [0:1] mux_tree_size2_0_sram ;
wire [0:1] mux_tree_size2_0_sram_inv ;

logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_2 logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0 ( 
    .prog_clk ( prog_clk ) , .frac_lut4_in ( frac_logic_in ) , 
    .ccff_head ( ccff_head ) ,
    .frac_lut4_lut3_out ( { 
        logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_frac_lut4_lut3_out[0] , 
        frac_logic_out[1] } ) ,
    
    .frac_lut4_lut4_out ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_frac_lut4_lut4_out ) , 
    .ccff_tail ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_ccff_tail ) ) ;
mux_tree_size2_26 mux_frac_logic_out_0 (
    .in ( { 
        logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_frac_lut4_lut4_out[0] , 
        logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_frac_lut4_lut3_out[0]
         } ) ,
    .sram ( mux_tree_size2_0_sram ) , 
    .sram_inv ( mux_tree_size2_0_sram_inv ) , .out ( frac_logic_out[0] ) , 
    .p1 ( p1 ) ) ;
mux_tree_size2_mem_26 mem_frac_logic_out_0 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_ccff_tail ) , 
    .ccff_tail ( ccff_tail ) , .mem_out ( mux_tree_size2_0_sram ) , 
    .mem_outb ( mux_tree_size2_0_sram_inv ) ) ;
direct_interc direct_interc_0_ (
    .in ( { SYNOPSYS_UNCONNECTED_1 } ) ,
    .out ( frac_logic_out[1] ) ) ;
direct_interc direct_interc_1_ (
    .in ( { SYNOPSYS_UNCONNECTED_2 } ) ,
    .out ( frac_logic_in[0] ) ) ;
direct_interc direct_interc_2_ (
    .in ( { SYNOPSYS_UNCONNECTED_3 } ) ,
    .out ( frac_logic_in[1] ) ) ;
direct_interc direct_interc_3_ (
    .in ( { SYNOPSYS_UNCONNECTED_4 } ) ,
    .out ( frac_logic_in[2] ) ) ;
direct_interc direct_interc_4_ (
    .in ( { SYNOPSYS_UNCONNECTED_5 } ) ,
    .out ( frac_logic_in[3] ) ) ;
endmodule


module logical_tile_clb_mode_default__fle_mode_physical__fabric_2 ( prog_clk , 
    Test_en , clk , fabric_in , fabric_regin , fabric_scin , fabric_clk , 
    ccff_head , fabric_out , fabric_regout , fabric_scout , ccff_tail , p1 ) ;
input  [0:0] prog_clk ;
input  [0:0] Test_en ;
input  [0:0] clk ;
input  [0:3] fabric_in ;
input  [0:0] fabric_regin ;
input  [0:0] fabric_scin ;
input  [0:0] fabric_clk ;
input  [0:0] ccff_head ;
output [0:1] fabric_out ;
output [0:0] fabric_regout ;
output [0:0] fabric_scout ;
output [0:0] ccff_tail ;
input  p1 ;

wire [0:0] logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0_ff_Q ;
wire [0:0] logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_ccff_tail ;
wire [0:1] logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_frac_logic_out ;
wire [0:1] mux_tree_size2_0_sram ;
wire [0:1] mux_tree_size2_0_sram_inv ;
wire [0:1] mux_tree_size2_1_sram ;
wire [0:1] mux_tree_size2_1_sram_inv ;
wire [0:0] mux_tree_size2_2_out ;
wire [0:1] mux_tree_size2_2_sram ;
wire [0:1] mux_tree_size2_2_sram_inv ;
wire [0:0] mux_tree_size2_mem_0_ccff_tail ;
wire [0:0] mux_tree_size2_mem_1_ccff_tail ;

assign fabric_regout[0] = fabric_scout[0] ;

logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_2 logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0 ( 
    .prog_clk ( prog_clk ) , .frac_logic_in ( fabric_in ) , 
    .ccff_head ( ccff_head ) , 
    .frac_logic_out ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_frac_logic_out ) , 
    .ccff_tail ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_ccff_tail ) , 
    .p1 ( p1 ) ) ;
logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_4 logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0 ( 
    .Test_en ( Test_en ) , .clk ( clk ) , .ff_D ( mux_tree_size2_2_out ) , 
    .ff_DI ( fabric_scin ) , 
    .ff_Q ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0_ff_Q ) ,
    .ff_clk ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_5 logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1 ( 
    .Test_en ( Test_en ) , .clk ( clk ) , 
    .ff_D ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_frac_logic_out[1] ) , 
    .ff_DI ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0_ff_Q ) , 
    .ff_Q ( fabric_scout ) ,
    .ff_clk ( { SYNOPSYS_UNCONNECTED_2 } ) ) ;
mux_tree_size2_6 mux_fabric_out_0 (
    .in ( { 
        logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0_ff_Q[0] , 
        logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_frac_logic_out[0]
         } ) ,
    .sram ( mux_tree_size2_0_sram ) , 
    .sram_inv ( mux_tree_size2_0_sram_inv ) , .out ( fabric_out[0] ) , 
    .p1 ( p1 ) ) ;
mux_tree_size2_7 mux_fabric_out_1 (
    .in ( { fabric_scout[0] , 
        logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_frac_logic_out[1]
         } ) ,
    .sram ( mux_tree_size2_1_sram ) , 
    .sram_inv ( mux_tree_size2_1_sram_inv ) , .out ( fabric_out[1] ) , 
    .p1 ( p1 ) ) ;
mux_tree_size2_8 mux_ff_0_D_0 (
    .in ( { 
        logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_frac_logic_out[0] , 
        fabric_regin[0] } ) ,
    .sram ( mux_tree_size2_2_sram ) , 
    .sram_inv ( mux_tree_size2_2_sram_inv ) , .out ( mux_tree_size2_2_out ) , 
    .p1 ( p1 ) ) ;
mux_tree_size2_mem_6 mem_fabric_out_0 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_size2_mem_0_ccff_tail ) , 
    .mem_out ( mux_tree_size2_0_sram ) , 
    .mem_outb ( mux_tree_size2_0_sram_inv ) ) ;
mux_tree_size2_mem_7 mem_fabric_out_1 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_size2_mem_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_size2_mem_1_ccff_tail ) , 
    .mem_out ( mux_tree_size2_1_sram ) , 
    .mem_outb ( mux_tree_size2_1_sram_inv ) ) ;
mux_tree_size2_mem_8 mem_ff_0_D_0 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_size2_mem_1_ccff_tail ) , .ccff_tail ( ccff_tail ) , 
    .mem_out ( mux_tree_size2_2_sram ) , 
    .mem_outb ( mux_tree_size2_2_sram_inv ) ) ;
direct_interc direct_interc_0_ (
    .in ( { SYNOPSYS_UNCONNECTED_3 } ) ,
    .out ( fabric_scout ) ) ;
direct_interc direct_interc_1_ (
    .in ( { SYNOPSYS_UNCONNECTED_4 } ) ,
    .out ( fabric_scout ) ) ;
direct_interc direct_interc_2_ (
    .in ( { SYNOPSYS_UNCONNECTED_5 } ) ,
    .out ( fabric_in[0] ) ) ;
direct_interc direct_interc_3_ (
    .in ( { SYNOPSYS_UNCONNECTED_6 } ) ,
    .out ( fabric_in[1] ) ) ;
direct_interc direct_interc_4_ (
    .in ( { SYNOPSYS_UNCONNECTED_7 } ) ,
    .out ( fabric_in[2] ) ) ;
direct_interc direct_interc_5_ (
    .in ( { SYNOPSYS_UNCONNECTED_8 } ) ,
    .out ( fabric_in[3] ) ) ;
direct_interc direct_interc_6_ (
    .in ( { SYNOPSYS_UNCONNECTED_9 } ) ,
    .out ( fabric_scin ) ) ;
direct_interc direct_interc_7_ (
    .in ( { SYNOPSYS_UNCONNECTED_10 } ) ,
    .out ( fabric_clk ) ) ;
direct_interc direct_interc_8_ (
    .in ( { SYNOPSYS_UNCONNECTED_11 } ) ,
    
    .out ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_frac_logic_out[1] ) ) ;
direct_interc direct_interc_9_ (
    .in ( { SYNOPSYS_UNCONNECTED_12 } ) ,
    
    .out ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0_ff_Q ) ) ;
direct_interc direct_interc_10_ (
    .in ( { SYNOPSYS_UNCONNECTED_13 } ) ,
    .out ( fabric_clk ) ) ;
endmodule


module logical_tile_clb_mode_default__fle_2 ( prog_clk , Test_en , clk , 
    fle_in , fle_regin , fle_scin , fle_clk , ccff_head , fle_out , 
    fle_regout , fle_scout , ccff_tail , p1 ) ;
input  [0:0] prog_clk ;
input  [0:0] Test_en ;
input  [0:0] clk ;
input  [0:3] fle_in ;
input  [0:0] fle_regin ;
input  [0:0] fle_scin ;
input  [0:0] fle_clk ;
input  [0:0] ccff_head ;
output [0:1] fle_out ;
output [0:0] fle_regout ;
output [0:0] fle_scout ;
output [0:0] ccff_tail ;
input  p1 ;

logical_tile_clb_mode_default__fle_mode_physical__fabric_2 logical_tile_clb_mode_default__fle_mode_physical__fabric_0 ( 
    .prog_clk ( prog_clk ) , .Test_en ( Test_en ) , .clk ( clk ) , 
    .fabric_in ( fle_in ) , .fabric_regin ( fle_regin ) , 
    .fabric_scin ( fle_scin ) , .fabric_clk ( fle_clk ) , 
    .ccff_head ( ccff_head ) , .fabric_out ( fle_out ) , 
    .fabric_regout ( fle_regout ) , .fabric_scout ( fle_scout ) , 
    .ccff_tail ( ccff_tail ) , .p1 ( p1 ) ) ;
direct_interc direct_interc_0_ (
    .in ( { SYNOPSYS_UNCONNECTED_1 } ) ,
    .out ( fle_out[0] ) ) ;
direct_interc direct_interc_1_ (
    .in ( { SYNOPSYS_UNCONNECTED_2 } ) ,
    .out ( fle_out[1] ) ) ;
direct_interc direct_interc_2_ (
    .in ( { SYNOPSYS_UNCONNECTED_3 } ) ,
    .out ( fle_regout ) ) ;
direct_interc direct_interc_3_ (
    .in ( { SYNOPSYS_UNCONNECTED_4 } ) ,
    .out ( fle_scout ) ) ;
direct_interc direct_interc_4_ (
    .in ( { SYNOPSYS_UNCONNECTED_5 } ) ,
    .out ( fle_in[0] ) ) ;
direct_interc direct_interc_5_ (
    .in ( { SYNOPSYS_UNCONNECTED_6 } ) ,
    .out ( fle_in[1] ) ) ;
direct_interc direct_interc_6_ (
    .in ( { SYNOPSYS_UNCONNECTED_7 } ) ,
    .out ( fle_in[2] ) ) ;
direct_interc direct_interc_7_ (
    .in ( { SYNOPSYS_UNCONNECTED_8 } ) ,
    .out ( fle_in[3] ) ) ;
direct_interc direct_interc_8_ (
    .in ( { SYNOPSYS_UNCONNECTED_9 } ) ,
    .out ( fle_regin ) ) ;
direct_interc direct_interc_9_ (
    .in ( { SYNOPSYS_UNCONNECTED_10 } ) ,
    .out ( fle_scin ) ) ;
direct_interc direct_interc_10_ (
    .in ( { SYNOPSYS_UNCONNECTED_11 } ) ,
    .out ( fle_clk ) ) ;
endmodule


module mux_tree_size2_mem_5 ( prog_clk , ccff_head , ccff_tail , mem_out , 
    mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_10__25 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_size2_mem_4 ( prog_clk , ccff_head , ccff_tail , mem_out , 
    mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_9__24 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_size2_mem_3 ( prog_clk , ccff_head , ccff_tail , mem_out , 
    mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_8__23 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_7 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_size2_5 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;

const1_7 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , .X ( out[0] ) ) ;
endmodule


module const1_6 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_size2_4 ( in , sram , sram_inv , out , p1 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p1 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;

const1_6 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p1 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , .X ( out[0] ) ) ;
endmodule


module const1_5 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_size2_3 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;

const1_5 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , .X ( out[0] ) ) ;
endmodule


module logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_3 ( 
    Test_en , clk , ff_D , ff_DI , ff_Q , ff_clk ) ;
input  [0:0] Test_en ;
input  [0:0] clk ;
input  [0:0] ff_D ;
input  [0:0] ff_DI ;
output [0:0] ff_Q ;
input  [0:0] ff_clk ;

sky130_fd_sc_hd__sdfxbp_1 sky130_fd_sc_hd__sdfxbp_1_0_ ( .D ( ff_D[0] ) , 
    .SCD ( ff_DI[0] ) , .SCE ( Test_en[0] ) , .CLK ( clk[0] ) , 
    .Q ( ff_Q[0] ) , .Q_N ( SYNOPSYS_UNCONNECTED_1 ) ) ;
endmodule


module logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_2 ( 
    Test_en , clk , ff_D , ff_DI , ff_Q , ff_clk ) ;
input  [0:0] Test_en ;
input  [0:0] clk ;
input  [0:0] ff_D ;
input  [0:0] ff_DI ;
output [0:0] ff_Q ;
input  [0:0] ff_clk ;

sky130_fd_sc_hd__sdfxbp_1 sky130_fd_sc_hd__sdfxbp_1_0_ ( .D ( ff_D[0] ) , 
    .SCD ( ff_DI[0] ) , .SCE ( Test_en[0] ) , .CLK ( clk[0] ) , 
    .Q ( ff_Q[0] ) , .Q_N ( SYNOPSYS_UNCONNECTED_1 ) ) ;
endmodule


module mux_tree_size2_mem_25 ( prog_clk , ccff_head , ccff_tail , mem_out , 
    mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_7__22 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_4 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_size2_25 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;

const1_4 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , .X ( out[0] ) ) ;
endmodule


module frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem_1 ( prog_clk , ccff_head , 
    ccff_tail , mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:16] mem_out ;
output [0:16] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_4_ ( .D ( mem_out[3] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[4] ) , .Q_N ( mem_outb[4] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_5_ ( .D ( mem_out[4] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[5] ) , .Q_N ( mem_outb[5] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_6_ ( .D ( mem_out[5] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[6] ) , .Q_N ( mem_outb[6] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_7_ ( .D ( mem_out[6] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[7] ) , .Q_N ( mem_outb[7] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_8_ ( .D ( mem_out[7] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[8] ) , .Q_N ( mem_outb[8] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_9_ ( .D ( mem_out[8] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[9] ) , .Q_N ( mem_outb[9] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_10_ ( .D ( mem_out[9] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[10] ) , .Q_N ( mem_outb[10] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_11_ ( .D ( mem_out[10] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[11] ) , .Q_N ( mem_outb[11] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_12_ ( .D ( mem_out[11] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[12] ) , .Q_N ( mem_outb[12] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_13_ ( .D ( mem_out[12] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[13] ) , .Q_N ( mem_outb[13] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_14_ ( .D ( mem_out[13] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[14] ) , .Q_N ( mem_outb[14] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_15_ ( .D ( mem_out[14] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[15] ) , .Q_N ( mem_outb[15] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_16_ ( .D ( mem_out[15] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[16] ) , .Q_N ( \_gOb1_mem_outb[16] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_6__21 ( .A ( mem_out[16] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module frac_lut4_mux_1 ( in , sram , sram_inv , lut3_out , lut4_out ) ;
input  [0:15] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:1] lut3_out ;
output [0:0] lut4_out ;

wire [0:0] sky130_fd_sc_hd__buf_2_3_X ;
wire [0:0] sky130_fd_sc_hd__buf_2_4_X ;
wire [0:0] sky130_fd_sc_hd__buf_2_5_X ;
wire [0:0] sky130_fd_sc_hd__buf_2_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_10_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_11_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_12_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_13_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_14_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_12_X[0] ) , .X ( lut3_out[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_1_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_13_X[0] ) , .X ( lut3_out[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_2_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_14_X[0] ) , .X ( lut4_out[0] ) ) ;
sky130_fd_sc_hd__buf_2 sky130_fd_sc_hd__buf_2_3_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .X ( sky130_fd_sc_hd__buf_2_3_X[0] ) ) ;
sky130_fd_sc_hd__buf_2 sky130_fd_sc_hd__buf_2_4_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , 
    .X ( sky130_fd_sc_hd__buf_2_4_X[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_5_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_10_X[0] ) , 
    .X ( sky130_fd_sc_hd__buf_2_5_X[0] ) ) ;
sky130_fd_sc_hd__buf_2 sky130_fd_sc_hd__buf_2_6_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_11_X[0] ) , 
    .X ( sky130_fd_sc_hd__buf_2_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_3_ ( .A0 ( in[7] ) , .A1 ( in[6] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_4_ ( .A0 ( in[9] ) , .A1 ( in[8] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_5_ ( .A0 ( in[11] ) , .A1 ( in[10] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_6_ ( .A0 ( in[13] ) , .A1 ( in[12] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_7_ ( .A0 ( in[15] ) , .A1 ( in[14] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_10_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_11_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( .A0 ( sky130_fd_sc_hd__buf_2_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__buf_2_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_12_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( .A0 ( sky130_fd_sc_hd__buf_2_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__buf_2_5_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_13_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_13_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_12_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_14_X[0] ) ) ;
endmodule


module frac_lut4_1 ( in , sram , sram_inv , mode , mode_inv , lut3_out , 
    lut4_out ) ;
input  [0:3] in ;
input  [0:15] sram ;
input  [0:15] sram_inv ;
input  [0:0] mode ;
input  [0:0] mode_inv ;
output [0:1] lut3_out ;
output [0:0] lut4_out ;

wire [0:0] sky130_fd_sc_hd__buf_2_0_X ;
wire [0:0] sky130_fd_sc_hd__buf_2_1_X ;
wire [0:0] sky130_fd_sc_hd__buf_2_2_X ;
wire [0:0] sky130_fd_sc_hd__buf_2_3_X ;
wire [0:0] sky130_fd_sc_hd__inv_1_0_Y ;
wire [0:0] sky130_fd_sc_hd__inv_1_1_Y ;
wire [0:0] sky130_fd_sc_hd__inv_1_2_Y ;
wire [0:0] sky130_fd_sc_hd__inv_1_3_Y ;
wire [0:0] sky130_fd_sc_hd__or2_1_0_X ;

sky130_fd_sc_hd__or2_0 sky130_fd_sc_hd__or2_1_0_ ( .A ( mode[0] ) , 
    .B ( in[3] ) , .X ( sky130_fd_sc_hd__or2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__inv_1 sky130_fd_sc_hd__inv_1_0_ ( .A ( in[0] ) , 
    .Y ( sky130_fd_sc_hd__inv_1_0_Y[0] ) ) ;
sky130_fd_sc_hd__inv_1 sky130_fd_sc_hd__inv_1_1_ ( .A ( in[1] ) , 
    .Y ( sky130_fd_sc_hd__inv_1_1_Y[0] ) ) ;
sky130_fd_sc_hd__inv_1 sky130_fd_sc_hd__inv_1_2_ ( .A ( in[2] ) , 
    .Y ( sky130_fd_sc_hd__inv_1_2_Y[0] ) ) ;
sky130_fd_sc_hd__inv_1 sky130_fd_sc_hd__inv_1_3_ ( 
    .A ( sky130_fd_sc_hd__or2_1_0_X[0] ) , 
    .Y ( sky130_fd_sc_hd__inv_1_3_Y[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_0_ ( .A ( in[0] ) , 
    .X ( sky130_fd_sc_hd__buf_2_0_X[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_1_ ( .A ( in[1] ) , 
    .X ( sky130_fd_sc_hd__buf_2_1_X[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_2_ ( .A ( in[2] ) , 
    .X ( sky130_fd_sc_hd__buf_2_2_X[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_3_ ( 
    .A ( sky130_fd_sc_hd__or2_1_0_X[0] ) , 
    .X ( sky130_fd_sc_hd__buf_2_3_X[0] ) ) ;
frac_lut4_mux_1 frac_lut4_mux_0_ ( .in ( sram ) ,
    .sram ( { sky130_fd_sc_hd__buf_2_0_X[0] , sky130_fd_sc_hd__buf_2_1_X[0] , 
        sky130_fd_sc_hd__buf_2_2_X[0] , sky130_fd_sc_hd__buf_2_3_X[0] } ) ,
    .sram_inv ( { sky130_fd_sc_hd__inv_1_0_Y[0] , 
        sky130_fd_sc_hd__inv_1_1_Y[0] , sky130_fd_sc_hd__inv_1_2_Y[0] , 
        sky130_fd_sc_hd__inv_1_3_Y[0] } ) ,
    .lut3_out ( lut3_out ) , .lut4_out ( lut4_out ) ) ;
endmodule


module logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_1 ( 
    prog_clk , frac_lut4_in , ccff_head , frac_lut4_lut3_out , 
    frac_lut4_lut4_out , ccff_tail ) ;
input  [0:0] prog_clk ;
input  [0:3] frac_lut4_in ;
input  [0:0] ccff_head ;
output [0:1] frac_lut4_lut3_out ;
output [0:0] frac_lut4_lut4_out ;
output [0:0] ccff_tail ;

wire [0:0] frac_lut4_0_mode ;
wire [0:15] frac_lut4_0_sram ;
wire [0:15] frac_lut4_0_sram_inv ;

frac_lut4_1 frac_lut4_0_ ( .in ( frac_lut4_in ) , .sram ( frac_lut4_0_sram ) , 
    .sram_inv ( frac_lut4_0_sram_inv ) , .mode ( frac_lut4_0_mode ) ,
    .mode_inv ( { SYNOPSYS_UNCONNECTED_1 } ) ,
    .lut3_out ( frac_lut4_lut3_out ) , .lut4_out ( frac_lut4_lut4_out ) ) ;
frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem_1 frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem ( 
    .prog_clk ( prog_clk ) , .ccff_head ( ccff_head ) , 
    .ccff_tail ( ccff_tail ) ,
    .mem_out ( { frac_lut4_0_sram[0] , frac_lut4_0_sram[1] , 
        frac_lut4_0_sram[2] , frac_lut4_0_sram[3] , frac_lut4_0_sram[4] , 
        frac_lut4_0_sram[5] , frac_lut4_0_sram[6] , frac_lut4_0_sram[7] , 
        frac_lut4_0_sram[8] , frac_lut4_0_sram[9] , frac_lut4_0_sram[10] , 
        frac_lut4_0_sram[11] , frac_lut4_0_sram[12] , frac_lut4_0_sram[13] , 
        frac_lut4_0_sram[14] , frac_lut4_0_sram[15] , frac_lut4_0_mode[0] } ) ,
    .mem_outb ( { frac_lut4_0_sram_inv[0] , frac_lut4_0_sram_inv[1] , 
        frac_lut4_0_sram_inv[2] , frac_lut4_0_sram_inv[3] , 
        frac_lut4_0_sram_inv[4] , frac_lut4_0_sram_inv[5] , 
        frac_lut4_0_sram_inv[6] , frac_lut4_0_sram_inv[7] , 
        frac_lut4_0_sram_inv[8] , frac_lut4_0_sram_inv[9] , 
        frac_lut4_0_sram_inv[10] , frac_lut4_0_sram_inv[11] , 
        frac_lut4_0_sram_inv[12] , frac_lut4_0_sram_inv[13] , 
        frac_lut4_0_sram_inv[14] , frac_lut4_0_sram_inv[15] , 
        SYNOPSYS_UNCONNECTED_2 } ) ) ;
endmodule


module logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_1 ( 
    prog_clk , frac_logic_in , ccff_head , frac_logic_out , ccff_tail , p0 ) ;
input  [0:0] prog_clk ;
input  [0:3] frac_logic_in ;
input  [0:0] ccff_head ;
output [0:1] frac_logic_out ;
output [0:0] ccff_tail ;
input  p0 ;

wire [0:0] logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_ccff_tail ;
wire [0:0] logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_frac_lut4_lut3_out ;
wire [0:0] logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_frac_lut4_lut4_out ;
wire [0:1] mux_tree_size2_0_sram ;
wire [0:1] mux_tree_size2_0_sram_inv ;

logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_1 logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0 ( 
    .prog_clk ( prog_clk ) , .frac_lut4_in ( frac_logic_in ) , 
    .ccff_head ( ccff_head ) ,
    .frac_lut4_lut3_out ( { 
        logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_frac_lut4_lut3_out[0] , 
        frac_logic_out[1] } ) ,
    
    .frac_lut4_lut4_out ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_frac_lut4_lut4_out ) , 
    .ccff_tail ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_ccff_tail ) ) ;
mux_tree_size2_25 mux_frac_logic_out_0 (
    .in ( { 
        logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_frac_lut4_lut4_out[0] , 
        logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_frac_lut4_lut3_out[0]
         } ) ,
    .sram ( mux_tree_size2_0_sram ) , 
    .sram_inv ( mux_tree_size2_0_sram_inv ) , .out ( frac_logic_out[0] ) , 
    .p0 ( p0 ) ) ;
mux_tree_size2_mem_25 mem_frac_logic_out_0 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_ccff_tail ) , 
    .ccff_tail ( ccff_tail ) , .mem_out ( mux_tree_size2_0_sram ) , 
    .mem_outb ( mux_tree_size2_0_sram_inv ) ) ;
direct_interc direct_interc_0_ (
    .in ( { SYNOPSYS_UNCONNECTED_1 } ) ,
    .out ( frac_logic_out[1] ) ) ;
direct_interc direct_interc_1_ (
    .in ( { SYNOPSYS_UNCONNECTED_2 } ) ,
    .out ( frac_logic_in[0] ) ) ;
direct_interc direct_interc_2_ (
    .in ( { SYNOPSYS_UNCONNECTED_3 } ) ,
    .out ( frac_logic_in[1] ) ) ;
direct_interc direct_interc_3_ (
    .in ( { SYNOPSYS_UNCONNECTED_4 } ) ,
    .out ( frac_logic_in[2] ) ) ;
direct_interc direct_interc_4_ (
    .in ( { SYNOPSYS_UNCONNECTED_5 } ) ,
    .out ( frac_logic_in[3] ) ) ;
endmodule


module logical_tile_clb_mode_default__fle_mode_physical__fabric_1 ( prog_clk , 
    Test_en , clk , fabric_in , fabric_regin , fabric_scin , fabric_clk , 
    ccff_head , fabric_out , fabric_regout , fabric_scout , ccff_tail , p0 , 
    p1 ) ;
input  [0:0] prog_clk ;
input  [0:0] Test_en ;
input  [0:0] clk ;
input  [0:3] fabric_in ;
input  [0:0] fabric_regin ;
input  [0:0] fabric_scin ;
input  [0:0] fabric_clk ;
input  [0:0] ccff_head ;
output [0:1] fabric_out ;
output [0:0] fabric_regout ;
output [0:0] fabric_scout ;
output [0:0] ccff_tail ;
input  p0 ;
input  p1 ;

wire [0:0] logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0_ff_Q ;
wire [0:0] logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_ccff_tail ;
wire [0:1] logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_frac_logic_out ;
wire [0:1] mux_tree_size2_0_sram ;
wire [0:1] mux_tree_size2_0_sram_inv ;
wire [0:1] mux_tree_size2_1_sram ;
wire [0:1] mux_tree_size2_1_sram_inv ;
wire [0:0] mux_tree_size2_2_out ;
wire [0:1] mux_tree_size2_2_sram ;
wire [0:1] mux_tree_size2_2_sram_inv ;
wire [0:0] mux_tree_size2_mem_0_ccff_tail ;
wire [0:0] mux_tree_size2_mem_1_ccff_tail ;

assign fabric_regout[0] = fabric_scout[0] ;

logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_1 logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0 ( 
    .prog_clk ( prog_clk ) , .frac_logic_in ( fabric_in ) , 
    .ccff_head ( ccff_head ) , 
    .frac_logic_out ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_frac_logic_out ) , 
    .ccff_tail ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_ccff_tail ) , 
    .p0 ( p0 ) ) ;
logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_2 logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0 ( 
    .Test_en ( Test_en ) , .clk ( clk ) , .ff_D ( mux_tree_size2_2_out ) , 
    .ff_DI ( fabric_scin ) , 
    .ff_Q ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0_ff_Q ) ,
    .ff_clk ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_3 logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1 ( 
    .Test_en ( Test_en ) , .clk ( clk ) , 
    .ff_D ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_frac_logic_out[1] ) , 
    .ff_DI ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0_ff_Q ) , 
    .ff_Q ( fabric_scout ) ,
    .ff_clk ( { SYNOPSYS_UNCONNECTED_2 } ) ) ;
mux_tree_size2_3 mux_fabric_out_0 (
    .in ( { 
        logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0_ff_Q[0] , 
        logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_frac_logic_out[0]
         } ) ,
    .sram ( mux_tree_size2_0_sram ) , 
    .sram_inv ( mux_tree_size2_0_sram_inv ) , .out ( fabric_out[0] ) , 
    .p0 ( p0 ) ) ;
mux_tree_size2_4 mux_fabric_out_1 (
    .in ( { fabric_scout[0] , 
        logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_frac_logic_out[1]
         } ) ,
    .sram ( mux_tree_size2_1_sram ) , 
    .sram_inv ( mux_tree_size2_1_sram_inv ) , .out ( fabric_out[1] ) , 
    .p1 ( p1 ) ) ;
mux_tree_size2_5 mux_ff_0_D_0 (
    .in ( { 
        logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_frac_logic_out[0] , 
        fabric_regin[0] } ) ,
    .sram ( mux_tree_size2_2_sram ) , 
    .sram_inv ( mux_tree_size2_2_sram_inv ) , .out ( mux_tree_size2_2_out ) , 
    .p0 ( p0 ) ) ;
mux_tree_size2_mem_3 mem_fabric_out_0 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_size2_mem_0_ccff_tail ) , 
    .mem_out ( mux_tree_size2_0_sram ) , 
    .mem_outb ( mux_tree_size2_0_sram_inv ) ) ;
mux_tree_size2_mem_4 mem_fabric_out_1 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_size2_mem_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_size2_mem_1_ccff_tail ) , 
    .mem_out ( mux_tree_size2_1_sram ) , 
    .mem_outb ( mux_tree_size2_1_sram_inv ) ) ;
mux_tree_size2_mem_5 mem_ff_0_D_0 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_size2_mem_1_ccff_tail ) , .ccff_tail ( ccff_tail ) , 
    .mem_out ( mux_tree_size2_2_sram ) , 
    .mem_outb ( mux_tree_size2_2_sram_inv ) ) ;
direct_interc direct_interc_0_ (
    .in ( { SYNOPSYS_UNCONNECTED_3 } ) ,
    .out ( fabric_scout ) ) ;
direct_interc direct_interc_1_ (
    .in ( { SYNOPSYS_UNCONNECTED_4 } ) ,
    .out ( fabric_scout ) ) ;
direct_interc direct_interc_2_ (
    .in ( { SYNOPSYS_UNCONNECTED_5 } ) ,
    .out ( fabric_in[0] ) ) ;
direct_interc direct_interc_3_ (
    .in ( { SYNOPSYS_UNCONNECTED_6 } ) ,
    .out ( fabric_in[1] ) ) ;
direct_interc direct_interc_4_ (
    .in ( { SYNOPSYS_UNCONNECTED_7 } ) ,
    .out ( fabric_in[2] ) ) ;
direct_interc direct_interc_5_ (
    .in ( { SYNOPSYS_UNCONNECTED_8 } ) ,
    .out ( fabric_in[3] ) ) ;
direct_interc direct_interc_6_ (
    .in ( { SYNOPSYS_UNCONNECTED_9 } ) ,
    .out ( fabric_scin ) ) ;
direct_interc direct_interc_7_ (
    .in ( { SYNOPSYS_UNCONNECTED_10 } ) ,
    .out ( fabric_clk ) ) ;
direct_interc direct_interc_8_ (
    .in ( { SYNOPSYS_UNCONNECTED_11 } ) ,
    
    .out ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_frac_logic_out[1] ) ) ;
direct_interc direct_interc_9_ (
    .in ( { SYNOPSYS_UNCONNECTED_12 } ) ,
    
    .out ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0_ff_Q ) ) ;
direct_interc direct_interc_10_ (
    .in ( { SYNOPSYS_UNCONNECTED_13 } ) ,
    .out ( fabric_clk ) ) ;
endmodule


module logical_tile_clb_mode_default__fle_1 ( prog_clk , Test_en , clk , 
    fle_in , fle_regin , fle_scin , fle_clk , ccff_head , fle_out , 
    fle_regout , fle_scout , ccff_tail , p0 , p1 ) ;
input  [0:0] prog_clk ;
input  [0:0] Test_en ;
input  [0:0] clk ;
input  [0:3] fle_in ;
input  [0:0] fle_regin ;
input  [0:0] fle_scin ;
input  [0:0] fle_clk ;
input  [0:0] ccff_head ;
output [0:1] fle_out ;
output [0:0] fle_regout ;
output [0:0] fle_scout ;
output [0:0] ccff_tail ;
input  p0 ;
input  p1 ;

logical_tile_clb_mode_default__fle_mode_physical__fabric_1 logical_tile_clb_mode_default__fle_mode_physical__fabric_0 ( 
    .prog_clk ( prog_clk ) , .Test_en ( Test_en ) , .clk ( clk ) , 
    .fabric_in ( fle_in ) , .fabric_regin ( fle_regin ) , 
    .fabric_scin ( fle_scin ) , .fabric_clk ( fle_clk ) , 
    .ccff_head ( ccff_head ) , .fabric_out ( fle_out ) , 
    .fabric_regout ( fle_regout ) , .fabric_scout ( fle_scout ) , 
    .ccff_tail ( ccff_tail ) , .p0 ( p0 ) , .p1 ( p1 ) ) ;
direct_interc direct_interc_0_ (
    .in ( { SYNOPSYS_UNCONNECTED_1 } ) ,
    .out ( fle_out[0] ) ) ;
direct_interc direct_interc_1_ (
    .in ( { SYNOPSYS_UNCONNECTED_2 } ) ,
    .out ( fle_out[1] ) ) ;
direct_interc direct_interc_2_ (
    .in ( { SYNOPSYS_UNCONNECTED_3 } ) ,
    .out ( fle_regout ) ) ;
direct_interc direct_interc_3_ (
    .in ( { SYNOPSYS_UNCONNECTED_4 } ) ,
    .out ( fle_scout ) ) ;
direct_interc direct_interc_4_ (
    .in ( { SYNOPSYS_UNCONNECTED_5 } ) ,
    .out ( fle_in[0] ) ) ;
direct_interc direct_interc_5_ (
    .in ( { SYNOPSYS_UNCONNECTED_6 } ) ,
    .out ( fle_in[1] ) ) ;
direct_interc direct_interc_6_ (
    .in ( { SYNOPSYS_UNCONNECTED_7 } ) ,
    .out ( fle_in[2] ) ) ;
direct_interc direct_interc_7_ (
    .in ( { SYNOPSYS_UNCONNECTED_8 } ) ,
    .out ( fle_in[3] ) ) ;
direct_interc direct_interc_8_ (
    .in ( { SYNOPSYS_UNCONNECTED_9 } ) ,
    .out ( fle_regin ) ) ;
direct_interc direct_interc_9_ (
    .in ( { SYNOPSYS_UNCONNECTED_10 } ) ,
    .out ( fle_scin ) ) ;
direct_interc direct_interc_10_ (
    .in ( { SYNOPSYS_UNCONNECTED_11 } ) ,
    .out ( fle_clk ) ) ;
endmodule


module mux_tree_size2_mem_2 ( prog_clk , ccff_head , ccff_tail , mem_out , 
    mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_5__20 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_size2_mem_1 ( prog_clk , ccff_head , ccff_tail , mem_out , 
    mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_4__19 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_size2_mem_0 ( prog_clk , ccff_head , ccff_tail , mem_out , 
    mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_3__18 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_3 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_size2_2 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;

const1_3 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , .X ( out[0] ) ) ;
endmodule


module const1_2 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_size2_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;

const1_2 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , .X ( out[0] ) ) ;
endmodule


module const1_1 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_size2_0 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;

const1_1 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , .X ( out[0] ) ) ;
endmodule


module logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1 ( 
    Test_en , clk , ff_D , ff_DI , ff_Q , ff_clk ) ;
input  [0:0] Test_en ;
input  [0:0] clk ;
input  [0:0] ff_D ;
input  [0:0] ff_DI ;
output [0:0] ff_Q ;
input  [0:0] ff_clk ;

sky130_fd_sc_hd__sdfxbp_1 sky130_fd_sc_hd__sdfxbp_1_0_ ( .D ( ff_D[0] ) , 
    .SCD ( ff_DI[0] ) , .SCE ( Test_en[0] ) , .CLK ( clk[0] ) , 
    .Q ( ff_Q[0] ) , .Q_N ( SYNOPSYS_UNCONNECTED_1 ) ) ;
endmodule


module logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0 ( 
    Test_en , clk , ff_D , ff_DI , ff_Q , ff_clk ) ;
input  [0:0] Test_en ;
input  [0:0] clk ;
input  [0:0] ff_D ;
input  [0:0] ff_DI ;
output [0:0] ff_Q ;
input  [0:0] ff_clk ;

sky130_fd_sc_hd__sdfxbp_1 sky130_fd_sc_hd__sdfxbp_1_0_ ( .D ( ff_D[0] ) , 
    .SCD ( ff_DI[0] ) , .SCE ( Test_en[0] ) , .CLK ( clk[0] ) , 
    .Q ( ff_Q[0] ) , .Q_N ( SYNOPSYS_UNCONNECTED_1 ) ) ;
endmodule


module direct_interc ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

assign out[0] = in[0] ;
endmodule


module mux_tree_size2_mem_24 ( prog_clk , ccff_head , ccff_tail , mem_out , 
    mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_2__17 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_0 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_size2_24 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;

const1_0 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , .X ( out[0] ) ) ;
endmodule


module frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem_0 ( prog_clk , ccff_head , 
    ccff_tail , mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:16] mem_out ;
output [0:16] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_4_ ( .D ( mem_out[3] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[4] ) , .Q_N ( mem_outb[4] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_5_ ( .D ( mem_out[4] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[5] ) , .Q_N ( mem_outb[5] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_6_ ( .D ( mem_out[5] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[6] ) , .Q_N ( mem_outb[6] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_7_ ( .D ( mem_out[6] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[7] ) , .Q_N ( mem_outb[7] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_8_ ( .D ( mem_out[7] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[8] ) , .Q_N ( mem_outb[8] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_9_ ( .D ( mem_out[8] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[9] ) , .Q_N ( mem_outb[9] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_10_ ( .D ( mem_out[9] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[10] ) , .Q_N ( mem_outb[10] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_11_ ( .D ( mem_out[10] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[11] ) , .Q_N ( mem_outb[11] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_12_ ( .D ( mem_out[11] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[12] ) , .Q_N ( mem_outb[12] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_13_ ( .D ( mem_out[12] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[13] ) , .Q_N ( mem_outb[13] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_14_ ( .D ( mem_out[13] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[14] ) , .Q_N ( mem_outb[14] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_15_ ( .D ( mem_out[14] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[15] ) , .Q_N ( mem_outb[15] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_16_ ( .D ( mem_out[15] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[16] ) , .Q_N ( \_gOb0_mem_outb[16] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_1__16 ( .A ( mem_out[16] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module frac_lut4_mux_0 ( in , sram , sram_inv , lut3_out , lut4_out ) ;
input  [0:15] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:1] lut3_out ;
output [0:0] lut4_out ;

wire [0:0] sky130_fd_sc_hd__buf_2_3_X ;
wire [0:0] sky130_fd_sc_hd__buf_2_4_X ;
wire [0:0] sky130_fd_sc_hd__buf_2_5_X ;
wire [0:0] sky130_fd_sc_hd__buf_2_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_10_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_11_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_12_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_13_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_14_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_12_X[0] ) , .X ( lut3_out[0] ) ) ;
sky130_fd_sc_hd__buf_2 sky130_fd_sc_hd__buf_2_1_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_13_X[0] ) , .X ( lut3_out[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_2_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_14_X[0] ) , .X ( lut4_out[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_3_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .X ( sky130_fd_sc_hd__buf_2_3_X[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_4_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , 
    .X ( sky130_fd_sc_hd__buf_2_4_X[0] ) ) ;
sky130_fd_sc_hd__buf_2 sky130_fd_sc_hd__buf_2_5_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_10_X[0] ) , 
    .X ( sky130_fd_sc_hd__buf_2_5_X[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_6_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_11_X[0] ) , 
    .X ( sky130_fd_sc_hd__buf_2_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_3_ ( .A0 ( in[7] ) , .A1 ( in[6] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_4_ ( .A0 ( in[9] ) , .A1 ( in[8] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_5_ ( .A0 ( in[11] ) , .A1 ( in[10] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_6_ ( .A0 ( in[13] ) , .A1 ( in[12] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_7_ ( .A0 ( in[15] ) , .A1 ( in[14] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_10_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_11_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( .A0 ( sky130_fd_sc_hd__buf_2_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__buf_2_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_12_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( .A0 ( sky130_fd_sc_hd__buf_2_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__buf_2_5_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_13_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_13_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_12_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_14_X[0] ) ) ;
endmodule


module frac_lut4_0 ( in , sram , sram_inv , mode , mode_inv , lut3_out , 
    lut4_out ) ;
input  [0:3] in ;
input  [0:15] sram ;
input  [0:15] sram_inv ;
input  [0:0] mode ;
input  [0:0] mode_inv ;
output [0:1] lut3_out ;
output [0:0] lut4_out ;

wire [0:0] sky130_fd_sc_hd__buf_2_0_X ;
wire [0:0] sky130_fd_sc_hd__buf_2_1_X ;
wire [0:0] sky130_fd_sc_hd__buf_2_2_X ;
wire [0:0] sky130_fd_sc_hd__buf_2_3_X ;
wire [0:0] sky130_fd_sc_hd__inv_1_0_Y ;
wire [0:0] sky130_fd_sc_hd__inv_1_1_Y ;
wire [0:0] sky130_fd_sc_hd__inv_1_2_Y ;
wire [0:0] sky130_fd_sc_hd__inv_1_3_Y ;
wire [0:0] sky130_fd_sc_hd__or2_1_0_X ;

sky130_fd_sc_hd__or2_0 sky130_fd_sc_hd__or2_1_0_ ( .A ( mode[0] ) , 
    .B ( in[3] ) , .X ( sky130_fd_sc_hd__or2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__inv_1 sky130_fd_sc_hd__inv_1_0_ ( .A ( in[0] ) , 
    .Y ( sky130_fd_sc_hd__inv_1_0_Y[0] ) ) ;
sky130_fd_sc_hd__inv_1 sky130_fd_sc_hd__inv_1_1_ ( .A ( in[1] ) , 
    .Y ( sky130_fd_sc_hd__inv_1_1_Y[0] ) ) ;
sky130_fd_sc_hd__inv_1 sky130_fd_sc_hd__inv_1_2_ ( .A ( in[2] ) , 
    .Y ( sky130_fd_sc_hd__inv_1_2_Y[0] ) ) ;
sky130_fd_sc_hd__inv_1 sky130_fd_sc_hd__inv_1_3_ ( 
    .A ( sky130_fd_sc_hd__or2_1_0_X[0] ) , 
    .Y ( sky130_fd_sc_hd__inv_1_3_Y[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_0_ ( .A ( in[0] ) , 
    .X ( sky130_fd_sc_hd__buf_2_0_X[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_1_ ( .A ( in[1] ) , 
    .X ( sky130_fd_sc_hd__buf_2_1_X[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_2_ ( .A ( in[2] ) , 
    .X ( sky130_fd_sc_hd__buf_2_2_X[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_3_ ( 
    .A ( sky130_fd_sc_hd__or2_1_0_X[0] ) , 
    .X ( sky130_fd_sc_hd__buf_2_3_X[0] ) ) ;
frac_lut4_mux_0 frac_lut4_mux_0_ ( .in ( sram ) ,
    .sram ( { sky130_fd_sc_hd__buf_2_0_X[0] , sky130_fd_sc_hd__buf_2_1_X[0] , 
        sky130_fd_sc_hd__buf_2_2_X[0] , sky130_fd_sc_hd__buf_2_3_X[0] } ) ,
    .sram_inv ( { sky130_fd_sc_hd__inv_1_0_Y[0] , 
        sky130_fd_sc_hd__inv_1_1_Y[0] , sky130_fd_sc_hd__inv_1_2_Y[0] , 
        sky130_fd_sc_hd__inv_1_3_Y[0] } ) ,
    .lut3_out ( lut3_out ) , .lut4_out ( lut4_out ) ) ;
endmodule


module logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0 ( 
    prog_clk , frac_lut4_in , ccff_head , frac_lut4_lut3_out , 
    frac_lut4_lut4_out , ccff_tail ) ;
input  [0:0] prog_clk ;
input  [0:3] frac_lut4_in ;
input  [0:0] ccff_head ;
output [0:1] frac_lut4_lut3_out ;
output [0:0] frac_lut4_lut4_out ;
output [0:0] ccff_tail ;

wire [0:0] frac_lut4_0_mode ;
wire [0:15] frac_lut4_0_sram ;
wire [0:15] frac_lut4_0_sram_inv ;

frac_lut4_0 frac_lut4_0_ ( .in ( frac_lut4_in ) , .sram ( frac_lut4_0_sram ) , 
    .sram_inv ( frac_lut4_0_sram_inv ) , .mode ( frac_lut4_0_mode ) ,
    .mode_inv ( { SYNOPSYS_UNCONNECTED_1 } ) ,
    .lut3_out ( frac_lut4_lut3_out ) , .lut4_out ( frac_lut4_lut4_out ) ) ;
frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem_0 frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem ( 
    .prog_clk ( prog_clk ) , .ccff_head ( ccff_head ) , 
    .ccff_tail ( ccff_tail ) ,
    .mem_out ( { frac_lut4_0_sram[0] , frac_lut4_0_sram[1] , 
        frac_lut4_0_sram[2] , frac_lut4_0_sram[3] , frac_lut4_0_sram[4] , 
        frac_lut4_0_sram[5] , frac_lut4_0_sram[6] , frac_lut4_0_sram[7] , 
        frac_lut4_0_sram[8] , frac_lut4_0_sram[9] , frac_lut4_0_sram[10] , 
        frac_lut4_0_sram[11] , frac_lut4_0_sram[12] , frac_lut4_0_sram[13] , 
        frac_lut4_0_sram[14] , frac_lut4_0_sram[15] , frac_lut4_0_mode[0] } ) ,
    .mem_outb ( { frac_lut4_0_sram_inv[0] , frac_lut4_0_sram_inv[1] , 
        frac_lut4_0_sram_inv[2] , frac_lut4_0_sram_inv[3] , 
        frac_lut4_0_sram_inv[4] , frac_lut4_0_sram_inv[5] , 
        frac_lut4_0_sram_inv[6] , frac_lut4_0_sram_inv[7] , 
        frac_lut4_0_sram_inv[8] , frac_lut4_0_sram_inv[9] , 
        frac_lut4_0_sram_inv[10] , frac_lut4_0_sram_inv[11] , 
        frac_lut4_0_sram_inv[12] , frac_lut4_0_sram_inv[13] , 
        frac_lut4_0_sram_inv[14] , frac_lut4_0_sram_inv[15] , 
        SYNOPSYS_UNCONNECTED_2 } ) ) ;
endmodule


module logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0 ( 
    prog_clk , frac_logic_in , ccff_head , frac_logic_out , ccff_tail , p0 ) ;
input  [0:0] prog_clk ;
input  [0:3] frac_logic_in ;
input  [0:0] ccff_head ;
output [0:1] frac_logic_out ;
output [0:0] ccff_tail ;
input  p0 ;

wire [0:0] logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_ccff_tail ;
wire [0:0] logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_frac_lut4_lut3_out ;
wire [0:0] logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_frac_lut4_lut4_out ;
wire [0:1] mux_tree_size2_0_sram ;
wire [0:1] mux_tree_size2_0_sram_inv ;

logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0 logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0 ( 
    .prog_clk ( prog_clk ) , .frac_lut4_in ( frac_logic_in ) , 
    .ccff_head ( ccff_head ) ,
    .frac_lut4_lut3_out ( { 
        logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_frac_lut4_lut3_out[0] , 
        frac_logic_out[1] } ) ,
    
    .frac_lut4_lut4_out ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_frac_lut4_lut4_out ) , 
    .ccff_tail ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_ccff_tail ) ) ;
mux_tree_size2_24 mux_frac_logic_out_0 (
    .in ( { 
        logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_frac_lut4_lut4_out[0] , 
        logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_frac_lut4_lut3_out[0]
         } ) ,
    .sram ( mux_tree_size2_0_sram ) , 
    .sram_inv ( mux_tree_size2_0_sram_inv ) , .out ( frac_logic_out[0] ) , 
    .p0 ( p0 ) ) ;
mux_tree_size2_mem_24 mem_frac_logic_out_0 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_ccff_tail ) , 
    .ccff_tail ( ccff_tail ) , .mem_out ( mux_tree_size2_0_sram ) , 
    .mem_outb ( mux_tree_size2_0_sram_inv ) ) ;
direct_interc direct_interc_0_ (
    .in ( { SYNOPSYS_UNCONNECTED_1 } ) ,
    .out ( frac_logic_out[1] ) ) ;
direct_interc direct_interc_1_ (
    .in ( { SYNOPSYS_UNCONNECTED_2 } ) ,
    .out ( frac_logic_in[0] ) ) ;
direct_interc direct_interc_2_ (
    .in ( { SYNOPSYS_UNCONNECTED_3 } ) ,
    .out ( frac_logic_in[1] ) ) ;
direct_interc direct_interc_3_ (
    .in ( { SYNOPSYS_UNCONNECTED_4 } ) ,
    .out ( frac_logic_in[2] ) ) ;
direct_interc direct_interc_4_ (
    .in ( { SYNOPSYS_UNCONNECTED_5 } ) ,
    .out ( frac_logic_in[3] ) ) ;
endmodule


module logical_tile_clb_mode_default__fle_mode_physical__fabric_0 ( prog_clk , 
    Test_en , clk , fabric_in , fabric_regin , fabric_scin , fabric_clk , 
    ccff_head , fabric_out , fabric_regout , fabric_scout , ccff_tail , p0 ) ;
input  [0:0] prog_clk ;
input  [0:0] Test_en ;
input  [0:0] clk ;
input  [0:3] fabric_in ;
input  [0:0] fabric_regin ;
input  [0:0] fabric_scin ;
input  [0:0] fabric_clk ;
input  [0:0] ccff_head ;
output [0:1] fabric_out ;
output [0:0] fabric_regout ;
output [0:0] fabric_scout ;
output [0:0] ccff_tail ;
input  p0 ;

wire [0:0] logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0_ff_Q ;
wire [0:0] logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_ccff_tail ;
wire [0:1] logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_frac_logic_out ;
wire [0:1] mux_tree_size2_0_sram ;
wire [0:1] mux_tree_size2_0_sram_inv ;
wire [0:1] mux_tree_size2_1_sram ;
wire [0:1] mux_tree_size2_1_sram_inv ;
wire [0:0] mux_tree_size2_2_out ;
wire [0:1] mux_tree_size2_2_sram ;
wire [0:1] mux_tree_size2_2_sram_inv ;
wire [0:0] mux_tree_size2_mem_0_ccff_tail ;
wire [0:0] mux_tree_size2_mem_1_ccff_tail ;

assign fabric_regout[0] = fabric_scout[0] ;

logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0 logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0 ( 
    .prog_clk ( prog_clk ) , .frac_logic_in ( fabric_in ) , 
    .ccff_head ( ccff_head ) , 
    .frac_logic_out ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_frac_logic_out ) , 
    .ccff_tail ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_ccff_tail ) , 
    .p0 ( p0 ) ) ;
logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0 logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0 ( 
    .Test_en ( Test_en ) , .clk ( clk ) , .ff_D ( mux_tree_size2_2_out ) , 
    .ff_DI ( fabric_scin ) , 
    .ff_Q ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0_ff_Q ) ,
    .ff_clk ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1 logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1 ( 
    .Test_en ( Test_en ) , .clk ( clk ) , 
    .ff_D ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_frac_logic_out[1] ) , 
    .ff_DI ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0_ff_Q ) , 
    .ff_Q ( fabric_scout ) ,
    .ff_clk ( { SYNOPSYS_UNCONNECTED_2 } ) ) ;
mux_tree_size2_0 mux_fabric_out_0 (
    .in ( { 
        logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0_ff_Q[0] , 
        logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_frac_logic_out[0]
         } ) ,
    .sram ( mux_tree_size2_0_sram ) , 
    .sram_inv ( mux_tree_size2_0_sram_inv ) , .out ( fabric_out[0] ) , 
    .p0 ( p0 ) ) ;
mux_tree_size2_1 mux_fabric_out_1 (
    .in ( { fabric_scout[0] , 
        logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_frac_logic_out[1]
         } ) ,
    .sram ( mux_tree_size2_1_sram ) , 
    .sram_inv ( mux_tree_size2_1_sram_inv ) , .out ( fabric_out[1] ) , 
    .p0 ( p0 ) ) ;
mux_tree_size2_2 mux_ff_0_D_0 (
    .in ( { 
        logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_frac_logic_out[0] , 
        fabric_regin[0] } ) ,
    .sram ( mux_tree_size2_2_sram ) , 
    .sram_inv ( mux_tree_size2_2_sram_inv ) , .out ( mux_tree_size2_2_out ) , 
    .p0 ( p0 ) ) ;
mux_tree_size2_mem_0 mem_fabric_out_0 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_size2_mem_0_ccff_tail ) , 
    .mem_out ( mux_tree_size2_0_sram ) , 
    .mem_outb ( mux_tree_size2_0_sram_inv ) ) ;
mux_tree_size2_mem_1 mem_fabric_out_1 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_size2_mem_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_size2_mem_1_ccff_tail ) , 
    .mem_out ( mux_tree_size2_1_sram ) , 
    .mem_outb ( mux_tree_size2_1_sram_inv ) ) ;
mux_tree_size2_mem_2 mem_ff_0_D_0 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_size2_mem_1_ccff_tail ) , .ccff_tail ( ccff_tail ) , 
    .mem_out ( mux_tree_size2_2_sram ) , 
    .mem_outb ( mux_tree_size2_2_sram_inv ) ) ;
direct_interc direct_interc_0_ (
    .in ( { SYNOPSYS_UNCONNECTED_3 } ) ,
    .out ( fabric_scout ) ) ;
direct_interc direct_interc_1_ (
    .in ( { SYNOPSYS_UNCONNECTED_4 } ) ,
    .out ( fabric_scout ) ) ;
direct_interc direct_interc_2_ (
    .in ( { SYNOPSYS_UNCONNECTED_5 } ) ,
    .out ( fabric_in[0] ) ) ;
direct_interc direct_interc_3_ (
    .in ( { SYNOPSYS_UNCONNECTED_6 } ) ,
    .out ( fabric_in[1] ) ) ;
direct_interc direct_interc_4_ (
    .in ( { SYNOPSYS_UNCONNECTED_7 } ) ,
    .out ( fabric_in[2] ) ) ;
direct_interc direct_interc_5_ (
    .in ( { SYNOPSYS_UNCONNECTED_8 } ) ,
    .out ( fabric_in[3] ) ) ;
direct_interc direct_interc_6_ (
    .in ( { SYNOPSYS_UNCONNECTED_9 } ) ,
    .out ( fabric_scin ) ) ;
direct_interc direct_interc_7_ (
    .in ( { SYNOPSYS_UNCONNECTED_10 } ) ,
    .out ( fabric_clk ) ) ;
direct_interc direct_interc_8_ (
    .in ( { SYNOPSYS_UNCONNECTED_11 } ) ,
    
    .out ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_frac_logic_out[1] ) ) ;
direct_interc direct_interc_9_ (
    .in ( { SYNOPSYS_UNCONNECTED_12 } ) ,
    
    .out ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0_ff_Q ) ) ;
direct_interc direct_interc_10_ (
    .in ( { SYNOPSYS_UNCONNECTED_13 } ) ,
    .out ( fabric_clk ) ) ;
endmodule


module logical_tile_clb_mode_default__fle_0 ( prog_clk , Test_en , clk , 
    fle_in , fle_regin , fle_scin , fle_clk , ccff_head , fle_out , 
    fle_regout , fle_scout , ccff_tail , p0 ) ;
input  [0:0] prog_clk ;
input  [0:0] Test_en ;
input  [0:0] clk ;
input  [0:3] fle_in ;
input  [0:0] fle_regin ;
input  [0:0] fle_scin ;
input  [0:0] fle_clk ;
input  [0:0] ccff_head ;
output [0:1] fle_out ;
output [0:0] fle_regout ;
output [0:0] fle_scout ;
output [0:0] ccff_tail ;
input  p0 ;

logical_tile_clb_mode_default__fle_mode_physical__fabric_0 logical_tile_clb_mode_default__fle_mode_physical__fabric_0 ( 
    .prog_clk ( prog_clk ) , .Test_en ( Test_en ) , .clk ( clk ) , 
    .fabric_in ( fle_in ) , .fabric_regin ( fle_regin ) , 
    .fabric_scin ( fle_scin ) , .fabric_clk ( fle_clk ) , 
    .ccff_head ( ccff_head ) , .fabric_out ( fle_out ) , 
    .fabric_regout ( fle_regout ) , .fabric_scout ( fle_scout ) , 
    .ccff_tail ( ccff_tail ) , .p0 ( p0 ) ) ;
direct_interc direct_interc_0_ (
    .in ( { SYNOPSYS_UNCONNECTED_1 } ) ,
    .out ( fle_out[0] ) ) ;
direct_interc direct_interc_1_ (
    .in ( { SYNOPSYS_UNCONNECTED_2 } ) ,
    .out ( fle_out[1] ) ) ;
direct_interc direct_interc_2_ (
    .in ( { SYNOPSYS_UNCONNECTED_3 } ) ,
    .out ( fle_regout ) ) ;
direct_interc direct_interc_3_ (
    .in ( { SYNOPSYS_UNCONNECTED_4 } ) ,
    .out ( fle_scout ) ) ;
direct_interc direct_interc_4_ (
    .in ( { SYNOPSYS_UNCONNECTED_5 } ) ,
    .out ( fle_in[0] ) ) ;
direct_interc direct_interc_5_ (
    .in ( { SYNOPSYS_UNCONNECTED_6 } ) ,
    .out ( fle_in[1] ) ) ;
direct_interc direct_interc_6_ (
    .in ( { SYNOPSYS_UNCONNECTED_7 } ) ,
    .out ( fle_in[2] ) ) ;
direct_interc direct_interc_7_ (
    .in ( { SYNOPSYS_UNCONNECTED_8 } ) ,
    .out ( fle_in[3] ) ) ;
direct_interc direct_interc_8_ (
    .in ( { SYNOPSYS_UNCONNECTED_9 } ) ,
    .out ( fle_regin ) ) ;
direct_interc direct_interc_9_ (
    .in ( { SYNOPSYS_UNCONNECTED_10 } ) ,
    .out ( fle_scin ) ) ;
direct_interc direct_interc_10_ (
    .in ( { SYNOPSYS_UNCONNECTED_11 } ) ,
    .out ( fle_clk ) ) ;
endmodule


module logical_tile_clb_mode_clb_ ( prog_clk , Test_en , clk , clb_I0 , 
    clb_I1 , clb_I2 , clb_I3 , clb_I4 , clb_I5 , clb_I6 , clb_I7 , clb_regin , 
    clb_scin , clb_clk , ccff_head , clb_O , clb_regout , clb_scout , 
    ccff_tail , p_abuf1 , p_abuf2 , p_abuf3 , p_abuf4 , p_abuf5 , p_abuf6 , 
    p_abuf7 , p_abuf8 , p_abuf9 , p_abuf10 , p_abuf11 , p_abuf12 , p_abuf13 , 
    p_abuf14 , p_abuf15 , p0 , p1 , p2 , p3 , p4 ) ;
input  [0:0] prog_clk ;
input  [0:0] Test_en ;
input  [0:0] clk ;
input  [0:3] clb_I0 ;
input  [0:3] clb_I1 ;
input  [0:3] clb_I2 ;
input  [0:3] clb_I3 ;
input  [0:3] clb_I4 ;
input  [0:3] clb_I5 ;
input  [0:3] clb_I6 ;
input  [0:3] clb_I7 ;
input  [0:0] clb_regin ;
input  [0:0] clb_scin ;
input  [0:0] clb_clk ;
input  [0:0] ccff_head ;
output [0:15] clb_O ;
output [0:0] clb_regout ;
output [0:0] clb_scout ;
output [0:0] ccff_tail ;
output p_abuf1 ;
output p_abuf2 ;
output p_abuf3 ;
output p_abuf4 ;
output p_abuf5 ;
output p_abuf6 ;
output p_abuf7 ;
output p_abuf8 ;
output p_abuf9 ;
output p_abuf10 ;
output p_abuf11 ;
output p_abuf12 ;
output p_abuf13 ;
output p_abuf14 ;
output p_abuf15 ;
input  p0 ;
input  p1 ;
input  p2 ;
input  p3 ;
input  p4 ;

wire [0:0] logical_tile_clb_mode_default__fle_0_ccff_tail ;
wire [0:0] logical_tile_clb_mode_default__fle_0_fle_out ;
wire [0:0] logical_tile_clb_mode_default__fle_0_fle_regout ;
wire [0:0] logical_tile_clb_mode_default__fle_0_fle_scout ;
wire [0:0] logical_tile_clb_mode_default__fle_1_ccff_tail ;
wire [0:0] logical_tile_clb_mode_default__fle_1_fle_out ;
wire [0:0] logical_tile_clb_mode_default__fle_1_fle_regout ;
wire [0:0] logical_tile_clb_mode_default__fle_1_fle_scout ;
wire [0:0] logical_tile_clb_mode_default__fle_2_ccff_tail ;
wire [0:0] logical_tile_clb_mode_default__fle_2_fle_regout ;
wire [0:0] logical_tile_clb_mode_default__fle_2_fle_scout ;
wire [0:0] logical_tile_clb_mode_default__fle_3_ccff_tail ;
wire [0:0] logical_tile_clb_mode_default__fle_3_fle_regout ;
wire [0:0] logical_tile_clb_mode_default__fle_3_fle_scout ;
wire [0:0] logical_tile_clb_mode_default__fle_4_ccff_tail ;
wire [0:1] logical_tile_clb_mode_default__fle_4_fle_out ;
wire [0:0] logical_tile_clb_mode_default__fle_4_fle_regout ;
wire [0:0] logical_tile_clb_mode_default__fle_4_fle_scout ;
wire [0:0] logical_tile_clb_mode_default__fle_5_ccff_tail ;
wire [0:0] logical_tile_clb_mode_default__fle_5_fle_regout ;
wire [0:0] logical_tile_clb_mode_default__fle_5_fle_scout ;
wire [0:0] logical_tile_clb_mode_default__fle_6_ccff_tail ;
wire [1:1] logical_tile_clb_mode_default__fle_6_fle_out ;
wire [0:0] logical_tile_clb_mode_default__fle_6_fle_regout ;
wire [0:0] logical_tile_clb_mode_default__fle_6_fle_scout ;
wire [1:1] logical_tile_clb_mode_default__fle_7_fle_out ;

logical_tile_clb_mode_default__fle_0 logical_tile_clb_mode_default__fle_0 ( 
    .prog_clk ( prog_clk ) , .Test_en ( Test_en ) , .clk ( clk ) , 
    .fle_in ( clb_I0 ) , .fle_regin ( clb_regin ) , .fle_scin ( clb_scin ) , 
    .fle_clk ( clb_clk ) , .ccff_head ( ccff_head ) ,
    .fle_out ( { logical_tile_clb_mode_default__fle_0_fle_out[0] , clb_O[0] } ) ,
    .fle_regout ( logical_tile_clb_mode_default__fle_0_fle_regout ) , 
    .fle_scout ( logical_tile_clb_mode_default__fle_0_fle_scout ) , 
    .ccff_tail ( logical_tile_clb_mode_default__fle_0_ccff_tail ) , 
    .p0 ( p1 ) ) ;
logical_tile_clb_mode_default__fle_1 logical_tile_clb_mode_default__fle_1 ( 
    .prog_clk ( prog_clk ) , .Test_en ( Test_en ) , .clk ( clk ) , 
    .fle_in ( clb_I1 ) , 
    .fle_regin ( logical_tile_clb_mode_default__fle_0_fle_regout ) , 
    .fle_scin ( logical_tile_clb_mode_default__fle_0_fle_scout ) , 
    .fle_clk ( clb_clk ) , 
    .ccff_head ( logical_tile_clb_mode_default__fle_0_ccff_tail ) ,
    .fle_out ( { logical_tile_clb_mode_default__fle_1_fle_out[0] , p_abuf3 } ) ,
    .fle_regout ( logical_tile_clb_mode_default__fle_1_fle_regout ) , 
    .fle_scout ( logical_tile_clb_mode_default__fle_1_fle_scout ) , 
    .ccff_tail ( logical_tile_clb_mode_default__fle_1_ccff_tail ) , 
    .p0 ( p0 ) , .p1 ( p2 ) ) ;
logical_tile_clb_mode_default__fle_2 logical_tile_clb_mode_default__fle_2 ( 
    .prog_clk ( prog_clk ) , .Test_en ( Test_en ) , .clk ( clk ) , 
    .fle_in ( clb_I2 ) , 
    .fle_regin ( logical_tile_clb_mode_default__fle_1_fle_regout ) , 
    .fle_scin ( logical_tile_clb_mode_default__fle_1_fle_scout ) , 
    .fle_clk ( clb_clk ) , 
    .ccff_head ( logical_tile_clb_mode_default__fle_1_ccff_tail ) ,
    .fle_out ( { clb_O[5] , p_abuf5 } ) ,
    .fle_regout ( logical_tile_clb_mode_default__fle_2_fle_regout ) , 
    .fle_scout ( logical_tile_clb_mode_default__fle_2_fle_scout ) , 
    .ccff_tail ( logical_tile_clb_mode_default__fle_2_ccff_tail ) , 
    .p1 ( p2 ) ) ;
logical_tile_clb_mode_default__fle_3 logical_tile_clb_mode_default__fle_3 ( 
    .prog_clk ( prog_clk ) , .Test_en ( Test_en ) , .clk ( clk ) , 
    .fle_in ( clb_I3 ) , 
    .fle_regin ( logical_tile_clb_mode_default__fle_2_fle_regout ) , 
    .fle_scin ( logical_tile_clb_mode_default__fle_2_fle_scout ) , 
    .fle_clk ( clb_clk ) , 
    .ccff_head ( logical_tile_clb_mode_default__fle_2_ccff_tail ) ,
    .fle_out ( { clb_O[7] , clb_O[6] } ) ,
    .fle_regout ( logical_tile_clb_mode_default__fle_3_fle_regout ) , 
    .fle_scout ( logical_tile_clb_mode_default__fle_3_fle_scout ) , 
    .ccff_tail ( logical_tile_clb_mode_default__fle_3_ccff_tail ) , 
    .p0 ( p0 ) ) ;
logical_tile_clb_mode_default__fle_4 logical_tile_clb_mode_default__fle_4 ( 
    .prog_clk ( prog_clk ) , .Test_en ( Test_en ) , .clk ( clk ) , 
    .fle_in ( clb_I4 ) , 
    .fle_regin ( logical_tile_clb_mode_default__fle_3_fle_regout ) , 
    .fle_scin ( logical_tile_clb_mode_default__fle_3_fle_scout ) , 
    .fle_clk ( clb_clk ) , 
    .ccff_head ( logical_tile_clb_mode_default__fle_3_ccff_tail ) , 
    .fle_out ( logical_tile_clb_mode_default__fle_4_fle_out ) , 
    .fle_regout ( logical_tile_clb_mode_default__fle_4_fle_regout ) , 
    .fle_scout ( logical_tile_clb_mode_default__fle_4_fle_scout ) , 
    .ccff_tail ( logical_tile_clb_mode_default__fle_4_ccff_tail ) , 
    .p0 ( p0 ) , .p2 ( p3 ) ) ;
logical_tile_clb_mode_default__fle_5 logical_tile_clb_mode_default__fle_5 ( 
    .prog_clk ( prog_clk ) , .Test_en ( Test_en ) , .clk ( clk ) , 
    .fle_in ( clb_I5 ) , 
    .fle_regin ( logical_tile_clb_mode_default__fle_4_fle_regout ) , 
    .fle_scin ( logical_tile_clb_mode_default__fle_4_fle_scout ) , 
    .fle_clk ( clb_clk ) , 
    .ccff_head ( logical_tile_clb_mode_default__fle_4_ccff_tail ) ,
    .fle_out ( { clb_O[11] , clb_O[10] } ) ,
    .fle_regout ( logical_tile_clb_mode_default__fle_5_fle_regout ) , 
    .fle_scout ( logical_tile_clb_mode_default__fle_5_fle_scout ) , 
    .ccff_tail ( logical_tile_clb_mode_default__fle_5_ccff_tail ) , 
    .p2 ( p3 ) ) ;
logical_tile_clb_mode_default__fle_6 logical_tile_clb_mode_default__fle_6 ( 
    .prog_clk ( prog_clk ) , .Test_en ( Test_en ) , .clk ( clk ) , 
    .fle_in ( clb_I6 ) , 
    .fle_regin ( logical_tile_clb_mode_default__fle_5_fle_regout ) , 
    .fle_scin ( logical_tile_clb_mode_default__fle_5_fle_scout ) , 
    .fle_clk ( clb_clk ) , 
    .ccff_head ( logical_tile_clb_mode_default__fle_5_ccff_tail ) ,
    .fle_out ( { clb_O[13] , logical_tile_clb_mode_default__fle_6_fle_out[1] } ) ,
    .fle_regout ( logical_tile_clb_mode_default__fle_6_fle_regout ) , 
    .fle_scout ( logical_tile_clb_mode_default__fle_6_fle_scout ) , 
    .ccff_tail ( logical_tile_clb_mode_default__fle_6_ccff_tail ) , 
    .p2 ( p3 ) , .p3 ( p4 ) ) ;
logical_tile_clb_mode_default__fle logical_tile_clb_mode_default__fle_7 ( 
    .prog_clk ( prog_clk ) , .Test_en ( Test_en ) , .clk ( clk ) , 
    .fle_in ( clb_I7 ) , 
    .fle_regin ( logical_tile_clb_mode_default__fle_6_fle_regout ) , 
    .fle_scin ( logical_tile_clb_mode_default__fle_6_fle_scout ) , 
    .fle_clk ( clb_clk ) , 
    .ccff_head ( logical_tile_clb_mode_default__fle_6_ccff_tail ) ,
    .fle_out ( { clb_O[15] , logical_tile_clb_mode_default__fle_7_fle_out[1] } ) ,
    .fle_regout ( clb_regout ) , .fle_scout ( clb_scout ) , 
    .ccff_tail ( ccff_tail ) , .p_abuf0 ( p_abuf16 ) , .p_abuf1 ( p_abuf17 ) , 
    .p3 ( p4 ) ) ;
direct_interc direct_interc_0_ (
    .in ( { SYNOPSYS_UNCONNECTED_1 } ) ,
    .out ( clb_O[0] ) ) ;
direct_interc direct_interc_1_ (
    .in ( { SYNOPSYS_UNCONNECTED_2 } ) ,
    .out ( logical_tile_clb_mode_default__fle_0_fle_out ) ) ;
direct_interc direct_interc_2_ (
    .in ( { SYNOPSYS_UNCONNECTED_3 } ) ,
    .out ( { p_abuf3 } ) ) ;
direct_interc direct_interc_3_ (
    .in ( { SYNOPSYS_UNCONNECTED_4 } ) ,
    .out ( logical_tile_clb_mode_default__fle_1_fle_out ) ) ;
direct_interc direct_interc_4_ (
    .in ( { SYNOPSYS_UNCONNECTED_5 } ) ,
    .out ( { p_abuf5 } ) ) ;
direct_interc direct_interc_5_ (
    .in ( { SYNOPSYS_UNCONNECTED_6 } ) ,
    .out ( clb_O[5] ) ) ;
direct_interc direct_interc_6_ (
    .in ( { SYNOPSYS_UNCONNECTED_7 } ) ,
    .out ( clb_O[6] ) ) ;
direct_interc direct_interc_7_ (
    .in ( { SYNOPSYS_UNCONNECTED_8 } ) ,
    .out ( clb_O[7] ) ) ;
direct_interc direct_interc_8_ (
    .in ( { SYNOPSYS_UNCONNECTED_9 } ) ,
    .out ( logical_tile_clb_mode_default__fle_4_fle_out[1] ) ) ;
direct_interc direct_interc_9_ (
    .in ( { SYNOPSYS_UNCONNECTED_10 } ) ,
    .out ( logical_tile_clb_mode_default__fle_4_fle_out[0] ) ) ;
direct_interc direct_interc_10_ (
    .in ( { SYNOPSYS_UNCONNECTED_11 } ) ,
    .out ( clb_O[10] ) ) ;
direct_interc direct_interc_11_ (
    .in ( { SYNOPSYS_UNCONNECTED_12 } ) ,
    .out ( clb_O[11] ) ) ;
direct_interc direct_interc_12_ (
    .in ( { SYNOPSYS_UNCONNECTED_13 } ) ,
    .out ( logical_tile_clb_mode_default__fle_6_fle_out ) ) ;
direct_interc direct_interc_13_ (
    .in ( { SYNOPSYS_UNCONNECTED_14 } ) ,
    .out ( clb_O[13] ) ) ;
direct_interc direct_interc_14_ (
    .in ( { SYNOPSYS_UNCONNECTED_15 } ) ,
    .out ( logical_tile_clb_mode_default__fle_7_fle_out ) ) ;
direct_interc direct_interc_15_ (
    .in ( { SYNOPSYS_UNCONNECTED_16 } ) ,
    .out ( clb_O[15] ) ) ;
direct_interc direct_interc_16_ (
    .in ( { SYNOPSYS_UNCONNECTED_17 } ) ,
    .out ( { p_abuf17 } ) ) ;
direct_interc direct_interc_17_ (
    .in ( { SYNOPSYS_UNCONNECTED_18 } ) ,
    .out ( { p_abuf16 } ) ) ;
direct_interc direct_interc_18_ (
    .in ( { SYNOPSYS_UNCONNECTED_19 } ) ,
    .out ( clb_I0[0] ) ) ;
direct_interc direct_interc_19_ (
    .in ( { SYNOPSYS_UNCONNECTED_20 } ) ,
    .out ( clb_I0[1] ) ) ;
direct_interc direct_interc_20_ (
    .in ( { SYNOPSYS_UNCONNECTED_21 } ) ,
    .out ( clb_I0[2] ) ) ;
direct_interc direct_interc_21_ (
    .in ( { SYNOPSYS_UNCONNECTED_22 } ) ,
    .out ( clb_I0[3] ) ) ;
direct_interc direct_interc_22_ (
    .in ( { SYNOPSYS_UNCONNECTED_23 } ) ,
    .out ( clb_regin ) ) ;
direct_interc direct_interc_23_ (
    .in ( { SYNOPSYS_UNCONNECTED_24 } ) ,
    .out ( clb_scin ) ) ;
direct_interc direct_interc_24_ (
    .in ( { SYNOPSYS_UNCONNECTED_25 } ) ,
    .out ( clb_clk ) ) ;
direct_interc direct_interc_25_ (
    .in ( { SYNOPSYS_UNCONNECTED_26 } ) ,
    .out ( clb_I1[0] ) ) ;
direct_interc direct_interc_26_ (
    .in ( { SYNOPSYS_UNCONNECTED_27 } ) ,
    .out ( clb_I1[1] ) ) ;
direct_interc direct_interc_27_ (
    .in ( { SYNOPSYS_UNCONNECTED_28 } ) ,
    .out ( clb_I1[2] ) ) ;
direct_interc direct_interc_28_ (
    .in ( { SYNOPSYS_UNCONNECTED_29 } ) ,
    .out ( clb_I1[3] ) ) ;
direct_interc direct_interc_29_ (
    .in ( { SYNOPSYS_UNCONNECTED_30 } ) ,
    .out ( logical_tile_clb_mode_default__fle_0_fle_regout ) ) ;
direct_interc direct_interc_30_ (
    .in ( { SYNOPSYS_UNCONNECTED_31 } ) ,
    .out ( logical_tile_clb_mode_default__fle_0_fle_scout ) ) ;
direct_interc direct_interc_31_ (
    .in ( { SYNOPSYS_UNCONNECTED_32 } ) ,
    .out ( clb_clk ) ) ;
direct_interc direct_interc_32_ (
    .in ( { SYNOPSYS_UNCONNECTED_33 } ) ,
    .out ( clb_I2[0] ) ) ;
direct_interc direct_interc_33_ (
    .in ( { SYNOPSYS_UNCONNECTED_34 } ) ,
    .out ( clb_I2[1] ) ) ;
direct_interc direct_interc_34_ (
    .in ( { SYNOPSYS_UNCONNECTED_35 } ) ,
    .out ( clb_I2[2] ) ) ;
direct_interc direct_interc_35_ (
    .in ( { SYNOPSYS_UNCONNECTED_36 } ) ,
    .out ( clb_I2[3] ) ) ;
direct_interc direct_interc_36_ (
    .in ( { SYNOPSYS_UNCONNECTED_37 } ) ,
    .out ( logical_tile_clb_mode_default__fle_1_fle_regout ) ) ;
direct_interc direct_interc_37_ (
    .in ( { SYNOPSYS_UNCONNECTED_38 } ) ,
    .out ( logical_tile_clb_mode_default__fle_1_fle_scout ) ) ;
direct_interc direct_interc_38_ (
    .in ( { SYNOPSYS_UNCONNECTED_39 } ) ,
    .out ( clb_clk ) ) ;
direct_interc direct_interc_39_ (
    .in ( { SYNOPSYS_UNCONNECTED_40 } ) ,
    .out ( clb_I3[0] ) ) ;
direct_interc direct_interc_40_ (
    .in ( { SYNOPSYS_UNCONNECTED_41 } ) ,
    .out ( clb_I3[1] ) ) ;
direct_interc direct_interc_41_ (
    .in ( { SYNOPSYS_UNCONNECTED_42 } ) ,
    .out ( clb_I3[2] ) ) ;
direct_interc direct_interc_42_ (
    .in ( { SYNOPSYS_UNCONNECTED_43 } ) ,
    .out ( clb_I3[3] ) ) ;
direct_interc direct_interc_43_ (
    .in ( { SYNOPSYS_UNCONNECTED_44 } ) ,
    .out ( logical_tile_clb_mode_default__fle_2_fle_regout ) ) ;
direct_interc direct_interc_44_ (
    .in ( { SYNOPSYS_UNCONNECTED_45 } ) ,
    .out ( logical_tile_clb_mode_default__fle_2_fle_scout ) ) ;
direct_interc direct_interc_45_ (
    .in ( { SYNOPSYS_UNCONNECTED_46 } ) ,
    .out ( clb_clk ) ) ;
direct_interc direct_interc_46_ (
    .in ( { SYNOPSYS_UNCONNECTED_47 } ) ,
    .out ( clb_I4[0] ) ) ;
direct_interc direct_interc_47_ (
    .in ( { SYNOPSYS_UNCONNECTED_48 } ) ,
    .out ( clb_I4[1] ) ) ;
direct_interc direct_interc_48_ (
    .in ( { SYNOPSYS_UNCONNECTED_49 } ) ,
    .out ( clb_I4[2] ) ) ;
direct_interc direct_interc_49_ (
    .in ( { SYNOPSYS_UNCONNECTED_50 } ) ,
    .out ( clb_I4[3] ) ) ;
direct_interc direct_interc_50_ (
    .in ( { SYNOPSYS_UNCONNECTED_51 } ) ,
    .out ( logical_tile_clb_mode_default__fle_3_fle_regout ) ) ;
direct_interc direct_interc_51_ (
    .in ( { SYNOPSYS_UNCONNECTED_52 } ) ,
    .out ( logical_tile_clb_mode_default__fle_3_fle_scout ) ) ;
direct_interc direct_interc_52_ (
    .in ( { SYNOPSYS_UNCONNECTED_53 } ) ,
    .out ( clb_clk ) ) ;
direct_interc direct_interc_53_ (
    .in ( { SYNOPSYS_UNCONNECTED_54 } ) ,
    .out ( clb_I5[0] ) ) ;
direct_interc direct_interc_54_ (
    .in ( { SYNOPSYS_UNCONNECTED_55 } ) ,
    .out ( clb_I5[1] ) ) ;
direct_interc direct_interc_55_ (
    .in ( { SYNOPSYS_UNCONNECTED_56 } ) ,
    .out ( clb_I5[2] ) ) ;
direct_interc direct_interc_56_ (
    .in ( { SYNOPSYS_UNCONNECTED_57 } ) ,
    .out ( clb_I5[3] ) ) ;
direct_interc direct_interc_57_ (
    .in ( { SYNOPSYS_UNCONNECTED_58 } ) ,
    .out ( logical_tile_clb_mode_default__fle_4_fle_regout ) ) ;
direct_interc direct_interc_58_ (
    .in ( { SYNOPSYS_UNCONNECTED_59 } ) ,
    .out ( logical_tile_clb_mode_default__fle_4_fle_scout ) ) ;
direct_interc direct_interc_59_ (
    .in ( { SYNOPSYS_UNCONNECTED_60 } ) ,
    .out ( clb_clk ) ) ;
direct_interc direct_interc_60_ (
    .in ( { SYNOPSYS_UNCONNECTED_61 } ) ,
    .out ( clb_I6[0] ) ) ;
direct_interc direct_interc_61_ (
    .in ( { SYNOPSYS_UNCONNECTED_62 } ) ,
    .out ( clb_I6[1] ) ) ;
direct_interc direct_interc_62_ (
    .in ( { SYNOPSYS_UNCONNECTED_63 } ) ,
    .out ( clb_I6[2] ) ) ;
direct_interc direct_interc_63_ (
    .in ( { SYNOPSYS_UNCONNECTED_64 } ) ,
    .out ( clb_I6[3] ) ) ;
direct_interc direct_interc_64_ (
    .in ( { SYNOPSYS_UNCONNECTED_65 } ) ,
    .out ( logical_tile_clb_mode_default__fle_5_fle_regout ) ) ;
direct_interc direct_interc_65_ (
    .in ( { SYNOPSYS_UNCONNECTED_66 } ) ,
    .out ( logical_tile_clb_mode_default__fle_5_fle_scout ) ) ;
direct_interc direct_interc_66_ (
    .in ( { SYNOPSYS_UNCONNECTED_67 } ) ,
    .out ( clb_clk ) ) ;
direct_interc direct_interc_67_ (
    .in ( { SYNOPSYS_UNCONNECTED_68 } ) ,
    .out ( clb_I7[0] ) ) ;
direct_interc direct_interc_68_ (
    .in ( { SYNOPSYS_UNCONNECTED_69 } ) ,
    .out ( clb_I7[1] ) ) ;
direct_interc direct_interc_69_ (
    .in ( { SYNOPSYS_UNCONNECTED_70 } ) ,
    .out ( clb_I7[2] ) ) ;
direct_interc direct_interc_70_ (
    .in ( { SYNOPSYS_UNCONNECTED_71 } ) ,
    .out ( clb_I7[3] ) ) ;
direct_interc direct_interc_71_ (
    .in ( { SYNOPSYS_UNCONNECTED_72 } ) ,
    .out ( logical_tile_clb_mode_default__fle_6_fle_regout ) ) ;
direct_interc direct_interc_72_ (
    .in ( { SYNOPSYS_UNCONNECTED_73 } ) ,
    .out ( logical_tile_clb_mode_default__fle_6_fle_scout ) ) ;
direct_interc direct_interc_73_ (
    .in ( { SYNOPSYS_UNCONNECTED_74 } ) ,
    .out ( clb_clk ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_57 ( 
    .A ( logical_tile_clb_mode_default__fle_0_fle_out[0] ) , .X ( clb_O[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_61 ( 
    .A ( logical_tile_clb_mode_default__fle_1_fle_out[0] ) , .X ( clb_O[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_60 ( .A ( clb_O[0] ) , .X ( p_abuf1 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_62 ( 
    .A ( logical_tile_clb_mode_default__fle_1_fle_out[0] ) , .X ( p_abuf2 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_63 ( .A ( p_abuf3 ) , .X ( clb_O[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_66 ( .A ( p_abuf5 ) , .X ( clb_O[4] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_65 ( .A ( clb_O[5] ) , 
    .X ( BUF_net_65 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_71 ( 
    .A ( logical_tile_clb_mode_default__fle_4_fle_out[0] ) , .X ( clb_O[9] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_68 ( .A ( clb_O[7] ) , 
    .X ( BUF_net_68 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_70 ( .A ( clb_O[6] ) , .X ( p_abuf7 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_72 ( 
    .A ( logical_tile_clb_mode_default__fle_4_fle_out[0] ) , 
    .X ( BUF_net_72 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_73 ( 
    .A ( logical_tile_clb_mode_default__fle_4_fle_out[1] ) , .X ( clb_O[8] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_74 ( 
    .A ( logical_tile_clb_mode_default__fle_4_fle_out[1] ) , 
    .X ( BUF_net_74 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_81 ( 
    .A ( logical_tile_clb_mode_default__fle_6_fle_out[1] ) , 
    .X ( clb_O[12] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_76 ( .A ( clb_O[11] ) , 
    .X ( BUF_net_76 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_78 ( .A ( clb_O[10] ) , 
    .X ( BUF_net_78 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_80 ( .A ( clb_O[13] ) , 
    .X ( BUF_net_80 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_82 ( 
    .A ( logical_tile_clb_mode_default__fle_6_fle_out[1] ) , 
    .X ( BUF_net_82 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_85 ( 
    .A ( logical_tile_clb_mode_default__fle_7_fle_out[1] ) , 
    .X ( clb_O[14] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_84 ( .A ( clb_O[15] ) , 
    .X ( BUF_net_84 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_86 ( 
    .A ( logical_tile_clb_mode_default__fle_7_fle_out[1] ) , 
    .X ( BUF_net_86 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_103 ( .A ( BUF_net_65 ) , 
    .X ( BUF_net_103 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_104 ( .A ( BUF_net_68 ) , 
    .X ( BUF_net_104 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_105 ( .A ( BUF_net_76 ) , 
    .X ( p_abuf10 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_106 ( .A ( BUF_net_82 ) , 
    .X ( p_abuf13 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_107 ( .A ( BUF_net_84 ) , 
    .X ( p_abuf14 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_108 ( .A ( BUF_net_86 ) , 
    .X ( p_abuf15 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_114 ( .A ( BUF_net_72 ) , 
    .X ( p_abuf8 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_115 ( .A ( BUF_net_74 ) , 
    .X ( p_abuf9 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_P_116 ( .A ( BUF_net_78 ) , 
    .X ( p_abuf11 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_P_117 ( .A ( BUF_net_80 ) , 
    .X ( p_abuf12 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_P_123 ( .A ( BUF_net_103 ) , 
    .X ( p_abuf4 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_124 ( .A ( BUF_net_104 ) , 
    .X ( p_abuf6 ) ) ;
endmodule


module grid_clb ( prog_clk , Test_en , clk , top_width_0_height_0__pin_32_ , 
    top_width_0_height_0__pin_33_ , right_width_0_height_0__pin_0_ , 
    right_width_0_height_0__pin_1_ , right_width_0_height_0__pin_2_ , 
    right_width_0_height_0__pin_3_ , right_width_0_height_0__pin_4_ , 
    right_width_0_height_0__pin_5_ , right_width_0_height_0__pin_6_ , 
    right_width_0_height_0__pin_7_ , right_width_0_height_0__pin_8_ , 
    right_width_0_height_0__pin_9_ , right_width_0_height_0__pin_10_ , 
    right_width_0_height_0__pin_11_ , right_width_0_height_0__pin_12_ , 
    right_width_0_height_0__pin_13_ , right_width_0_height_0__pin_14_ , 
    right_width_0_height_0__pin_15_ , bottom_width_0_height_0__pin_16_ , 
    bottom_width_0_height_0__pin_17_ , bottom_width_0_height_0__pin_18_ , 
    bottom_width_0_height_0__pin_19_ , bottom_width_0_height_0__pin_20_ , 
    bottom_width_0_height_0__pin_21_ , bottom_width_0_height_0__pin_22_ , 
    bottom_width_0_height_0__pin_23_ , bottom_width_0_height_0__pin_24_ , 
    bottom_width_0_height_0__pin_25_ , bottom_width_0_height_0__pin_26_ , 
    bottom_width_0_height_0__pin_27_ , bottom_width_0_height_0__pin_28_ , 
    bottom_width_0_height_0__pin_29_ , bottom_width_0_height_0__pin_30_ , 
    bottom_width_0_height_0__pin_31_ , left_width_0_height_0__pin_52_ , 
    ccff_head , right_width_0_height_0__pin_34_upper , 
    right_width_0_height_0__pin_34_lower , 
    right_width_0_height_0__pin_35_upper , 
    right_width_0_height_0__pin_35_lower , 
    right_width_0_height_0__pin_36_upper , 
    right_width_0_height_0__pin_36_lower , 
    right_width_0_height_0__pin_37_upper , 
    right_width_0_height_0__pin_37_lower , 
    right_width_0_height_0__pin_38_upper , 
    right_width_0_height_0__pin_38_lower , 
    right_width_0_height_0__pin_39_upper , 
    right_width_0_height_0__pin_39_lower , 
    right_width_0_height_0__pin_40_upper , 
    right_width_0_height_0__pin_40_lower , 
    right_width_0_height_0__pin_41_upper , 
    right_width_0_height_0__pin_41_lower , 
    bottom_width_0_height_0__pin_42_upper , 
    bottom_width_0_height_0__pin_42_lower , 
    bottom_width_0_height_0__pin_43_upper , 
    bottom_width_0_height_0__pin_43_lower , 
    bottom_width_0_height_0__pin_44_upper , 
    bottom_width_0_height_0__pin_44_lower , 
    bottom_width_0_height_0__pin_45_upper , 
    bottom_width_0_height_0__pin_45_lower , 
    bottom_width_0_height_0__pin_46_upper , 
    bottom_width_0_height_0__pin_46_lower , 
    bottom_width_0_height_0__pin_47_upper , 
    bottom_width_0_height_0__pin_47_lower , 
    bottom_width_0_height_0__pin_48_upper , 
    bottom_width_0_height_0__pin_48_lower , 
    bottom_width_0_height_0__pin_49_upper , 
    bottom_width_0_height_0__pin_49_lower , bottom_width_0_height_0__pin_50_ , 
    bottom_width_0_height_0__pin_51_ , ccff_tail ) ;
input  [0:0] prog_clk ;
input  [0:0] Test_en ;
input  [0:0] clk ;
input  [0:0] top_width_0_height_0__pin_32_ ;
input  [0:0] top_width_0_height_0__pin_33_ ;
input  [0:0] right_width_0_height_0__pin_0_ ;
input  [0:0] right_width_0_height_0__pin_1_ ;
input  [0:0] right_width_0_height_0__pin_2_ ;
input  [0:0] right_width_0_height_0__pin_3_ ;
input  [0:0] right_width_0_height_0__pin_4_ ;
input  [0:0] right_width_0_height_0__pin_5_ ;
input  [0:0] right_width_0_height_0__pin_6_ ;
input  [0:0] right_width_0_height_0__pin_7_ ;
input  [0:0] right_width_0_height_0__pin_8_ ;
input  [0:0] right_width_0_height_0__pin_9_ ;
input  [0:0] right_width_0_height_0__pin_10_ ;
input  [0:0] right_width_0_height_0__pin_11_ ;
input  [0:0] right_width_0_height_0__pin_12_ ;
input  [0:0] right_width_0_height_0__pin_13_ ;
input  [0:0] right_width_0_height_0__pin_14_ ;
input  [0:0] right_width_0_height_0__pin_15_ ;
input  [0:0] bottom_width_0_height_0__pin_16_ ;
input  [0:0] bottom_width_0_height_0__pin_17_ ;
input  [0:0] bottom_width_0_height_0__pin_18_ ;
input  [0:0] bottom_width_0_height_0__pin_19_ ;
input  [0:0] bottom_width_0_height_0__pin_20_ ;
input  [0:0] bottom_width_0_height_0__pin_21_ ;
input  [0:0] bottom_width_0_height_0__pin_22_ ;
input  [0:0] bottom_width_0_height_0__pin_23_ ;
input  [0:0] bottom_width_0_height_0__pin_24_ ;
input  [0:0] bottom_width_0_height_0__pin_25_ ;
input  [0:0] bottom_width_0_height_0__pin_26_ ;
input  [0:0] bottom_width_0_height_0__pin_27_ ;
input  [0:0] bottom_width_0_height_0__pin_28_ ;
input  [0:0] bottom_width_0_height_0__pin_29_ ;
input  [0:0] bottom_width_0_height_0__pin_30_ ;
input  [0:0] bottom_width_0_height_0__pin_31_ ;
input  [0:0] left_width_0_height_0__pin_52_ ;
input  [0:0] ccff_head ;
output [0:0] right_width_0_height_0__pin_34_upper ;
output [0:0] right_width_0_height_0__pin_34_lower ;
output [0:0] right_width_0_height_0__pin_35_upper ;
output [0:0] right_width_0_height_0__pin_35_lower ;
output [0:0] right_width_0_height_0__pin_36_upper ;
output [0:0] right_width_0_height_0__pin_36_lower ;
output [0:0] right_width_0_height_0__pin_37_upper ;
output [0:0] right_width_0_height_0__pin_37_lower ;
output [0:0] right_width_0_height_0__pin_38_upper ;
output [0:0] right_width_0_height_0__pin_38_lower ;
output [0:0] right_width_0_height_0__pin_39_upper ;
output [0:0] right_width_0_height_0__pin_39_lower ;
output [0:0] right_width_0_height_0__pin_40_upper ;
output [0:0] right_width_0_height_0__pin_40_lower ;
output [0:0] right_width_0_height_0__pin_41_upper ;
output [0:0] right_width_0_height_0__pin_41_lower ;
output [0:0] bottom_width_0_height_0__pin_42_upper ;
output [0:0] bottom_width_0_height_0__pin_42_lower ;
output [0:0] bottom_width_0_height_0__pin_43_upper ;
output [0:0] bottom_width_0_height_0__pin_43_lower ;
output [0:0] bottom_width_0_height_0__pin_44_upper ;
output [0:0] bottom_width_0_height_0__pin_44_lower ;
output [0:0] bottom_width_0_height_0__pin_45_upper ;
output [0:0] bottom_width_0_height_0__pin_45_lower ;
output [0:0] bottom_width_0_height_0__pin_46_upper ;
output [0:0] bottom_width_0_height_0__pin_46_lower ;
output [0:0] bottom_width_0_height_0__pin_47_upper ;
output [0:0] bottom_width_0_height_0__pin_47_lower ;
output [0:0] bottom_width_0_height_0__pin_48_upper ;
output [0:0] bottom_width_0_height_0__pin_48_lower ;
output [0:0] bottom_width_0_height_0__pin_49_upper ;
output [0:0] bottom_width_0_height_0__pin_49_lower ;
output [0:0] bottom_width_0_height_0__pin_50_ ;
output [0:0] bottom_width_0_height_0__pin_51_ ;
output [0:0] ccff_tail ;

wire p_abuf3 ;
wire ropt_net_141 ;
wire p_abuf5 ;
wire ropt_net_149 ;
wire ropt_net_154 ;
wire ropt_net_142 ;
wire ropt_net_137 ;
wire ropt_net_138 ;
wire ropt_net_150 ;
wire ropt_net_152 ;
wire ropt_net_140 ;

logical_tile_clb_mode_clb_ logical_tile_clb_mode_clb__0 ( 
    .prog_clk ( prog_clk ) , .Test_en ( Test_en ) , .clk ( clk ) ,
    .clb_I0 ( { right_width_0_height_0__pin_0_[0] , 
        right_width_0_height_0__pin_1_[0] , 
        right_width_0_height_0__pin_2_[0] , 
        right_width_0_height_0__pin_3_[0] } ) ,
    .clb_I1 ( { right_width_0_height_0__pin_4_[0] , 
        right_width_0_height_0__pin_5_[0] , 
        right_width_0_height_0__pin_6_[0] , 
        right_width_0_height_0__pin_7_[0] } ) ,
    .clb_I2 ( { right_width_0_height_0__pin_8_[0] , 
        right_width_0_height_0__pin_9_[0] , 
        right_width_0_height_0__pin_10_[0] , 
        right_width_0_height_0__pin_11_[0] } ) ,
    .clb_I3 ( { right_width_0_height_0__pin_12_[0] , 
        right_width_0_height_0__pin_13_[0] , 
        right_width_0_height_0__pin_14_[0] , 
        right_width_0_height_0__pin_15_[0] } ) ,
    .clb_I4 ( { bottom_width_0_height_0__pin_16_[0] , 
        bottom_width_0_height_0__pin_17_[0] , 
        bottom_width_0_height_0__pin_18_[0] , 
        bottom_width_0_height_0__pin_19_[0] } ) ,
    .clb_I5 ( { bottom_width_0_height_0__pin_20_[0] , 
        bottom_width_0_height_0__pin_21_[0] , 
        bottom_width_0_height_0__pin_22_[0] , 
        bottom_width_0_height_0__pin_23_[0] } ) ,
    .clb_I6 ( { bottom_width_0_height_0__pin_24_[0] , 
        bottom_width_0_height_0__pin_25_[0] , 
        bottom_width_0_height_0__pin_26_[0] , 
        bottom_width_0_height_0__pin_27_[0] } ) ,
    .clb_I7 ( { bottom_width_0_height_0__pin_28_[0] , 
        bottom_width_0_height_0__pin_29_[0] , 
        bottom_width_0_height_0__pin_30_[0] , 
        bottom_width_0_height_0__pin_31_[0] } ) ,
    .clb_regin ( top_width_0_height_0__pin_32_ ) , 
    .clb_scin ( top_width_0_height_0__pin_33_ ) , 
    .clb_clk ( left_width_0_height_0__pin_52_ ) , .ccff_head ( ccff_head ) ,
    .clb_O ( { aps_rename_129_ , ropt_net_132 , ropt_net_139 , 
        aps_rename_133_ , right_width_0_height_0__pin_38_upper[0] , 
        aps_rename_136_ , aps_rename_138_ , aps_rename_140_ , 
        aps_rename_142_ , aps_rename_144_ , aps_rename_146_ , 
        aps_rename_148_ , aps_rename_150_ , aps_rename_151_ , 
        aps_rename_153_ , aps_rename_154_ } ) ,
    .clb_regout ( bottom_width_0_height_0__pin_50_ ) , 
    .clb_scout ( bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( ccff_tail ) , 
    .p_abuf1 ( right_width_0_height_0__pin_34_upper[0] ) , 
    .p_abuf2 ( ropt_net_141 ) , .p_abuf3 ( p_abuf3 ) , 
    .p_abuf4 ( right_width_0_height_0__pin_39_upper[0] ) , 
    .p_abuf5 ( p_abuf5 ) , .p_abuf6 ( ropt_net_154 ) , 
    .p_abuf7 ( ropt_net_149 ) , .p_abuf8 ( ropt_net_137 ) , 
    .p_abuf9 ( ropt_net_142 ) , .p_abuf10 ( ropt_net_138 ) , 
    .p_abuf11 ( bottom_width_0_height_0__pin_44_upper[0] ) , 
    .p_abuf12 ( bottom_width_0_height_0__pin_47_upper[0] ) , 
    .p_abuf13 ( ropt_net_150 ) , .p_abuf14 ( ropt_net_140 ) , 
    .p_abuf15 ( ropt_net_152 ) , .p0 ( optlc_net_126 ) , 
    .p1 ( optlc_net_127 ) , .p2 ( optlc_net_128 ) , .p3 ( optlc_net_129 ) , 
    .p4 ( optlc_net_130 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_1__0 ( .A ( aps_rename_129_ ) , 
    .X ( aps_rename_130_ ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_2__1 ( .A ( ropt_net_132 ) , 
    .X ( aps_rename_131_ ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_3__2 ( .A ( p_abuf3 ) , 
    .X ( aps_rename_132_ ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_4__3 ( .A ( aps_rename_133_ ) , 
    .X ( aps_rename_134_ ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_5__4 ( .A ( p_abuf5 ) , 
    .X ( aps_rename_135_ ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_6__5 ( .A ( aps_rename_136_ ) , 
    .X ( aps_rename_137_ ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_7__6 ( .A ( aps_rename_138_ ) , 
    .X ( aps_rename_139_ ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_8__7 ( .A ( aps_rename_140_ ) , 
    .X ( aps_rename_141_ ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_9__8 ( .A ( aps_rename_142_ ) , 
    .X ( aps_rename_143_ ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_10__9 ( .A ( aps_rename_144_ ) , 
    .X ( aps_rename_145_ ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_11__10 ( .A ( aps_rename_146_ ) , 
    .X ( aps_rename_147_ ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_12__11 ( .A ( aps_rename_148_ ) , 
    .X ( aps_rename_149_ ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_13__12 ( .A ( aps_rename_150_ ) , 
    .X ( ropt_net_134 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_14__13 ( .A ( aps_rename_151_ ) , 
    .X ( aps_rename_152_ ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_15__14 ( .A ( aps_rename_153_ ) , 
    .X ( ropt_net_135 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_16__15 ( .A ( aps_rename_154_ ) , 
    .X ( aps_rename_155_ ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_89 ( .A ( aps_rename_130_ ) , 
    .X ( right_width_0_height_0__pin_34_lower[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_90 ( .A ( aps_rename_131_ ) , 
    .X ( BUF_net_90 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_91 ( .A ( aps_rename_132_ ) , 
    .X ( BUF_net_91 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_92 ( .A ( aps_rename_134_ ) , 
    .X ( BUF_net_92 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_93 ( .A ( aps_rename_135_ ) , 
    .X ( right_width_0_height_0__pin_38_lower[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_94 ( .A ( aps_rename_137_ ) , 
    .X ( right_width_0_height_0__pin_39_lower[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_95 ( .A ( aps_rename_139_ ) , 
    .X ( right_width_0_height_0__pin_40_lower[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_96 ( .A ( aps_rename_141_ ) , 
    .X ( right_width_0_height_0__pin_41_lower[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_97 ( .A ( aps_rename_143_ ) , 
    .X ( ropt_net_133 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_98 ( .A ( aps_rename_145_ ) , 
    .X ( ropt_net_136 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_99 ( .A ( aps_rename_147_ ) , 
    .X ( ropt_net_147 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_100 ( .A ( aps_rename_149_ ) , 
    .X ( BUF_net_100 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_101 ( .A ( aps_rename_152_ ) , 
    .X ( ropt_net_145 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_102 ( .A ( aps_rename_155_ ) , 
    .X ( ropt_net_146 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_119 ( .A ( BUF_net_90 ) , 
    .X ( ropt_net_144 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_120 ( .A ( BUF_net_91 ) , 
    .X ( ropt_net_143 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_P_121 ( .A ( BUF_net_92 ) , 
    .X ( right_width_0_height_0__pin_37_lower[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_P_122 ( .A ( BUF_net_100 ) , 
    .X ( ropt_net_148 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_127 ( .LO ( SYNOPSYS_UNCONNECTED_1 ) , 
    .HI ( optlc_net_126 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_130 ( .LO ( SYNOPSYS_UNCONNECTED_2 ) , 
    .HI ( optlc_net_127 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_132 ( .LO ( SYNOPSYS_UNCONNECTED_3 ) , 
    .HI ( optlc_net_128 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_134 ( .LO ( SYNOPSYS_UNCONNECTED_4 ) , 
    .HI ( optlc_net_129 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_136 ( .LO ( SYNOPSYS_UNCONNECTED_5 ) , 
    .HI ( optlc_net_130 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 ropt_mt_inst_885 ( .A ( ropt_net_132 ) , 
    .X ( right_width_0_height_0__pin_35_upper[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 ropt_mt_inst_886 ( .A ( ropt_net_133 ) , 
    .X ( bottom_width_0_height_0__pin_42_lower[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 ropt_mt_inst_887 ( .A ( ropt_net_134 ) , 
    .X ( bottom_width_0_height_0__pin_46_lower[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 ropt_mt_inst_888 ( .A ( ropt_net_135 ) , 
    .X ( bottom_width_0_height_0__pin_48_lower[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 ropt_mt_inst_891 ( .A ( ropt_net_136 ) , 
    .X ( bottom_width_0_height_0__pin_43_lower[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 ropt_mt_inst_893 ( .A ( ropt_net_137 ) , 
    .X ( bottom_width_0_height_0__pin_43_upper[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 ropt_mt_inst_894 ( .A ( ropt_net_138 ) , 
    .X ( bottom_width_0_height_0__pin_45_upper[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 ropt_mt_inst_895 ( .A ( ropt_net_139 ) , 
    .X ( right_width_0_height_0__pin_36_upper[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 ropt_mt_inst_899 ( .A ( ropt_net_140 ) , 
    .X ( ropt_net_151 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 ropt_mt_inst_900 ( .A ( ropt_net_141 ) , 
    .X ( ropt_net_153 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 ropt_mt_inst_901 ( .A ( ropt_net_142 ) , 
    .X ( bottom_width_0_height_0__pin_42_upper[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 ropt_mt_inst_911 ( .A ( ropt_net_143 ) , 
    .X ( right_width_0_height_0__pin_36_lower[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 ropt_mt_inst_913 ( .A ( ropt_net_144 ) , 
    .X ( right_width_0_height_0__pin_35_lower[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 ropt_mt_inst_914 ( .A ( ropt_net_145 ) , 
    .X ( bottom_width_0_height_0__pin_47_lower[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 ropt_mt_inst_915 ( .A ( ropt_net_146 ) , 
    .X ( bottom_width_0_height_0__pin_49_lower[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 ropt_mt_inst_916 ( .A ( ropt_net_147 ) , 
    .X ( bottom_width_0_height_0__pin_44_lower[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 ropt_mt_inst_917 ( .A ( ropt_net_148 ) , 
    .X ( bottom_width_0_height_0__pin_45_lower[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 ropt_mt_inst_927 ( .A ( ropt_net_149 ) , 
    .X ( right_width_0_height_0__pin_40_upper[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 ropt_mt_inst_928 ( .A ( ropt_net_150 ) , 
    .X ( bottom_width_0_height_0__pin_46_upper[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 ropt_mt_inst_930 ( .A ( ropt_net_151 ) , 
    .X ( bottom_width_0_height_0__pin_49_upper[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 ropt_mt_inst_936 ( .A ( ropt_net_152 ) , 
    .X ( bottom_width_0_height_0__pin_48_upper[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 ropt_mt_inst_938 ( .A ( ropt_net_153 ) , 
    .X ( right_width_0_height_0__pin_37_upper[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 ropt_mt_inst_939 ( .A ( ropt_net_154 ) , 
    .X ( right_width_0_height_0__pin_41_upper[0] ) ) ;
endmodule


module fpga_core ( prog_clk , Test_en , clk , gfpga_pad_GPIO_A , 
    gfpga_pad_GPIO_IE , gfpga_pad_GPIO_OE , gfpga_pad_GPIO_Y , ccff_head , 
    ccff_tail ) ;
input  [0:0] prog_clk ;
input  [0:0] Test_en ;
input  [0:0] clk ;
output [0:47] gfpga_pad_GPIO_A ;
output [0:47] gfpga_pad_GPIO_IE ;
output [0:47] gfpga_pad_GPIO_OE ;
inout  [0:47] gfpga_pad_GPIO_Y ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;

wire [0:0] cbx_1__0__0_bottom_grid_pin_0_ ;
wire [0:0] cbx_1__0__0_ccff_tail ;
wire [0:19] cbx_1__0__0_chanx_left_out ;
wire [0:19] cbx_1__0__0_chanx_right_out ;
wire [0:0] cbx_1__0__0_top_grid_pin_16_ ;
wire [0:0] cbx_1__0__0_top_grid_pin_17_ ;
wire [0:0] cbx_1__0__0_top_grid_pin_18_ ;
wire [0:0] cbx_1__0__0_top_grid_pin_19_ ;
wire [0:0] cbx_1__0__0_top_grid_pin_20_ ;
wire [0:0] cbx_1__0__0_top_grid_pin_21_ ;
wire [0:0] cbx_1__0__0_top_grid_pin_22_ ;
wire [0:0] cbx_1__0__0_top_grid_pin_23_ ;
wire [0:0] cbx_1__0__0_top_grid_pin_24_ ;
wire [0:0] cbx_1__0__0_top_grid_pin_25_ ;
wire [0:0] cbx_1__0__0_top_grid_pin_26_ ;
wire [0:0] cbx_1__0__0_top_grid_pin_27_ ;
wire [0:0] cbx_1__0__0_top_grid_pin_28_ ;
wire [0:0] cbx_1__0__0_top_grid_pin_29_ ;
wire [0:0] cbx_1__0__0_top_grid_pin_30_ ;
wire [0:0] cbx_1__0__0_top_grid_pin_31_ ;
wire [0:0] cbx_1__0__10_bottom_grid_pin_0_ ;
wire [0:0] cbx_1__0__10_ccff_tail ;
wire [0:19] cbx_1__0__10_chanx_left_out ;
wire [0:19] cbx_1__0__10_chanx_right_out ;
wire [0:0] cbx_1__0__10_top_grid_pin_16_ ;
wire [0:0] cbx_1__0__10_top_grid_pin_17_ ;
wire [0:0] cbx_1__0__10_top_grid_pin_18_ ;
wire [0:0] cbx_1__0__10_top_grid_pin_19_ ;
wire [0:0] cbx_1__0__10_top_grid_pin_20_ ;
wire [0:0] cbx_1__0__10_top_grid_pin_21_ ;
wire [0:0] cbx_1__0__10_top_grid_pin_22_ ;
wire [0:0] cbx_1__0__10_top_grid_pin_23_ ;
wire [0:0] cbx_1__0__10_top_grid_pin_24_ ;
wire [0:0] cbx_1__0__10_top_grid_pin_25_ ;
wire [0:0] cbx_1__0__10_top_grid_pin_26_ ;
wire [0:0] cbx_1__0__10_top_grid_pin_27_ ;
wire [0:0] cbx_1__0__10_top_grid_pin_28_ ;
wire [0:0] cbx_1__0__10_top_grid_pin_29_ ;
wire [0:0] cbx_1__0__10_top_grid_pin_30_ ;
wire [0:0] cbx_1__0__10_top_grid_pin_31_ ;
wire [0:0] cbx_1__0__11_bottom_grid_pin_0_ ;
wire [0:0] cbx_1__0__11_ccff_tail ;
wire [0:19] cbx_1__0__11_chanx_left_out ;
wire [0:19] cbx_1__0__11_chanx_right_out ;
wire [0:0] cbx_1__0__11_top_grid_pin_16_ ;
wire [0:0] cbx_1__0__11_top_grid_pin_17_ ;
wire [0:0] cbx_1__0__11_top_grid_pin_18_ ;
wire [0:0] cbx_1__0__11_top_grid_pin_19_ ;
wire [0:0] cbx_1__0__11_top_grid_pin_20_ ;
wire [0:0] cbx_1__0__11_top_grid_pin_21_ ;
wire [0:0] cbx_1__0__11_top_grid_pin_22_ ;
wire [0:0] cbx_1__0__11_top_grid_pin_23_ ;
wire [0:0] cbx_1__0__11_top_grid_pin_24_ ;
wire [0:0] cbx_1__0__11_top_grid_pin_25_ ;
wire [0:0] cbx_1__0__11_top_grid_pin_26_ ;
wire [0:0] cbx_1__0__11_top_grid_pin_27_ ;
wire [0:0] cbx_1__0__11_top_grid_pin_28_ ;
wire [0:0] cbx_1__0__11_top_grid_pin_29_ ;
wire [0:0] cbx_1__0__11_top_grid_pin_30_ ;
wire [0:0] cbx_1__0__11_top_grid_pin_31_ ;
wire [0:0] cbx_1__0__1_bottom_grid_pin_0_ ;
wire [0:0] cbx_1__0__1_ccff_tail ;
wire [0:19] cbx_1__0__1_chanx_left_out ;
wire [0:19] cbx_1__0__1_chanx_right_out ;
wire [0:0] cbx_1__0__1_top_grid_pin_16_ ;
wire [0:0] cbx_1__0__1_top_grid_pin_17_ ;
wire [0:0] cbx_1__0__1_top_grid_pin_18_ ;
wire [0:0] cbx_1__0__1_top_grid_pin_19_ ;
wire [0:0] cbx_1__0__1_top_grid_pin_20_ ;
wire [0:0] cbx_1__0__1_top_grid_pin_21_ ;
wire [0:0] cbx_1__0__1_top_grid_pin_22_ ;
wire [0:0] cbx_1__0__1_top_grid_pin_23_ ;
wire [0:0] cbx_1__0__1_top_grid_pin_24_ ;
wire [0:0] cbx_1__0__1_top_grid_pin_25_ ;
wire [0:0] cbx_1__0__1_top_grid_pin_26_ ;
wire [0:0] cbx_1__0__1_top_grid_pin_27_ ;
wire [0:0] cbx_1__0__1_top_grid_pin_28_ ;
wire [0:0] cbx_1__0__1_top_grid_pin_29_ ;
wire [0:0] cbx_1__0__1_top_grid_pin_30_ ;
wire [0:0] cbx_1__0__1_top_grid_pin_31_ ;
wire [0:0] cbx_1__0__2_bottom_grid_pin_0_ ;
wire [0:0] cbx_1__0__2_ccff_tail ;
wire [0:19] cbx_1__0__2_chanx_left_out ;
wire [0:19] cbx_1__0__2_chanx_right_out ;
wire [0:0] cbx_1__0__2_top_grid_pin_16_ ;
wire [0:0] cbx_1__0__2_top_grid_pin_17_ ;
wire [0:0] cbx_1__0__2_top_grid_pin_18_ ;
wire [0:0] cbx_1__0__2_top_grid_pin_19_ ;
wire [0:0] cbx_1__0__2_top_grid_pin_20_ ;
wire [0:0] cbx_1__0__2_top_grid_pin_21_ ;
wire [0:0] cbx_1__0__2_top_grid_pin_22_ ;
wire [0:0] cbx_1__0__2_top_grid_pin_23_ ;
wire [0:0] cbx_1__0__2_top_grid_pin_24_ ;
wire [0:0] cbx_1__0__2_top_grid_pin_25_ ;
wire [0:0] cbx_1__0__2_top_grid_pin_26_ ;
wire [0:0] cbx_1__0__2_top_grid_pin_27_ ;
wire [0:0] cbx_1__0__2_top_grid_pin_28_ ;
wire [0:0] cbx_1__0__2_top_grid_pin_29_ ;
wire [0:0] cbx_1__0__2_top_grid_pin_30_ ;
wire [0:0] cbx_1__0__2_top_grid_pin_31_ ;
wire [0:0] cbx_1__0__3_bottom_grid_pin_0_ ;
wire [0:0] cbx_1__0__3_ccff_tail ;
wire [0:19] cbx_1__0__3_chanx_left_out ;
wire [0:19] cbx_1__0__3_chanx_right_out ;
wire [0:0] cbx_1__0__3_top_grid_pin_16_ ;
wire [0:0] cbx_1__0__3_top_grid_pin_17_ ;
wire [0:0] cbx_1__0__3_top_grid_pin_18_ ;
wire [0:0] cbx_1__0__3_top_grid_pin_19_ ;
wire [0:0] cbx_1__0__3_top_grid_pin_20_ ;
wire [0:0] cbx_1__0__3_top_grid_pin_21_ ;
wire [0:0] cbx_1__0__3_top_grid_pin_22_ ;
wire [0:0] cbx_1__0__3_top_grid_pin_23_ ;
wire [0:0] cbx_1__0__3_top_grid_pin_24_ ;
wire [0:0] cbx_1__0__3_top_grid_pin_25_ ;
wire [0:0] cbx_1__0__3_top_grid_pin_26_ ;
wire [0:0] cbx_1__0__3_top_grid_pin_27_ ;
wire [0:0] cbx_1__0__3_top_grid_pin_28_ ;
wire [0:0] cbx_1__0__3_top_grid_pin_29_ ;
wire [0:0] cbx_1__0__3_top_grid_pin_30_ ;
wire [0:0] cbx_1__0__3_top_grid_pin_31_ ;
wire [0:0] cbx_1__0__4_bottom_grid_pin_0_ ;
wire [0:0] cbx_1__0__4_ccff_tail ;
wire [0:19] cbx_1__0__4_chanx_left_out ;
wire [0:19] cbx_1__0__4_chanx_right_out ;
wire [0:0] cbx_1__0__4_top_grid_pin_16_ ;
wire [0:0] cbx_1__0__4_top_grid_pin_17_ ;
wire [0:0] cbx_1__0__4_top_grid_pin_18_ ;
wire [0:0] cbx_1__0__4_top_grid_pin_19_ ;
wire [0:0] cbx_1__0__4_top_grid_pin_20_ ;
wire [0:0] cbx_1__0__4_top_grid_pin_21_ ;
wire [0:0] cbx_1__0__4_top_grid_pin_22_ ;
wire [0:0] cbx_1__0__4_top_grid_pin_23_ ;
wire [0:0] cbx_1__0__4_top_grid_pin_24_ ;
wire [0:0] cbx_1__0__4_top_grid_pin_25_ ;
wire [0:0] cbx_1__0__4_top_grid_pin_26_ ;
wire [0:0] cbx_1__0__4_top_grid_pin_27_ ;
wire [0:0] cbx_1__0__4_top_grid_pin_28_ ;
wire [0:0] cbx_1__0__4_top_grid_pin_29_ ;
wire [0:0] cbx_1__0__4_top_grid_pin_30_ ;
wire [0:0] cbx_1__0__4_top_grid_pin_31_ ;
wire [0:0] cbx_1__0__5_bottom_grid_pin_0_ ;
wire [0:0] cbx_1__0__5_ccff_tail ;
wire [0:19] cbx_1__0__5_chanx_left_out ;
wire [0:19] cbx_1__0__5_chanx_right_out ;
wire [0:0] cbx_1__0__5_top_grid_pin_16_ ;
wire [0:0] cbx_1__0__5_top_grid_pin_17_ ;
wire [0:0] cbx_1__0__5_top_grid_pin_18_ ;
wire [0:0] cbx_1__0__5_top_grid_pin_19_ ;
wire [0:0] cbx_1__0__5_top_grid_pin_20_ ;
wire [0:0] cbx_1__0__5_top_grid_pin_21_ ;
wire [0:0] cbx_1__0__5_top_grid_pin_22_ ;
wire [0:0] cbx_1__0__5_top_grid_pin_23_ ;
wire [0:0] cbx_1__0__5_top_grid_pin_24_ ;
wire [0:0] cbx_1__0__5_top_grid_pin_25_ ;
wire [0:0] cbx_1__0__5_top_grid_pin_26_ ;
wire [0:0] cbx_1__0__5_top_grid_pin_27_ ;
wire [0:0] cbx_1__0__5_top_grid_pin_28_ ;
wire [0:0] cbx_1__0__5_top_grid_pin_29_ ;
wire [0:0] cbx_1__0__5_top_grid_pin_30_ ;
wire [0:0] cbx_1__0__5_top_grid_pin_31_ ;
wire [0:0] cbx_1__0__6_bottom_grid_pin_0_ ;
wire [0:0] cbx_1__0__6_ccff_tail ;
wire [0:19] cbx_1__0__6_chanx_left_out ;
wire [0:19] cbx_1__0__6_chanx_right_out ;
wire [0:0] cbx_1__0__6_top_grid_pin_16_ ;
wire [0:0] cbx_1__0__6_top_grid_pin_17_ ;
wire [0:0] cbx_1__0__6_top_grid_pin_18_ ;
wire [0:0] cbx_1__0__6_top_grid_pin_19_ ;
wire [0:0] cbx_1__0__6_top_grid_pin_20_ ;
wire [0:0] cbx_1__0__6_top_grid_pin_21_ ;
wire [0:0] cbx_1__0__6_top_grid_pin_22_ ;
wire [0:0] cbx_1__0__6_top_grid_pin_23_ ;
wire [0:0] cbx_1__0__6_top_grid_pin_24_ ;
wire [0:0] cbx_1__0__6_top_grid_pin_25_ ;
wire [0:0] cbx_1__0__6_top_grid_pin_26_ ;
wire [0:0] cbx_1__0__6_top_grid_pin_27_ ;
wire [0:0] cbx_1__0__6_top_grid_pin_28_ ;
wire [0:0] cbx_1__0__6_top_grid_pin_29_ ;
wire [0:0] cbx_1__0__6_top_grid_pin_30_ ;
wire [0:0] cbx_1__0__6_top_grid_pin_31_ ;
wire [0:0] cbx_1__0__7_bottom_grid_pin_0_ ;
wire [0:0] cbx_1__0__7_ccff_tail ;
wire [0:19] cbx_1__0__7_chanx_left_out ;
wire [0:19] cbx_1__0__7_chanx_right_out ;
wire [0:0] cbx_1__0__7_top_grid_pin_16_ ;
wire [0:0] cbx_1__0__7_top_grid_pin_17_ ;
wire [0:0] cbx_1__0__7_top_grid_pin_18_ ;
wire [0:0] cbx_1__0__7_top_grid_pin_19_ ;
wire [0:0] cbx_1__0__7_top_grid_pin_20_ ;
wire [0:0] cbx_1__0__7_top_grid_pin_21_ ;
wire [0:0] cbx_1__0__7_top_grid_pin_22_ ;
wire [0:0] cbx_1__0__7_top_grid_pin_23_ ;
wire [0:0] cbx_1__0__7_top_grid_pin_24_ ;
wire [0:0] cbx_1__0__7_top_grid_pin_25_ ;
wire [0:0] cbx_1__0__7_top_grid_pin_26_ ;
wire [0:0] cbx_1__0__7_top_grid_pin_27_ ;
wire [0:0] cbx_1__0__7_top_grid_pin_28_ ;
wire [0:0] cbx_1__0__7_top_grid_pin_29_ ;
wire [0:0] cbx_1__0__7_top_grid_pin_30_ ;
wire [0:0] cbx_1__0__7_top_grid_pin_31_ ;
wire [0:0] cbx_1__0__8_bottom_grid_pin_0_ ;
wire [0:0] cbx_1__0__8_ccff_tail ;
wire [0:19] cbx_1__0__8_chanx_left_out ;
wire [0:19] cbx_1__0__8_chanx_right_out ;
wire [0:0] cbx_1__0__8_top_grid_pin_16_ ;
wire [0:0] cbx_1__0__8_top_grid_pin_17_ ;
wire [0:0] cbx_1__0__8_top_grid_pin_18_ ;
wire [0:0] cbx_1__0__8_top_grid_pin_19_ ;
wire [0:0] cbx_1__0__8_top_grid_pin_20_ ;
wire [0:0] cbx_1__0__8_top_grid_pin_21_ ;
wire [0:0] cbx_1__0__8_top_grid_pin_22_ ;
wire [0:0] cbx_1__0__8_top_grid_pin_23_ ;
wire [0:0] cbx_1__0__8_top_grid_pin_24_ ;
wire [0:0] cbx_1__0__8_top_grid_pin_25_ ;
wire [0:0] cbx_1__0__8_top_grid_pin_26_ ;
wire [0:0] cbx_1__0__8_top_grid_pin_27_ ;
wire [0:0] cbx_1__0__8_top_grid_pin_28_ ;
wire [0:0] cbx_1__0__8_top_grid_pin_29_ ;
wire [0:0] cbx_1__0__8_top_grid_pin_30_ ;
wire [0:0] cbx_1__0__8_top_grid_pin_31_ ;
wire [0:0] cbx_1__0__9_bottom_grid_pin_0_ ;
wire [0:0] cbx_1__0__9_ccff_tail ;
wire [0:19] cbx_1__0__9_chanx_left_out ;
wire [0:19] cbx_1__0__9_chanx_right_out ;
wire [0:0] cbx_1__0__9_top_grid_pin_16_ ;
wire [0:0] cbx_1__0__9_top_grid_pin_17_ ;
wire [0:0] cbx_1__0__9_top_grid_pin_18_ ;
wire [0:0] cbx_1__0__9_top_grid_pin_19_ ;
wire [0:0] cbx_1__0__9_top_grid_pin_20_ ;
wire [0:0] cbx_1__0__9_top_grid_pin_21_ ;
wire [0:0] cbx_1__0__9_top_grid_pin_22_ ;
wire [0:0] cbx_1__0__9_top_grid_pin_23_ ;
wire [0:0] cbx_1__0__9_top_grid_pin_24_ ;
wire [0:0] cbx_1__0__9_top_grid_pin_25_ ;
wire [0:0] cbx_1__0__9_top_grid_pin_26_ ;
wire [0:0] cbx_1__0__9_top_grid_pin_27_ ;
wire [0:0] cbx_1__0__9_top_grid_pin_28_ ;
wire [0:0] cbx_1__0__9_top_grid_pin_29_ ;
wire [0:0] cbx_1__0__9_top_grid_pin_30_ ;
wire [0:0] cbx_1__0__9_top_grid_pin_31_ ;
wire [0:0] cbx_1__12__0_ccff_tail ;
wire [0:19] cbx_1__12__0_chanx_left_out ;
wire [0:19] cbx_1__12__0_chanx_right_out ;
wire [0:0] cbx_1__12__0_top_grid_pin_0_ ;
wire [0:0] cbx_1__12__10_ccff_tail ;
wire [0:19] cbx_1__12__10_chanx_left_out ;
wire [0:19] cbx_1__12__10_chanx_right_out ;
wire [0:0] cbx_1__12__10_top_grid_pin_0_ ;
wire [0:0] cbx_1__12__11_ccff_tail ;
wire [0:19] cbx_1__12__11_chanx_left_out ;
wire [0:19] cbx_1__12__11_chanx_right_out ;
wire [0:0] cbx_1__12__11_top_grid_pin_0_ ;
wire [0:0] cbx_1__12__1_ccff_tail ;
wire [0:19] cbx_1__12__1_chanx_left_out ;
wire [0:19] cbx_1__12__1_chanx_right_out ;
wire [0:0] cbx_1__12__1_top_grid_pin_0_ ;
wire [0:0] cbx_1__12__2_ccff_tail ;
wire [0:19] cbx_1__12__2_chanx_left_out ;
wire [0:19] cbx_1__12__2_chanx_right_out ;
wire [0:0] cbx_1__12__2_top_grid_pin_0_ ;
wire [0:0] cbx_1__12__3_ccff_tail ;
wire [0:19] cbx_1__12__3_chanx_left_out ;
wire [0:19] cbx_1__12__3_chanx_right_out ;
wire [0:0] cbx_1__12__3_top_grid_pin_0_ ;
wire [0:0] cbx_1__12__4_ccff_tail ;
wire [0:19] cbx_1__12__4_chanx_left_out ;
wire [0:19] cbx_1__12__4_chanx_right_out ;
wire [0:0] cbx_1__12__4_top_grid_pin_0_ ;
wire [0:0] cbx_1__12__5_ccff_tail ;
wire [0:19] cbx_1__12__5_chanx_left_out ;
wire [0:19] cbx_1__12__5_chanx_right_out ;
wire [0:0] cbx_1__12__5_top_grid_pin_0_ ;
wire [0:0] cbx_1__12__6_ccff_tail ;
wire [0:19] cbx_1__12__6_chanx_left_out ;
wire [0:19] cbx_1__12__6_chanx_right_out ;
wire [0:0] cbx_1__12__6_top_grid_pin_0_ ;
wire [0:0] cbx_1__12__7_ccff_tail ;
wire [0:19] cbx_1__12__7_chanx_left_out ;
wire [0:19] cbx_1__12__7_chanx_right_out ;
wire [0:0] cbx_1__12__7_top_grid_pin_0_ ;
wire [0:0] cbx_1__12__8_ccff_tail ;
wire [0:19] cbx_1__12__8_chanx_left_out ;
wire [0:19] cbx_1__12__8_chanx_right_out ;
wire [0:0] cbx_1__12__8_top_grid_pin_0_ ;
wire [0:0] cbx_1__12__9_ccff_tail ;
wire [0:19] cbx_1__12__9_chanx_left_out ;
wire [0:19] cbx_1__12__9_chanx_right_out ;
wire [0:0] cbx_1__12__9_top_grid_pin_0_ ;
wire [0:0] cbx_1__1__0_ccff_tail ;
wire [0:19] cbx_1__1__0_chanx_left_out ;
wire [0:19] cbx_1__1__0_chanx_right_out ;
wire [0:0] cbx_1__1__0_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__0_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__0_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__0_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__0_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__0_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__0_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__0_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__0_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__0_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__0_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__0_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__0_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__0_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__0_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__0_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__100_ccff_tail ;
wire [0:19] cbx_1__1__100_chanx_left_out ;
wire [0:19] cbx_1__1__100_chanx_right_out ;
wire [0:0] cbx_1__1__100_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__100_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__100_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__100_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__100_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__100_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__100_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__100_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__100_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__100_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__100_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__100_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__100_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__100_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__100_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__100_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__101_ccff_tail ;
wire [0:19] cbx_1__1__101_chanx_left_out ;
wire [0:19] cbx_1__1__101_chanx_right_out ;
wire [0:0] cbx_1__1__101_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__101_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__101_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__101_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__101_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__101_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__101_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__101_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__101_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__101_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__101_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__101_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__101_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__101_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__101_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__101_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__102_ccff_tail ;
wire [0:19] cbx_1__1__102_chanx_left_out ;
wire [0:19] cbx_1__1__102_chanx_right_out ;
wire [0:0] cbx_1__1__102_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__102_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__102_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__102_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__102_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__102_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__102_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__102_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__102_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__102_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__102_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__102_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__102_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__102_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__102_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__102_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__103_ccff_tail ;
wire [0:19] cbx_1__1__103_chanx_left_out ;
wire [0:19] cbx_1__1__103_chanx_right_out ;
wire [0:0] cbx_1__1__103_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__103_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__103_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__103_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__103_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__103_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__103_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__103_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__103_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__103_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__103_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__103_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__103_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__103_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__103_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__103_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__104_ccff_tail ;
wire [0:19] cbx_1__1__104_chanx_left_out ;
wire [0:19] cbx_1__1__104_chanx_right_out ;
wire [0:0] cbx_1__1__104_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__104_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__104_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__104_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__104_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__104_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__104_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__104_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__104_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__104_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__104_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__104_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__104_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__104_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__104_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__104_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__105_ccff_tail ;
wire [0:19] cbx_1__1__105_chanx_left_out ;
wire [0:19] cbx_1__1__105_chanx_right_out ;
wire [0:0] cbx_1__1__105_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__105_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__105_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__105_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__105_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__105_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__105_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__105_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__105_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__105_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__105_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__105_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__105_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__105_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__105_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__105_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__106_ccff_tail ;
wire [0:19] cbx_1__1__106_chanx_left_out ;
wire [0:19] cbx_1__1__106_chanx_right_out ;
wire [0:0] cbx_1__1__106_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__106_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__106_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__106_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__106_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__106_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__106_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__106_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__106_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__106_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__106_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__106_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__106_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__106_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__106_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__106_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__107_ccff_tail ;
wire [0:19] cbx_1__1__107_chanx_left_out ;
wire [0:19] cbx_1__1__107_chanx_right_out ;
wire [0:0] cbx_1__1__107_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__107_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__107_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__107_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__107_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__107_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__107_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__107_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__107_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__107_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__107_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__107_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__107_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__107_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__107_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__107_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__108_ccff_tail ;
wire [0:19] cbx_1__1__108_chanx_left_out ;
wire [0:19] cbx_1__1__108_chanx_right_out ;
wire [0:0] cbx_1__1__108_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__108_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__108_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__108_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__108_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__108_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__108_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__108_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__108_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__108_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__108_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__108_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__108_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__108_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__108_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__108_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__109_ccff_tail ;
wire [0:19] cbx_1__1__109_chanx_left_out ;
wire [0:19] cbx_1__1__109_chanx_right_out ;
wire [0:0] cbx_1__1__109_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__109_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__109_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__109_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__109_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__109_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__109_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__109_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__109_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__109_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__109_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__109_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__109_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__109_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__109_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__109_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__10_ccff_tail ;
wire [0:19] cbx_1__1__10_chanx_left_out ;
wire [0:19] cbx_1__1__10_chanx_right_out ;
wire [0:0] cbx_1__1__10_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__10_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__10_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__10_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__10_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__10_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__10_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__10_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__10_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__10_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__10_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__10_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__10_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__10_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__10_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__10_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__110_ccff_tail ;
wire [0:19] cbx_1__1__110_chanx_left_out ;
wire [0:19] cbx_1__1__110_chanx_right_out ;
wire [0:0] cbx_1__1__110_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__110_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__110_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__110_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__110_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__110_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__110_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__110_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__110_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__110_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__110_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__110_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__110_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__110_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__110_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__110_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__111_ccff_tail ;
wire [0:19] cbx_1__1__111_chanx_left_out ;
wire [0:19] cbx_1__1__111_chanx_right_out ;
wire [0:0] cbx_1__1__111_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__111_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__111_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__111_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__111_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__111_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__111_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__111_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__111_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__111_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__111_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__111_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__111_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__111_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__111_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__111_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__112_ccff_tail ;
wire [0:19] cbx_1__1__112_chanx_left_out ;
wire [0:19] cbx_1__1__112_chanx_right_out ;
wire [0:0] cbx_1__1__112_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__112_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__112_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__112_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__112_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__112_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__112_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__112_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__112_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__112_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__112_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__112_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__112_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__112_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__112_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__112_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__113_ccff_tail ;
wire [0:19] cbx_1__1__113_chanx_left_out ;
wire [0:19] cbx_1__1__113_chanx_right_out ;
wire [0:0] cbx_1__1__113_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__113_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__113_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__113_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__113_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__113_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__113_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__113_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__113_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__113_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__113_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__113_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__113_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__113_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__113_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__113_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__114_ccff_tail ;
wire [0:19] cbx_1__1__114_chanx_left_out ;
wire [0:19] cbx_1__1__114_chanx_right_out ;
wire [0:0] cbx_1__1__114_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__114_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__114_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__114_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__114_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__114_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__114_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__114_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__114_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__114_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__114_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__114_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__114_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__114_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__114_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__114_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__115_ccff_tail ;
wire [0:19] cbx_1__1__115_chanx_left_out ;
wire [0:19] cbx_1__1__115_chanx_right_out ;
wire [0:0] cbx_1__1__115_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__115_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__115_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__115_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__115_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__115_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__115_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__115_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__115_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__115_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__115_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__115_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__115_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__115_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__115_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__115_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__116_ccff_tail ;
wire [0:19] cbx_1__1__116_chanx_left_out ;
wire [0:19] cbx_1__1__116_chanx_right_out ;
wire [0:0] cbx_1__1__116_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__116_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__116_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__116_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__116_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__116_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__116_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__116_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__116_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__116_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__116_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__116_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__116_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__116_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__116_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__116_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__117_ccff_tail ;
wire [0:19] cbx_1__1__117_chanx_left_out ;
wire [0:19] cbx_1__1__117_chanx_right_out ;
wire [0:0] cbx_1__1__117_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__117_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__117_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__117_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__117_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__117_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__117_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__117_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__117_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__117_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__117_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__117_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__117_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__117_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__117_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__117_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__118_ccff_tail ;
wire [0:19] cbx_1__1__118_chanx_left_out ;
wire [0:19] cbx_1__1__118_chanx_right_out ;
wire [0:0] cbx_1__1__118_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__118_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__118_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__118_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__118_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__118_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__118_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__118_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__118_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__118_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__118_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__118_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__118_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__118_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__118_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__118_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__119_ccff_tail ;
wire [0:19] cbx_1__1__119_chanx_left_out ;
wire [0:19] cbx_1__1__119_chanx_right_out ;
wire [0:0] cbx_1__1__119_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__119_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__119_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__119_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__119_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__119_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__119_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__119_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__119_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__119_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__119_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__119_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__119_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__119_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__119_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__119_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__11_ccff_tail ;
wire [0:19] cbx_1__1__11_chanx_left_out ;
wire [0:19] cbx_1__1__11_chanx_right_out ;
wire [0:0] cbx_1__1__11_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__11_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__11_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__11_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__11_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__11_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__11_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__11_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__11_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__11_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__11_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__11_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__11_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__11_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__11_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__11_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__120_ccff_tail ;
wire [0:19] cbx_1__1__120_chanx_left_out ;
wire [0:19] cbx_1__1__120_chanx_right_out ;
wire [0:0] cbx_1__1__120_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__120_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__120_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__120_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__120_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__120_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__120_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__120_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__120_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__120_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__120_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__120_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__120_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__120_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__120_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__120_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__121_ccff_tail ;
wire [0:19] cbx_1__1__121_chanx_left_out ;
wire [0:19] cbx_1__1__121_chanx_right_out ;
wire [0:0] cbx_1__1__121_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__121_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__121_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__121_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__121_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__121_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__121_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__121_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__121_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__121_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__121_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__121_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__121_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__121_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__121_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__121_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__122_ccff_tail ;
wire [0:19] cbx_1__1__122_chanx_left_out ;
wire [0:19] cbx_1__1__122_chanx_right_out ;
wire [0:0] cbx_1__1__122_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__122_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__122_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__122_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__122_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__122_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__122_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__122_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__122_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__122_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__122_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__122_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__122_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__122_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__122_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__122_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__123_ccff_tail ;
wire [0:19] cbx_1__1__123_chanx_left_out ;
wire [0:19] cbx_1__1__123_chanx_right_out ;
wire [0:0] cbx_1__1__123_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__123_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__123_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__123_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__123_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__123_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__123_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__123_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__123_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__123_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__123_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__123_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__123_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__123_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__123_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__123_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__124_ccff_tail ;
wire [0:19] cbx_1__1__124_chanx_left_out ;
wire [0:19] cbx_1__1__124_chanx_right_out ;
wire [0:0] cbx_1__1__124_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__124_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__124_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__124_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__124_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__124_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__124_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__124_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__124_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__124_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__124_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__124_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__124_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__124_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__124_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__124_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__125_ccff_tail ;
wire [0:19] cbx_1__1__125_chanx_left_out ;
wire [0:19] cbx_1__1__125_chanx_right_out ;
wire [0:0] cbx_1__1__125_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__125_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__125_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__125_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__125_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__125_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__125_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__125_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__125_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__125_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__125_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__125_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__125_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__125_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__125_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__125_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__126_ccff_tail ;
wire [0:19] cbx_1__1__126_chanx_left_out ;
wire [0:19] cbx_1__1__126_chanx_right_out ;
wire [0:0] cbx_1__1__126_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__126_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__126_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__126_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__126_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__126_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__126_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__126_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__126_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__126_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__126_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__126_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__126_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__126_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__126_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__126_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__127_ccff_tail ;
wire [0:19] cbx_1__1__127_chanx_left_out ;
wire [0:19] cbx_1__1__127_chanx_right_out ;
wire [0:0] cbx_1__1__127_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__127_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__127_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__127_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__127_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__127_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__127_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__127_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__127_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__127_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__127_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__127_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__127_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__127_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__127_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__127_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__128_ccff_tail ;
wire [0:19] cbx_1__1__128_chanx_left_out ;
wire [0:19] cbx_1__1__128_chanx_right_out ;
wire [0:0] cbx_1__1__128_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__128_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__128_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__128_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__128_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__128_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__128_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__128_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__128_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__128_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__128_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__128_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__128_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__128_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__128_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__128_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__129_ccff_tail ;
wire [0:19] cbx_1__1__129_chanx_left_out ;
wire [0:19] cbx_1__1__129_chanx_right_out ;
wire [0:0] cbx_1__1__129_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__129_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__129_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__129_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__129_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__129_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__129_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__129_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__129_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__129_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__129_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__129_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__129_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__129_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__129_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__129_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__12_ccff_tail ;
wire [0:19] cbx_1__1__12_chanx_left_out ;
wire [0:19] cbx_1__1__12_chanx_right_out ;
wire [0:0] cbx_1__1__12_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__12_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__12_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__12_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__12_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__12_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__12_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__12_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__12_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__12_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__12_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__12_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__12_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__12_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__12_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__12_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__130_ccff_tail ;
wire [0:19] cbx_1__1__130_chanx_left_out ;
wire [0:19] cbx_1__1__130_chanx_right_out ;
wire [0:0] cbx_1__1__130_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__130_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__130_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__130_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__130_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__130_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__130_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__130_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__130_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__130_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__130_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__130_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__130_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__130_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__130_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__130_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__131_ccff_tail ;
wire [0:19] cbx_1__1__131_chanx_left_out ;
wire [0:19] cbx_1__1__131_chanx_right_out ;
wire [0:0] cbx_1__1__131_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__131_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__131_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__131_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__131_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__131_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__131_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__131_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__131_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__131_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__131_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__131_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__131_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__131_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__131_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__131_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__13_ccff_tail ;
wire [0:19] cbx_1__1__13_chanx_left_out ;
wire [0:19] cbx_1__1__13_chanx_right_out ;
wire [0:0] cbx_1__1__13_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__13_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__13_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__13_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__13_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__13_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__13_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__13_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__13_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__13_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__13_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__13_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__13_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__13_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__13_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__13_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__14_ccff_tail ;
wire [0:19] cbx_1__1__14_chanx_left_out ;
wire [0:19] cbx_1__1__14_chanx_right_out ;
wire [0:0] cbx_1__1__14_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__14_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__14_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__14_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__14_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__14_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__14_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__14_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__14_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__14_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__14_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__14_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__14_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__14_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__14_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__14_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__15_ccff_tail ;
wire [0:19] cbx_1__1__15_chanx_left_out ;
wire [0:19] cbx_1__1__15_chanx_right_out ;
wire [0:0] cbx_1__1__15_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__15_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__15_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__15_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__15_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__15_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__15_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__15_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__15_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__15_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__15_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__15_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__15_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__15_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__15_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__15_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__16_ccff_tail ;
wire [0:19] cbx_1__1__16_chanx_left_out ;
wire [0:19] cbx_1__1__16_chanx_right_out ;
wire [0:0] cbx_1__1__16_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__16_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__16_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__16_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__16_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__16_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__16_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__16_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__16_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__16_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__16_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__16_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__16_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__16_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__16_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__16_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__17_ccff_tail ;
wire [0:19] cbx_1__1__17_chanx_left_out ;
wire [0:19] cbx_1__1__17_chanx_right_out ;
wire [0:0] cbx_1__1__17_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__17_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__17_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__17_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__17_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__17_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__17_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__17_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__17_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__17_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__17_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__17_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__17_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__17_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__17_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__17_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__18_ccff_tail ;
wire [0:19] cbx_1__1__18_chanx_left_out ;
wire [0:19] cbx_1__1__18_chanx_right_out ;
wire [0:0] cbx_1__1__18_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__18_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__18_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__18_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__18_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__18_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__18_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__18_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__18_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__18_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__18_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__18_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__18_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__18_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__18_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__18_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__19_ccff_tail ;
wire [0:19] cbx_1__1__19_chanx_left_out ;
wire [0:19] cbx_1__1__19_chanx_right_out ;
wire [0:0] cbx_1__1__19_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__19_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__19_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__19_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__19_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__19_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__19_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__19_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__19_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__19_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__19_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__19_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__19_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__19_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__19_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__19_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__1_ccff_tail ;
wire [0:19] cbx_1__1__1_chanx_left_out ;
wire [0:19] cbx_1__1__1_chanx_right_out ;
wire [0:0] cbx_1__1__1_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__1_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__1_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__1_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__1_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__1_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__1_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__1_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__1_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__1_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__1_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__1_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__1_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__1_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__1_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__1_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__20_ccff_tail ;
wire [0:19] cbx_1__1__20_chanx_left_out ;
wire [0:19] cbx_1__1__20_chanx_right_out ;
wire [0:0] cbx_1__1__20_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__20_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__20_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__20_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__20_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__20_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__20_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__20_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__20_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__20_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__20_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__20_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__20_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__20_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__20_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__20_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__21_ccff_tail ;
wire [0:19] cbx_1__1__21_chanx_left_out ;
wire [0:19] cbx_1__1__21_chanx_right_out ;
wire [0:0] cbx_1__1__21_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__21_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__21_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__21_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__21_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__21_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__21_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__21_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__21_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__21_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__21_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__21_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__21_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__21_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__21_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__21_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__22_ccff_tail ;
wire [0:19] cbx_1__1__22_chanx_left_out ;
wire [0:19] cbx_1__1__22_chanx_right_out ;
wire [0:0] cbx_1__1__22_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__22_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__22_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__22_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__22_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__22_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__22_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__22_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__22_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__22_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__22_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__22_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__22_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__22_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__22_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__22_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__23_ccff_tail ;
wire [0:19] cbx_1__1__23_chanx_left_out ;
wire [0:19] cbx_1__1__23_chanx_right_out ;
wire [0:0] cbx_1__1__23_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__23_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__23_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__23_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__23_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__23_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__23_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__23_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__23_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__23_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__23_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__23_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__23_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__23_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__23_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__23_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__24_ccff_tail ;
wire [0:19] cbx_1__1__24_chanx_left_out ;
wire [0:19] cbx_1__1__24_chanx_right_out ;
wire [0:0] cbx_1__1__24_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__24_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__24_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__24_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__24_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__24_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__24_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__24_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__24_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__24_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__24_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__24_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__24_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__24_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__24_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__24_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__25_ccff_tail ;
wire [0:19] cbx_1__1__25_chanx_left_out ;
wire [0:19] cbx_1__1__25_chanx_right_out ;
wire [0:0] cbx_1__1__25_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__25_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__25_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__25_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__25_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__25_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__25_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__25_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__25_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__25_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__25_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__25_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__25_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__25_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__25_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__25_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__26_ccff_tail ;
wire [0:19] cbx_1__1__26_chanx_left_out ;
wire [0:19] cbx_1__1__26_chanx_right_out ;
wire [0:0] cbx_1__1__26_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__26_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__26_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__26_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__26_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__26_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__26_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__26_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__26_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__26_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__26_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__26_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__26_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__26_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__26_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__26_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__27_ccff_tail ;
wire [0:19] cbx_1__1__27_chanx_left_out ;
wire [0:19] cbx_1__1__27_chanx_right_out ;
wire [0:0] cbx_1__1__27_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__27_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__27_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__27_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__27_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__27_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__27_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__27_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__27_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__27_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__27_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__27_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__27_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__27_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__27_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__27_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__28_ccff_tail ;
wire [0:19] cbx_1__1__28_chanx_left_out ;
wire [0:19] cbx_1__1__28_chanx_right_out ;
wire [0:0] cbx_1__1__28_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__28_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__28_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__28_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__28_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__28_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__28_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__28_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__28_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__28_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__28_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__28_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__28_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__28_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__28_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__28_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__29_ccff_tail ;
wire [0:19] cbx_1__1__29_chanx_left_out ;
wire [0:19] cbx_1__1__29_chanx_right_out ;
wire [0:0] cbx_1__1__29_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__29_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__29_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__29_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__29_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__29_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__29_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__29_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__29_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__29_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__29_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__29_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__29_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__29_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__29_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__29_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__2_ccff_tail ;
wire [0:19] cbx_1__1__2_chanx_left_out ;
wire [0:19] cbx_1__1__2_chanx_right_out ;
wire [0:0] cbx_1__1__2_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__2_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__2_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__2_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__2_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__2_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__2_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__2_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__2_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__2_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__2_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__2_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__2_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__2_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__2_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__2_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__30_ccff_tail ;
wire [0:19] cbx_1__1__30_chanx_left_out ;
wire [0:19] cbx_1__1__30_chanx_right_out ;
wire [0:0] cbx_1__1__30_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__30_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__30_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__30_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__30_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__30_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__30_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__30_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__30_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__30_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__30_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__30_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__30_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__30_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__30_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__30_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__31_ccff_tail ;
wire [0:19] cbx_1__1__31_chanx_left_out ;
wire [0:19] cbx_1__1__31_chanx_right_out ;
wire [0:0] cbx_1__1__31_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__31_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__31_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__31_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__31_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__31_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__31_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__31_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__31_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__31_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__31_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__31_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__31_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__31_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__31_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__31_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__32_ccff_tail ;
wire [0:19] cbx_1__1__32_chanx_left_out ;
wire [0:19] cbx_1__1__32_chanx_right_out ;
wire [0:0] cbx_1__1__32_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__32_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__32_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__32_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__32_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__32_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__32_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__32_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__32_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__32_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__32_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__32_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__32_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__32_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__32_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__32_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__33_ccff_tail ;
wire [0:19] cbx_1__1__33_chanx_left_out ;
wire [0:19] cbx_1__1__33_chanx_right_out ;
wire [0:0] cbx_1__1__33_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__33_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__33_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__33_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__33_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__33_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__33_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__33_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__33_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__33_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__33_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__33_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__33_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__33_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__33_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__33_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__34_ccff_tail ;
wire [0:19] cbx_1__1__34_chanx_left_out ;
wire [0:19] cbx_1__1__34_chanx_right_out ;
wire [0:0] cbx_1__1__34_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__34_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__34_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__34_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__34_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__34_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__34_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__34_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__34_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__34_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__34_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__34_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__34_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__34_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__34_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__34_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__35_ccff_tail ;
wire [0:19] cbx_1__1__35_chanx_left_out ;
wire [0:19] cbx_1__1__35_chanx_right_out ;
wire [0:0] cbx_1__1__35_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__35_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__35_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__35_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__35_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__35_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__35_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__35_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__35_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__35_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__35_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__35_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__35_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__35_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__35_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__35_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__36_ccff_tail ;
wire [0:19] cbx_1__1__36_chanx_left_out ;
wire [0:19] cbx_1__1__36_chanx_right_out ;
wire [0:0] cbx_1__1__36_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__36_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__36_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__36_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__36_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__36_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__36_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__36_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__36_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__36_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__36_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__36_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__36_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__36_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__36_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__36_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__37_ccff_tail ;
wire [0:19] cbx_1__1__37_chanx_left_out ;
wire [0:19] cbx_1__1__37_chanx_right_out ;
wire [0:0] cbx_1__1__37_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__37_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__37_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__37_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__37_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__37_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__37_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__37_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__37_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__37_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__37_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__37_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__37_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__37_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__37_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__37_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__38_ccff_tail ;
wire [0:19] cbx_1__1__38_chanx_left_out ;
wire [0:19] cbx_1__1__38_chanx_right_out ;
wire [0:0] cbx_1__1__38_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__38_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__38_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__38_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__38_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__38_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__38_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__38_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__38_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__38_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__38_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__38_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__38_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__38_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__38_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__38_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__39_ccff_tail ;
wire [0:19] cbx_1__1__39_chanx_left_out ;
wire [0:19] cbx_1__1__39_chanx_right_out ;
wire [0:0] cbx_1__1__39_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__39_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__39_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__39_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__39_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__39_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__39_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__39_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__39_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__39_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__39_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__39_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__39_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__39_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__39_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__39_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__3_ccff_tail ;
wire [0:19] cbx_1__1__3_chanx_left_out ;
wire [0:19] cbx_1__1__3_chanx_right_out ;
wire [0:0] cbx_1__1__3_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__3_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__3_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__3_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__3_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__3_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__3_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__3_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__3_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__3_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__3_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__3_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__3_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__3_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__3_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__3_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__40_ccff_tail ;
wire [0:19] cbx_1__1__40_chanx_left_out ;
wire [0:19] cbx_1__1__40_chanx_right_out ;
wire [0:0] cbx_1__1__40_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__40_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__40_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__40_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__40_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__40_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__40_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__40_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__40_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__40_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__40_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__40_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__40_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__40_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__40_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__40_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__41_ccff_tail ;
wire [0:19] cbx_1__1__41_chanx_left_out ;
wire [0:19] cbx_1__1__41_chanx_right_out ;
wire [0:0] cbx_1__1__41_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__41_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__41_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__41_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__41_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__41_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__41_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__41_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__41_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__41_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__41_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__41_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__41_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__41_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__41_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__41_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__42_ccff_tail ;
wire [0:19] cbx_1__1__42_chanx_left_out ;
wire [0:19] cbx_1__1__42_chanx_right_out ;
wire [0:0] cbx_1__1__42_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__42_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__42_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__42_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__42_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__42_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__42_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__42_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__42_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__42_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__42_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__42_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__42_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__42_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__42_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__42_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__43_ccff_tail ;
wire [0:19] cbx_1__1__43_chanx_left_out ;
wire [0:19] cbx_1__1__43_chanx_right_out ;
wire [0:0] cbx_1__1__43_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__43_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__43_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__43_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__43_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__43_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__43_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__43_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__43_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__43_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__43_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__43_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__43_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__43_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__43_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__43_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__44_ccff_tail ;
wire [0:19] cbx_1__1__44_chanx_left_out ;
wire [0:19] cbx_1__1__44_chanx_right_out ;
wire [0:0] cbx_1__1__44_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__44_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__44_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__44_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__44_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__44_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__44_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__44_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__44_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__44_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__44_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__44_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__44_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__44_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__44_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__44_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__45_ccff_tail ;
wire [0:19] cbx_1__1__45_chanx_left_out ;
wire [0:19] cbx_1__1__45_chanx_right_out ;
wire [0:0] cbx_1__1__45_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__45_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__45_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__45_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__45_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__45_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__45_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__45_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__45_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__45_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__45_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__45_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__45_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__45_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__45_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__45_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__46_ccff_tail ;
wire [0:19] cbx_1__1__46_chanx_left_out ;
wire [0:19] cbx_1__1__46_chanx_right_out ;
wire [0:0] cbx_1__1__46_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__46_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__46_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__46_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__46_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__46_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__46_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__46_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__46_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__46_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__46_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__46_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__46_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__46_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__46_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__46_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__47_ccff_tail ;
wire [0:19] cbx_1__1__47_chanx_left_out ;
wire [0:19] cbx_1__1__47_chanx_right_out ;
wire [0:0] cbx_1__1__47_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__47_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__47_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__47_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__47_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__47_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__47_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__47_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__47_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__47_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__47_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__47_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__47_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__47_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__47_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__47_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__48_ccff_tail ;
wire [0:19] cbx_1__1__48_chanx_left_out ;
wire [0:19] cbx_1__1__48_chanx_right_out ;
wire [0:0] cbx_1__1__48_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__48_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__48_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__48_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__48_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__48_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__48_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__48_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__48_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__48_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__48_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__48_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__48_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__48_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__48_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__48_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__49_ccff_tail ;
wire [0:19] cbx_1__1__49_chanx_left_out ;
wire [0:19] cbx_1__1__49_chanx_right_out ;
wire [0:0] cbx_1__1__49_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__49_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__49_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__49_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__49_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__49_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__49_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__49_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__49_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__49_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__49_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__49_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__49_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__49_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__49_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__49_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__4_ccff_tail ;
wire [0:19] cbx_1__1__4_chanx_left_out ;
wire [0:19] cbx_1__1__4_chanx_right_out ;
wire [0:0] cbx_1__1__4_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__4_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__4_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__4_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__4_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__4_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__4_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__4_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__4_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__4_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__4_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__4_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__4_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__4_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__4_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__4_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__50_ccff_tail ;
wire [0:19] cbx_1__1__50_chanx_left_out ;
wire [0:19] cbx_1__1__50_chanx_right_out ;
wire [0:0] cbx_1__1__50_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__50_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__50_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__50_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__50_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__50_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__50_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__50_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__50_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__50_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__50_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__50_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__50_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__50_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__50_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__50_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__51_ccff_tail ;
wire [0:19] cbx_1__1__51_chanx_left_out ;
wire [0:19] cbx_1__1__51_chanx_right_out ;
wire [0:0] cbx_1__1__51_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__51_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__51_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__51_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__51_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__51_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__51_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__51_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__51_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__51_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__51_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__51_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__51_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__51_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__51_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__51_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__52_ccff_tail ;
wire [0:19] cbx_1__1__52_chanx_left_out ;
wire [0:19] cbx_1__1__52_chanx_right_out ;
wire [0:0] cbx_1__1__52_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__52_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__52_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__52_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__52_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__52_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__52_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__52_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__52_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__52_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__52_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__52_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__52_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__52_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__52_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__52_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__53_ccff_tail ;
wire [0:19] cbx_1__1__53_chanx_left_out ;
wire [0:19] cbx_1__1__53_chanx_right_out ;
wire [0:0] cbx_1__1__53_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__53_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__53_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__53_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__53_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__53_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__53_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__53_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__53_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__53_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__53_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__53_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__53_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__53_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__53_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__53_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__54_ccff_tail ;
wire [0:19] cbx_1__1__54_chanx_left_out ;
wire [0:19] cbx_1__1__54_chanx_right_out ;
wire [0:0] cbx_1__1__54_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__54_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__54_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__54_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__54_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__54_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__54_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__54_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__54_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__54_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__54_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__54_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__54_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__54_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__54_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__54_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__55_ccff_tail ;
wire [0:19] cbx_1__1__55_chanx_left_out ;
wire [0:19] cbx_1__1__55_chanx_right_out ;
wire [0:0] cbx_1__1__55_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__55_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__55_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__55_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__55_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__55_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__55_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__55_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__55_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__55_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__55_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__55_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__55_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__55_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__55_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__55_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__56_ccff_tail ;
wire [0:19] cbx_1__1__56_chanx_left_out ;
wire [0:19] cbx_1__1__56_chanx_right_out ;
wire [0:0] cbx_1__1__56_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__56_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__56_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__56_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__56_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__56_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__56_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__56_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__56_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__56_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__56_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__56_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__56_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__56_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__56_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__56_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__57_ccff_tail ;
wire [0:19] cbx_1__1__57_chanx_left_out ;
wire [0:19] cbx_1__1__57_chanx_right_out ;
wire [0:0] cbx_1__1__57_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__57_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__57_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__57_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__57_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__57_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__57_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__57_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__57_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__57_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__57_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__57_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__57_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__57_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__57_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__57_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__58_ccff_tail ;
wire [0:19] cbx_1__1__58_chanx_left_out ;
wire [0:19] cbx_1__1__58_chanx_right_out ;
wire [0:0] cbx_1__1__58_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__58_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__58_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__58_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__58_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__58_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__58_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__58_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__58_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__58_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__58_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__58_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__58_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__58_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__58_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__58_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__59_ccff_tail ;
wire [0:19] cbx_1__1__59_chanx_left_out ;
wire [0:19] cbx_1__1__59_chanx_right_out ;
wire [0:0] cbx_1__1__59_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__59_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__59_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__59_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__59_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__59_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__59_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__59_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__59_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__59_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__59_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__59_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__59_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__59_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__59_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__59_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__5_ccff_tail ;
wire [0:19] cbx_1__1__5_chanx_left_out ;
wire [0:19] cbx_1__1__5_chanx_right_out ;
wire [0:0] cbx_1__1__5_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__5_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__5_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__5_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__5_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__5_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__5_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__5_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__5_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__5_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__5_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__5_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__5_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__5_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__5_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__5_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__60_ccff_tail ;
wire [0:19] cbx_1__1__60_chanx_left_out ;
wire [0:19] cbx_1__1__60_chanx_right_out ;
wire [0:0] cbx_1__1__60_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__60_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__60_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__60_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__60_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__60_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__60_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__60_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__60_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__60_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__60_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__60_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__60_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__60_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__60_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__60_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__61_ccff_tail ;
wire [0:19] cbx_1__1__61_chanx_left_out ;
wire [0:19] cbx_1__1__61_chanx_right_out ;
wire [0:0] cbx_1__1__61_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__61_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__61_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__61_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__61_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__61_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__61_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__61_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__61_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__61_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__61_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__61_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__61_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__61_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__61_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__61_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__62_ccff_tail ;
wire [0:19] cbx_1__1__62_chanx_left_out ;
wire [0:19] cbx_1__1__62_chanx_right_out ;
wire [0:0] cbx_1__1__62_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__62_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__62_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__62_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__62_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__62_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__62_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__62_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__62_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__62_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__62_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__62_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__62_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__62_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__62_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__62_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__63_ccff_tail ;
wire [0:19] cbx_1__1__63_chanx_left_out ;
wire [0:19] cbx_1__1__63_chanx_right_out ;
wire [0:0] cbx_1__1__63_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__63_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__63_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__63_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__63_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__63_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__63_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__63_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__63_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__63_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__63_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__63_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__63_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__63_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__63_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__63_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__64_ccff_tail ;
wire [0:19] cbx_1__1__64_chanx_left_out ;
wire [0:19] cbx_1__1__64_chanx_right_out ;
wire [0:0] cbx_1__1__64_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__64_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__64_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__64_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__64_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__64_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__64_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__64_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__64_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__64_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__64_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__64_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__64_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__64_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__64_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__64_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__65_ccff_tail ;
wire [0:19] cbx_1__1__65_chanx_left_out ;
wire [0:19] cbx_1__1__65_chanx_right_out ;
wire [0:0] cbx_1__1__65_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__65_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__65_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__65_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__65_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__65_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__65_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__65_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__65_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__65_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__65_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__65_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__65_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__65_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__65_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__65_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__66_ccff_tail ;
wire [0:19] cbx_1__1__66_chanx_left_out ;
wire [0:19] cbx_1__1__66_chanx_right_out ;
wire [0:0] cbx_1__1__66_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__66_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__66_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__66_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__66_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__66_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__66_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__66_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__66_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__66_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__66_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__66_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__66_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__66_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__66_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__66_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__67_ccff_tail ;
wire [0:19] cbx_1__1__67_chanx_left_out ;
wire [0:19] cbx_1__1__67_chanx_right_out ;
wire [0:0] cbx_1__1__67_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__67_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__67_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__67_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__67_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__67_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__67_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__67_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__67_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__67_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__67_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__67_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__67_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__67_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__67_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__67_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__68_ccff_tail ;
wire [0:19] cbx_1__1__68_chanx_left_out ;
wire [0:19] cbx_1__1__68_chanx_right_out ;
wire [0:0] cbx_1__1__68_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__68_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__68_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__68_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__68_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__68_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__68_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__68_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__68_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__68_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__68_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__68_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__68_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__68_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__68_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__68_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__69_ccff_tail ;
wire [0:19] cbx_1__1__69_chanx_left_out ;
wire [0:19] cbx_1__1__69_chanx_right_out ;
wire [0:0] cbx_1__1__69_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__69_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__69_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__69_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__69_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__69_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__69_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__69_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__69_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__69_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__69_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__69_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__69_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__69_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__69_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__69_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__6_ccff_tail ;
wire [0:19] cbx_1__1__6_chanx_left_out ;
wire [0:19] cbx_1__1__6_chanx_right_out ;
wire [0:0] cbx_1__1__6_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__6_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__6_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__6_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__6_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__6_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__6_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__6_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__6_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__6_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__6_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__6_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__6_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__6_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__6_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__6_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__70_ccff_tail ;
wire [0:19] cbx_1__1__70_chanx_left_out ;
wire [0:19] cbx_1__1__70_chanx_right_out ;
wire [0:0] cbx_1__1__70_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__70_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__70_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__70_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__70_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__70_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__70_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__70_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__70_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__70_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__70_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__70_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__70_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__70_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__70_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__70_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__71_ccff_tail ;
wire [0:19] cbx_1__1__71_chanx_left_out ;
wire [0:19] cbx_1__1__71_chanx_right_out ;
wire [0:0] cbx_1__1__71_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__71_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__71_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__71_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__71_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__71_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__71_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__71_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__71_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__71_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__71_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__71_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__71_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__71_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__71_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__71_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__72_ccff_tail ;
wire [0:19] cbx_1__1__72_chanx_left_out ;
wire [0:19] cbx_1__1__72_chanx_right_out ;
wire [0:0] cbx_1__1__72_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__72_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__72_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__72_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__72_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__72_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__72_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__72_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__72_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__72_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__72_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__72_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__72_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__72_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__72_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__72_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__73_ccff_tail ;
wire [0:19] cbx_1__1__73_chanx_left_out ;
wire [0:19] cbx_1__1__73_chanx_right_out ;
wire [0:0] cbx_1__1__73_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__73_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__73_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__73_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__73_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__73_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__73_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__73_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__73_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__73_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__73_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__73_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__73_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__73_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__73_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__73_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__74_ccff_tail ;
wire [0:19] cbx_1__1__74_chanx_left_out ;
wire [0:19] cbx_1__1__74_chanx_right_out ;
wire [0:0] cbx_1__1__74_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__74_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__74_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__74_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__74_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__74_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__74_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__74_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__74_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__74_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__74_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__74_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__74_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__74_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__74_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__74_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__75_ccff_tail ;
wire [0:19] cbx_1__1__75_chanx_left_out ;
wire [0:19] cbx_1__1__75_chanx_right_out ;
wire [0:0] cbx_1__1__75_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__75_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__75_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__75_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__75_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__75_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__75_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__75_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__75_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__75_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__75_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__75_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__75_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__75_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__75_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__75_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__76_ccff_tail ;
wire [0:19] cbx_1__1__76_chanx_left_out ;
wire [0:19] cbx_1__1__76_chanx_right_out ;
wire [0:0] cbx_1__1__76_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__76_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__76_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__76_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__76_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__76_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__76_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__76_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__76_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__76_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__76_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__76_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__76_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__76_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__76_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__76_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__77_ccff_tail ;
wire [0:19] cbx_1__1__77_chanx_left_out ;
wire [0:19] cbx_1__1__77_chanx_right_out ;
wire [0:0] cbx_1__1__77_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__77_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__77_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__77_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__77_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__77_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__77_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__77_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__77_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__77_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__77_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__77_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__77_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__77_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__77_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__77_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__78_ccff_tail ;
wire [0:19] cbx_1__1__78_chanx_left_out ;
wire [0:19] cbx_1__1__78_chanx_right_out ;
wire [0:0] cbx_1__1__78_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__78_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__78_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__78_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__78_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__78_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__78_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__78_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__78_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__78_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__78_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__78_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__78_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__78_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__78_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__78_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__79_ccff_tail ;
wire [0:19] cbx_1__1__79_chanx_left_out ;
wire [0:19] cbx_1__1__79_chanx_right_out ;
wire [0:0] cbx_1__1__79_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__79_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__79_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__79_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__79_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__79_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__79_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__79_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__79_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__79_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__79_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__79_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__79_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__79_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__79_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__79_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__7_ccff_tail ;
wire [0:19] cbx_1__1__7_chanx_left_out ;
wire [0:19] cbx_1__1__7_chanx_right_out ;
wire [0:0] cbx_1__1__7_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__7_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__7_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__7_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__7_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__7_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__7_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__7_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__7_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__7_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__7_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__7_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__7_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__7_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__7_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__7_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__80_ccff_tail ;
wire [0:19] cbx_1__1__80_chanx_left_out ;
wire [0:19] cbx_1__1__80_chanx_right_out ;
wire [0:0] cbx_1__1__80_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__80_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__80_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__80_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__80_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__80_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__80_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__80_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__80_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__80_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__80_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__80_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__80_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__80_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__80_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__80_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__81_ccff_tail ;
wire [0:19] cbx_1__1__81_chanx_left_out ;
wire [0:19] cbx_1__1__81_chanx_right_out ;
wire [0:0] cbx_1__1__81_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__81_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__81_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__81_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__81_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__81_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__81_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__81_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__81_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__81_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__81_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__81_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__81_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__81_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__81_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__81_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__82_ccff_tail ;
wire [0:19] cbx_1__1__82_chanx_left_out ;
wire [0:19] cbx_1__1__82_chanx_right_out ;
wire [0:0] cbx_1__1__82_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__82_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__82_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__82_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__82_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__82_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__82_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__82_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__82_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__82_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__82_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__82_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__82_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__82_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__82_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__82_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__83_ccff_tail ;
wire [0:19] cbx_1__1__83_chanx_left_out ;
wire [0:19] cbx_1__1__83_chanx_right_out ;
wire [0:0] cbx_1__1__83_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__83_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__83_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__83_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__83_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__83_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__83_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__83_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__83_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__83_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__83_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__83_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__83_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__83_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__83_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__83_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__84_ccff_tail ;
wire [0:19] cbx_1__1__84_chanx_left_out ;
wire [0:19] cbx_1__1__84_chanx_right_out ;
wire [0:0] cbx_1__1__84_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__84_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__84_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__84_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__84_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__84_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__84_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__84_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__84_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__84_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__84_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__84_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__84_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__84_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__84_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__84_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__85_ccff_tail ;
wire [0:19] cbx_1__1__85_chanx_left_out ;
wire [0:19] cbx_1__1__85_chanx_right_out ;
wire [0:0] cbx_1__1__85_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__85_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__85_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__85_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__85_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__85_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__85_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__85_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__85_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__85_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__85_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__85_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__85_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__85_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__85_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__85_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__86_ccff_tail ;
wire [0:19] cbx_1__1__86_chanx_left_out ;
wire [0:19] cbx_1__1__86_chanx_right_out ;
wire [0:0] cbx_1__1__86_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__86_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__86_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__86_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__86_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__86_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__86_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__86_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__86_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__86_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__86_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__86_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__86_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__86_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__86_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__86_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__87_ccff_tail ;
wire [0:19] cbx_1__1__87_chanx_left_out ;
wire [0:19] cbx_1__1__87_chanx_right_out ;
wire [0:0] cbx_1__1__87_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__87_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__87_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__87_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__87_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__87_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__87_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__87_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__87_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__87_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__87_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__87_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__87_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__87_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__87_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__87_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__88_ccff_tail ;
wire [0:19] cbx_1__1__88_chanx_left_out ;
wire [0:19] cbx_1__1__88_chanx_right_out ;
wire [0:0] cbx_1__1__88_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__88_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__88_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__88_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__88_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__88_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__88_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__88_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__88_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__88_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__88_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__88_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__88_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__88_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__88_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__88_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__89_ccff_tail ;
wire [0:19] cbx_1__1__89_chanx_left_out ;
wire [0:19] cbx_1__1__89_chanx_right_out ;
wire [0:0] cbx_1__1__89_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__89_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__89_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__89_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__89_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__89_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__89_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__89_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__89_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__89_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__89_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__89_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__89_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__89_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__89_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__89_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__8_ccff_tail ;
wire [0:19] cbx_1__1__8_chanx_left_out ;
wire [0:19] cbx_1__1__8_chanx_right_out ;
wire [0:0] cbx_1__1__8_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__8_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__8_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__8_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__8_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__8_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__8_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__8_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__8_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__8_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__8_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__8_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__8_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__8_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__8_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__8_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__90_ccff_tail ;
wire [0:19] cbx_1__1__90_chanx_left_out ;
wire [0:19] cbx_1__1__90_chanx_right_out ;
wire [0:0] cbx_1__1__90_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__90_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__90_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__90_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__90_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__90_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__90_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__90_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__90_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__90_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__90_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__90_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__90_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__90_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__90_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__90_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__91_ccff_tail ;
wire [0:19] cbx_1__1__91_chanx_left_out ;
wire [0:19] cbx_1__1__91_chanx_right_out ;
wire [0:0] cbx_1__1__91_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__91_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__91_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__91_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__91_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__91_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__91_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__91_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__91_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__91_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__91_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__91_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__91_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__91_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__91_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__91_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__92_ccff_tail ;
wire [0:19] cbx_1__1__92_chanx_left_out ;
wire [0:19] cbx_1__1__92_chanx_right_out ;
wire [0:0] cbx_1__1__92_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__92_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__92_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__92_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__92_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__92_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__92_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__92_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__92_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__92_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__92_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__92_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__92_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__92_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__92_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__92_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__93_ccff_tail ;
wire [0:19] cbx_1__1__93_chanx_left_out ;
wire [0:19] cbx_1__1__93_chanx_right_out ;
wire [0:0] cbx_1__1__93_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__93_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__93_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__93_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__93_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__93_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__93_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__93_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__93_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__93_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__93_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__93_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__93_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__93_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__93_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__93_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__94_ccff_tail ;
wire [0:19] cbx_1__1__94_chanx_left_out ;
wire [0:19] cbx_1__1__94_chanx_right_out ;
wire [0:0] cbx_1__1__94_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__94_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__94_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__94_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__94_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__94_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__94_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__94_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__94_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__94_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__94_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__94_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__94_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__94_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__94_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__94_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__95_ccff_tail ;
wire [0:19] cbx_1__1__95_chanx_left_out ;
wire [0:19] cbx_1__1__95_chanx_right_out ;
wire [0:0] cbx_1__1__95_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__95_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__95_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__95_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__95_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__95_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__95_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__95_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__95_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__95_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__95_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__95_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__95_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__95_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__95_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__95_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__96_ccff_tail ;
wire [0:19] cbx_1__1__96_chanx_left_out ;
wire [0:19] cbx_1__1__96_chanx_right_out ;
wire [0:0] cbx_1__1__96_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__96_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__96_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__96_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__96_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__96_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__96_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__96_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__96_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__96_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__96_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__96_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__96_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__96_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__96_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__96_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__97_ccff_tail ;
wire [0:19] cbx_1__1__97_chanx_left_out ;
wire [0:19] cbx_1__1__97_chanx_right_out ;
wire [0:0] cbx_1__1__97_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__97_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__97_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__97_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__97_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__97_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__97_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__97_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__97_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__97_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__97_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__97_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__97_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__97_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__97_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__97_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__98_ccff_tail ;
wire [0:19] cbx_1__1__98_chanx_left_out ;
wire [0:19] cbx_1__1__98_chanx_right_out ;
wire [0:0] cbx_1__1__98_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__98_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__98_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__98_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__98_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__98_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__98_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__98_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__98_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__98_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__98_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__98_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__98_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__98_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__98_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__98_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__99_ccff_tail ;
wire [0:19] cbx_1__1__99_chanx_left_out ;
wire [0:19] cbx_1__1__99_chanx_right_out ;
wire [0:0] cbx_1__1__99_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__99_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__99_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__99_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__99_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__99_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__99_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__99_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__99_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__99_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__99_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__99_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__99_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__99_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__99_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__99_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__9_ccff_tail ;
wire [0:19] cbx_1__1__9_chanx_left_out ;
wire [0:19] cbx_1__1__9_chanx_right_out ;
wire [0:0] cbx_1__1__9_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__9_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__9_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__9_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__9_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__9_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__9_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__9_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__9_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__9_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__9_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__9_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__9_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__9_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__9_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__9_top_grid_pin_31_ ;
wire [0:0] cby_0__1__0_ccff_tail ;
wire [0:19] cby_0__1__0_chany_bottom_out ;
wire [0:19] cby_0__1__0_chany_top_out ;
wire [0:0] cby_0__1__0_left_grid_pin_0_ ;
wire [0:0] cby_0__1__0_right_grid_pin_52_ ;
wire [0:0] cby_0__1__10_ccff_tail ;
wire [0:19] cby_0__1__10_chany_bottom_out ;
wire [0:19] cby_0__1__10_chany_top_out ;
wire [0:0] cby_0__1__10_left_grid_pin_0_ ;
wire [0:0] cby_0__1__10_right_grid_pin_52_ ;
wire [0:0] cby_0__1__11_ccff_tail ;
wire [0:19] cby_0__1__11_chany_bottom_out ;
wire [0:19] cby_0__1__11_chany_top_out ;
wire [0:0] cby_0__1__11_left_grid_pin_0_ ;
wire [0:0] cby_0__1__11_right_grid_pin_52_ ;
wire [0:0] cby_0__1__1_ccff_tail ;
wire [0:19] cby_0__1__1_chany_bottom_out ;
wire [0:19] cby_0__1__1_chany_top_out ;
wire [0:0] cby_0__1__1_left_grid_pin_0_ ;
wire [0:0] cby_0__1__1_right_grid_pin_52_ ;
wire [0:0] cby_0__1__2_ccff_tail ;
wire [0:19] cby_0__1__2_chany_bottom_out ;
wire [0:19] cby_0__1__2_chany_top_out ;
wire [0:0] cby_0__1__2_left_grid_pin_0_ ;
wire [0:0] cby_0__1__2_right_grid_pin_52_ ;
wire [0:0] cby_0__1__3_ccff_tail ;
wire [0:19] cby_0__1__3_chany_bottom_out ;
wire [0:19] cby_0__1__3_chany_top_out ;
wire [0:0] cby_0__1__3_left_grid_pin_0_ ;
wire [0:0] cby_0__1__3_right_grid_pin_52_ ;
wire [0:0] cby_0__1__4_ccff_tail ;
wire [0:19] cby_0__1__4_chany_bottom_out ;
wire [0:19] cby_0__1__4_chany_top_out ;
wire [0:0] cby_0__1__4_left_grid_pin_0_ ;
wire [0:0] cby_0__1__4_right_grid_pin_52_ ;
wire [0:0] cby_0__1__5_ccff_tail ;
wire [0:19] cby_0__1__5_chany_bottom_out ;
wire [0:19] cby_0__1__5_chany_top_out ;
wire [0:0] cby_0__1__5_left_grid_pin_0_ ;
wire [0:0] cby_0__1__5_right_grid_pin_52_ ;
wire [0:0] cby_0__1__6_ccff_tail ;
wire [0:19] cby_0__1__6_chany_bottom_out ;
wire [0:19] cby_0__1__6_chany_top_out ;
wire [0:0] cby_0__1__6_left_grid_pin_0_ ;
wire [0:0] cby_0__1__6_right_grid_pin_52_ ;
wire [0:0] cby_0__1__7_ccff_tail ;
wire [0:19] cby_0__1__7_chany_bottom_out ;
wire [0:19] cby_0__1__7_chany_top_out ;
wire [0:0] cby_0__1__7_left_grid_pin_0_ ;
wire [0:0] cby_0__1__7_right_grid_pin_52_ ;
wire [0:0] cby_0__1__8_ccff_tail ;
wire [0:19] cby_0__1__8_chany_bottom_out ;
wire [0:19] cby_0__1__8_chany_top_out ;
wire [0:0] cby_0__1__8_left_grid_pin_0_ ;
wire [0:0] cby_0__1__8_right_grid_pin_52_ ;
wire [0:0] cby_0__1__9_ccff_tail ;
wire [0:19] cby_0__1__9_chany_bottom_out ;
wire [0:19] cby_0__1__9_chany_top_out ;
wire [0:0] cby_0__1__9_left_grid_pin_0_ ;
wire [0:0] cby_0__1__9_right_grid_pin_52_ ;
wire [0:0] cby_1__1__0_ccff_tail ;
wire [0:19] cby_1__1__0_chany_bottom_out ;
wire [0:19] cby_1__1__0_chany_top_out ;
wire [0:0] cby_1__1__0_left_grid_pin_0_ ;
wire [0:0] cby_1__1__0_left_grid_pin_10_ ;
wire [0:0] cby_1__1__0_left_grid_pin_11_ ;
wire [0:0] cby_1__1__0_left_grid_pin_12_ ;
wire [0:0] cby_1__1__0_left_grid_pin_13_ ;
wire [0:0] cby_1__1__0_left_grid_pin_14_ ;
wire [0:0] cby_1__1__0_left_grid_pin_15_ ;
wire [0:0] cby_1__1__0_left_grid_pin_1_ ;
wire [0:0] cby_1__1__0_left_grid_pin_2_ ;
wire [0:0] cby_1__1__0_left_grid_pin_3_ ;
wire [0:0] cby_1__1__0_left_grid_pin_4_ ;
wire [0:0] cby_1__1__0_left_grid_pin_5_ ;
wire [0:0] cby_1__1__0_left_grid_pin_6_ ;
wire [0:0] cby_1__1__0_left_grid_pin_7_ ;
wire [0:0] cby_1__1__0_left_grid_pin_8_ ;
wire [0:0] cby_1__1__0_left_grid_pin_9_ ;
wire [0:0] cby_1__1__0_right_grid_pin_52_ ;
wire [0:0] cby_1__1__100_ccff_tail ;
wire [0:19] cby_1__1__100_chany_bottom_out ;
wire [0:19] cby_1__1__100_chany_top_out ;
wire [0:0] cby_1__1__100_left_grid_pin_0_ ;
wire [0:0] cby_1__1__100_left_grid_pin_10_ ;
wire [0:0] cby_1__1__100_left_grid_pin_11_ ;
wire [0:0] cby_1__1__100_left_grid_pin_12_ ;
wire [0:0] cby_1__1__100_left_grid_pin_13_ ;
wire [0:0] cby_1__1__100_left_grid_pin_14_ ;
wire [0:0] cby_1__1__100_left_grid_pin_15_ ;
wire [0:0] cby_1__1__100_left_grid_pin_1_ ;
wire [0:0] cby_1__1__100_left_grid_pin_2_ ;
wire [0:0] cby_1__1__100_left_grid_pin_3_ ;
wire [0:0] cby_1__1__100_left_grid_pin_4_ ;
wire [0:0] cby_1__1__100_left_grid_pin_5_ ;
wire [0:0] cby_1__1__100_left_grid_pin_6_ ;
wire [0:0] cby_1__1__100_left_grid_pin_7_ ;
wire [0:0] cby_1__1__100_left_grid_pin_8_ ;
wire [0:0] cby_1__1__100_left_grid_pin_9_ ;
wire [0:0] cby_1__1__100_right_grid_pin_52_ ;
wire [0:0] cby_1__1__101_ccff_tail ;
wire [0:19] cby_1__1__101_chany_bottom_out ;
wire [0:19] cby_1__1__101_chany_top_out ;
wire [0:0] cby_1__1__101_left_grid_pin_0_ ;
wire [0:0] cby_1__1__101_left_grid_pin_10_ ;
wire [0:0] cby_1__1__101_left_grid_pin_11_ ;
wire [0:0] cby_1__1__101_left_grid_pin_12_ ;
wire [0:0] cby_1__1__101_left_grid_pin_13_ ;
wire [0:0] cby_1__1__101_left_grid_pin_14_ ;
wire [0:0] cby_1__1__101_left_grid_pin_15_ ;
wire [0:0] cby_1__1__101_left_grid_pin_1_ ;
wire [0:0] cby_1__1__101_left_grid_pin_2_ ;
wire [0:0] cby_1__1__101_left_grid_pin_3_ ;
wire [0:0] cby_1__1__101_left_grid_pin_4_ ;
wire [0:0] cby_1__1__101_left_grid_pin_5_ ;
wire [0:0] cby_1__1__101_left_grid_pin_6_ ;
wire [0:0] cby_1__1__101_left_grid_pin_7_ ;
wire [0:0] cby_1__1__101_left_grid_pin_8_ ;
wire [0:0] cby_1__1__101_left_grid_pin_9_ ;
wire [0:0] cby_1__1__101_right_grid_pin_52_ ;
wire [0:0] cby_1__1__102_ccff_tail ;
wire [0:19] cby_1__1__102_chany_bottom_out ;
wire [0:19] cby_1__1__102_chany_top_out ;
wire [0:0] cby_1__1__102_left_grid_pin_0_ ;
wire [0:0] cby_1__1__102_left_grid_pin_10_ ;
wire [0:0] cby_1__1__102_left_grid_pin_11_ ;
wire [0:0] cby_1__1__102_left_grid_pin_12_ ;
wire [0:0] cby_1__1__102_left_grid_pin_13_ ;
wire [0:0] cby_1__1__102_left_grid_pin_14_ ;
wire [0:0] cby_1__1__102_left_grid_pin_15_ ;
wire [0:0] cby_1__1__102_left_grid_pin_1_ ;
wire [0:0] cby_1__1__102_left_grid_pin_2_ ;
wire [0:0] cby_1__1__102_left_grid_pin_3_ ;
wire [0:0] cby_1__1__102_left_grid_pin_4_ ;
wire [0:0] cby_1__1__102_left_grid_pin_5_ ;
wire [0:0] cby_1__1__102_left_grid_pin_6_ ;
wire [0:0] cby_1__1__102_left_grid_pin_7_ ;
wire [0:0] cby_1__1__102_left_grid_pin_8_ ;
wire [0:0] cby_1__1__102_left_grid_pin_9_ ;
wire [0:0] cby_1__1__102_right_grid_pin_52_ ;
wire [0:0] cby_1__1__103_ccff_tail ;
wire [0:19] cby_1__1__103_chany_bottom_out ;
wire [0:19] cby_1__1__103_chany_top_out ;
wire [0:0] cby_1__1__103_left_grid_pin_0_ ;
wire [0:0] cby_1__1__103_left_grid_pin_10_ ;
wire [0:0] cby_1__1__103_left_grid_pin_11_ ;
wire [0:0] cby_1__1__103_left_grid_pin_12_ ;
wire [0:0] cby_1__1__103_left_grid_pin_13_ ;
wire [0:0] cby_1__1__103_left_grid_pin_14_ ;
wire [0:0] cby_1__1__103_left_grid_pin_15_ ;
wire [0:0] cby_1__1__103_left_grid_pin_1_ ;
wire [0:0] cby_1__1__103_left_grid_pin_2_ ;
wire [0:0] cby_1__1__103_left_grid_pin_3_ ;
wire [0:0] cby_1__1__103_left_grid_pin_4_ ;
wire [0:0] cby_1__1__103_left_grid_pin_5_ ;
wire [0:0] cby_1__1__103_left_grid_pin_6_ ;
wire [0:0] cby_1__1__103_left_grid_pin_7_ ;
wire [0:0] cby_1__1__103_left_grid_pin_8_ ;
wire [0:0] cby_1__1__103_left_grid_pin_9_ ;
wire [0:0] cby_1__1__103_right_grid_pin_52_ ;
wire [0:0] cby_1__1__104_ccff_tail ;
wire [0:19] cby_1__1__104_chany_bottom_out ;
wire [0:19] cby_1__1__104_chany_top_out ;
wire [0:0] cby_1__1__104_left_grid_pin_0_ ;
wire [0:0] cby_1__1__104_left_grid_pin_10_ ;
wire [0:0] cby_1__1__104_left_grid_pin_11_ ;
wire [0:0] cby_1__1__104_left_grid_pin_12_ ;
wire [0:0] cby_1__1__104_left_grid_pin_13_ ;
wire [0:0] cby_1__1__104_left_grid_pin_14_ ;
wire [0:0] cby_1__1__104_left_grid_pin_15_ ;
wire [0:0] cby_1__1__104_left_grid_pin_1_ ;
wire [0:0] cby_1__1__104_left_grid_pin_2_ ;
wire [0:0] cby_1__1__104_left_grid_pin_3_ ;
wire [0:0] cby_1__1__104_left_grid_pin_4_ ;
wire [0:0] cby_1__1__104_left_grid_pin_5_ ;
wire [0:0] cby_1__1__104_left_grid_pin_6_ ;
wire [0:0] cby_1__1__104_left_grid_pin_7_ ;
wire [0:0] cby_1__1__104_left_grid_pin_8_ ;
wire [0:0] cby_1__1__104_left_grid_pin_9_ ;
wire [0:0] cby_1__1__104_right_grid_pin_52_ ;
wire [0:0] cby_1__1__105_ccff_tail ;
wire [0:19] cby_1__1__105_chany_bottom_out ;
wire [0:19] cby_1__1__105_chany_top_out ;
wire [0:0] cby_1__1__105_left_grid_pin_0_ ;
wire [0:0] cby_1__1__105_left_grid_pin_10_ ;
wire [0:0] cby_1__1__105_left_grid_pin_11_ ;
wire [0:0] cby_1__1__105_left_grid_pin_12_ ;
wire [0:0] cby_1__1__105_left_grid_pin_13_ ;
wire [0:0] cby_1__1__105_left_grid_pin_14_ ;
wire [0:0] cby_1__1__105_left_grid_pin_15_ ;
wire [0:0] cby_1__1__105_left_grid_pin_1_ ;
wire [0:0] cby_1__1__105_left_grid_pin_2_ ;
wire [0:0] cby_1__1__105_left_grid_pin_3_ ;
wire [0:0] cby_1__1__105_left_grid_pin_4_ ;
wire [0:0] cby_1__1__105_left_grid_pin_5_ ;
wire [0:0] cby_1__1__105_left_grid_pin_6_ ;
wire [0:0] cby_1__1__105_left_grid_pin_7_ ;
wire [0:0] cby_1__1__105_left_grid_pin_8_ ;
wire [0:0] cby_1__1__105_left_grid_pin_9_ ;
wire [0:0] cby_1__1__105_right_grid_pin_52_ ;
wire [0:0] cby_1__1__106_ccff_tail ;
wire [0:19] cby_1__1__106_chany_bottom_out ;
wire [0:19] cby_1__1__106_chany_top_out ;
wire [0:0] cby_1__1__106_left_grid_pin_0_ ;
wire [0:0] cby_1__1__106_left_grid_pin_10_ ;
wire [0:0] cby_1__1__106_left_grid_pin_11_ ;
wire [0:0] cby_1__1__106_left_grid_pin_12_ ;
wire [0:0] cby_1__1__106_left_grid_pin_13_ ;
wire [0:0] cby_1__1__106_left_grid_pin_14_ ;
wire [0:0] cby_1__1__106_left_grid_pin_15_ ;
wire [0:0] cby_1__1__106_left_grid_pin_1_ ;
wire [0:0] cby_1__1__106_left_grid_pin_2_ ;
wire [0:0] cby_1__1__106_left_grid_pin_3_ ;
wire [0:0] cby_1__1__106_left_grid_pin_4_ ;
wire [0:0] cby_1__1__106_left_grid_pin_5_ ;
wire [0:0] cby_1__1__106_left_grid_pin_6_ ;
wire [0:0] cby_1__1__106_left_grid_pin_7_ ;
wire [0:0] cby_1__1__106_left_grid_pin_8_ ;
wire [0:0] cby_1__1__106_left_grid_pin_9_ ;
wire [0:0] cby_1__1__106_right_grid_pin_52_ ;
wire [0:0] cby_1__1__107_ccff_tail ;
wire [0:19] cby_1__1__107_chany_bottom_out ;
wire [0:19] cby_1__1__107_chany_top_out ;
wire [0:0] cby_1__1__107_left_grid_pin_0_ ;
wire [0:0] cby_1__1__107_left_grid_pin_10_ ;
wire [0:0] cby_1__1__107_left_grid_pin_11_ ;
wire [0:0] cby_1__1__107_left_grid_pin_12_ ;
wire [0:0] cby_1__1__107_left_grid_pin_13_ ;
wire [0:0] cby_1__1__107_left_grid_pin_14_ ;
wire [0:0] cby_1__1__107_left_grid_pin_15_ ;
wire [0:0] cby_1__1__107_left_grid_pin_1_ ;
wire [0:0] cby_1__1__107_left_grid_pin_2_ ;
wire [0:0] cby_1__1__107_left_grid_pin_3_ ;
wire [0:0] cby_1__1__107_left_grid_pin_4_ ;
wire [0:0] cby_1__1__107_left_grid_pin_5_ ;
wire [0:0] cby_1__1__107_left_grid_pin_6_ ;
wire [0:0] cby_1__1__107_left_grid_pin_7_ ;
wire [0:0] cby_1__1__107_left_grid_pin_8_ ;
wire [0:0] cby_1__1__107_left_grid_pin_9_ ;
wire [0:0] cby_1__1__107_right_grid_pin_52_ ;
wire [0:0] cby_1__1__108_ccff_tail ;
wire [0:19] cby_1__1__108_chany_bottom_out ;
wire [0:19] cby_1__1__108_chany_top_out ;
wire [0:0] cby_1__1__108_left_grid_pin_0_ ;
wire [0:0] cby_1__1__108_left_grid_pin_10_ ;
wire [0:0] cby_1__1__108_left_grid_pin_11_ ;
wire [0:0] cby_1__1__108_left_grid_pin_12_ ;
wire [0:0] cby_1__1__108_left_grid_pin_13_ ;
wire [0:0] cby_1__1__108_left_grid_pin_14_ ;
wire [0:0] cby_1__1__108_left_grid_pin_15_ ;
wire [0:0] cby_1__1__108_left_grid_pin_1_ ;
wire [0:0] cby_1__1__108_left_grid_pin_2_ ;
wire [0:0] cby_1__1__108_left_grid_pin_3_ ;
wire [0:0] cby_1__1__108_left_grid_pin_4_ ;
wire [0:0] cby_1__1__108_left_grid_pin_5_ ;
wire [0:0] cby_1__1__108_left_grid_pin_6_ ;
wire [0:0] cby_1__1__108_left_grid_pin_7_ ;
wire [0:0] cby_1__1__108_left_grid_pin_8_ ;
wire [0:0] cby_1__1__108_left_grid_pin_9_ ;
wire [0:0] cby_1__1__108_right_grid_pin_52_ ;
wire [0:0] cby_1__1__109_ccff_tail ;
wire [0:19] cby_1__1__109_chany_bottom_out ;
wire [0:19] cby_1__1__109_chany_top_out ;
wire [0:0] cby_1__1__109_left_grid_pin_0_ ;
wire [0:0] cby_1__1__109_left_grid_pin_10_ ;
wire [0:0] cby_1__1__109_left_grid_pin_11_ ;
wire [0:0] cby_1__1__109_left_grid_pin_12_ ;
wire [0:0] cby_1__1__109_left_grid_pin_13_ ;
wire [0:0] cby_1__1__109_left_grid_pin_14_ ;
wire [0:0] cby_1__1__109_left_grid_pin_15_ ;
wire [0:0] cby_1__1__109_left_grid_pin_1_ ;
wire [0:0] cby_1__1__109_left_grid_pin_2_ ;
wire [0:0] cby_1__1__109_left_grid_pin_3_ ;
wire [0:0] cby_1__1__109_left_grid_pin_4_ ;
wire [0:0] cby_1__1__109_left_grid_pin_5_ ;
wire [0:0] cby_1__1__109_left_grid_pin_6_ ;
wire [0:0] cby_1__1__109_left_grid_pin_7_ ;
wire [0:0] cby_1__1__109_left_grid_pin_8_ ;
wire [0:0] cby_1__1__109_left_grid_pin_9_ ;
wire [0:0] cby_1__1__109_right_grid_pin_52_ ;
wire [0:0] cby_1__1__10_ccff_tail ;
wire [0:19] cby_1__1__10_chany_bottom_out ;
wire [0:19] cby_1__1__10_chany_top_out ;
wire [0:0] cby_1__1__10_left_grid_pin_0_ ;
wire [0:0] cby_1__1__10_left_grid_pin_10_ ;
wire [0:0] cby_1__1__10_left_grid_pin_11_ ;
wire [0:0] cby_1__1__10_left_grid_pin_12_ ;
wire [0:0] cby_1__1__10_left_grid_pin_13_ ;
wire [0:0] cby_1__1__10_left_grid_pin_14_ ;
wire [0:0] cby_1__1__10_left_grid_pin_15_ ;
wire [0:0] cby_1__1__10_left_grid_pin_1_ ;
wire [0:0] cby_1__1__10_left_grid_pin_2_ ;
wire [0:0] cby_1__1__10_left_grid_pin_3_ ;
wire [0:0] cby_1__1__10_left_grid_pin_4_ ;
wire [0:0] cby_1__1__10_left_grid_pin_5_ ;
wire [0:0] cby_1__1__10_left_grid_pin_6_ ;
wire [0:0] cby_1__1__10_left_grid_pin_7_ ;
wire [0:0] cby_1__1__10_left_grid_pin_8_ ;
wire [0:0] cby_1__1__10_left_grid_pin_9_ ;
wire [0:0] cby_1__1__10_right_grid_pin_52_ ;
wire [0:0] cby_1__1__110_ccff_tail ;
wire [0:19] cby_1__1__110_chany_bottom_out ;
wire [0:19] cby_1__1__110_chany_top_out ;
wire [0:0] cby_1__1__110_left_grid_pin_0_ ;
wire [0:0] cby_1__1__110_left_grid_pin_10_ ;
wire [0:0] cby_1__1__110_left_grid_pin_11_ ;
wire [0:0] cby_1__1__110_left_grid_pin_12_ ;
wire [0:0] cby_1__1__110_left_grid_pin_13_ ;
wire [0:0] cby_1__1__110_left_grid_pin_14_ ;
wire [0:0] cby_1__1__110_left_grid_pin_15_ ;
wire [0:0] cby_1__1__110_left_grid_pin_1_ ;
wire [0:0] cby_1__1__110_left_grid_pin_2_ ;
wire [0:0] cby_1__1__110_left_grid_pin_3_ ;
wire [0:0] cby_1__1__110_left_grid_pin_4_ ;
wire [0:0] cby_1__1__110_left_grid_pin_5_ ;
wire [0:0] cby_1__1__110_left_grid_pin_6_ ;
wire [0:0] cby_1__1__110_left_grid_pin_7_ ;
wire [0:0] cby_1__1__110_left_grid_pin_8_ ;
wire [0:0] cby_1__1__110_left_grid_pin_9_ ;
wire [0:0] cby_1__1__110_right_grid_pin_52_ ;
wire [0:0] cby_1__1__111_ccff_tail ;
wire [0:19] cby_1__1__111_chany_bottom_out ;
wire [0:19] cby_1__1__111_chany_top_out ;
wire [0:0] cby_1__1__111_left_grid_pin_0_ ;
wire [0:0] cby_1__1__111_left_grid_pin_10_ ;
wire [0:0] cby_1__1__111_left_grid_pin_11_ ;
wire [0:0] cby_1__1__111_left_grid_pin_12_ ;
wire [0:0] cby_1__1__111_left_grid_pin_13_ ;
wire [0:0] cby_1__1__111_left_grid_pin_14_ ;
wire [0:0] cby_1__1__111_left_grid_pin_15_ ;
wire [0:0] cby_1__1__111_left_grid_pin_1_ ;
wire [0:0] cby_1__1__111_left_grid_pin_2_ ;
wire [0:0] cby_1__1__111_left_grid_pin_3_ ;
wire [0:0] cby_1__1__111_left_grid_pin_4_ ;
wire [0:0] cby_1__1__111_left_grid_pin_5_ ;
wire [0:0] cby_1__1__111_left_grid_pin_6_ ;
wire [0:0] cby_1__1__111_left_grid_pin_7_ ;
wire [0:0] cby_1__1__111_left_grid_pin_8_ ;
wire [0:0] cby_1__1__111_left_grid_pin_9_ ;
wire [0:0] cby_1__1__111_right_grid_pin_52_ ;
wire [0:0] cby_1__1__112_ccff_tail ;
wire [0:19] cby_1__1__112_chany_bottom_out ;
wire [0:19] cby_1__1__112_chany_top_out ;
wire [0:0] cby_1__1__112_left_grid_pin_0_ ;
wire [0:0] cby_1__1__112_left_grid_pin_10_ ;
wire [0:0] cby_1__1__112_left_grid_pin_11_ ;
wire [0:0] cby_1__1__112_left_grid_pin_12_ ;
wire [0:0] cby_1__1__112_left_grid_pin_13_ ;
wire [0:0] cby_1__1__112_left_grid_pin_14_ ;
wire [0:0] cby_1__1__112_left_grid_pin_15_ ;
wire [0:0] cby_1__1__112_left_grid_pin_1_ ;
wire [0:0] cby_1__1__112_left_grid_pin_2_ ;
wire [0:0] cby_1__1__112_left_grid_pin_3_ ;
wire [0:0] cby_1__1__112_left_grid_pin_4_ ;
wire [0:0] cby_1__1__112_left_grid_pin_5_ ;
wire [0:0] cby_1__1__112_left_grid_pin_6_ ;
wire [0:0] cby_1__1__112_left_grid_pin_7_ ;
wire [0:0] cby_1__1__112_left_grid_pin_8_ ;
wire [0:0] cby_1__1__112_left_grid_pin_9_ ;
wire [0:0] cby_1__1__112_right_grid_pin_52_ ;
wire [0:0] cby_1__1__113_ccff_tail ;
wire [0:19] cby_1__1__113_chany_bottom_out ;
wire [0:19] cby_1__1__113_chany_top_out ;
wire [0:0] cby_1__1__113_left_grid_pin_0_ ;
wire [0:0] cby_1__1__113_left_grid_pin_10_ ;
wire [0:0] cby_1__1__113_left_grid_pin_11_ ;
wire [0:0] cby_1__1__113_left_grid_pin_12_ ;
wire [0:0] cby_1__1__113_left_grid_pin_13_ ;
wire [0:0] cby_1__1__113_left_grid_pin_14_ ;
wire [0:0] cby_1__1__113_left_grid_pin_15_ ;
wire [0:0] cby_1__1__113_left_grid_pin_1_ ;
wire [0:0] cby_1__1__113_left_grid_pin_2_ ;
wire [0:0] cby_1__1__113_left_grid_pin_3_ ;
wire [0:0] cby_1__1__113_left_grid_pin_4_ ;
wire [0:0] cby_1__1__113_left_grid_pin_5_ ;
wire [0:0] cby_1__1__113_left_grid_pin_6_ ;
wire [0:0] cby_1__1__113_left_grid_pin_7_ ;
wire [0:0] cby_1__1__113_left_grid_pin_8_ ;
wire [0:0] cby_1__1__113_left_grid_pin_9_ ;
wire [0:0] cby_1__1__113_right_grid_pin_52_ ;
wire [0:0] cby_1__1__114_ccff_tail ;
wire [0:19] cby_1__1__114_chany_bottom_out ;
wire [0:19] cby_1__1__114_chany_top_out ;
wire [0:0] cby_1__1__114_left_grid_pin_0_ ;
wire [0:0] cby_1__1__114_left_grid_pin_10_ ;
wire [0:0] cby_1__1__114_left_grid_pin_11_ ;
wire [0:0] cby_1__1__114_left_grid_pin_12_ ;
wire [0:0] cby_1__1__114_left_grid_pin_13_ ;
wire [0:0] cby_1__1__114_left_grid_pin_14_ ;
wire [0:0] cby_1__1__114_left_grid_pin_15_ ;
wire [0:0] cby_1__1__114_left_grid_pin_1_ ;
wire [0:0] cby_1__1__114_left_grid_pin_2_ ;
wire [0:0] cby_1__1__114_left_grid_pin_3_ ;
wire [0:0] cby_1__1__114_left_grid_pin_4_ ;
wire [0:0] cby_1__1__114_left_grid_pin_5_ ;
wire [0:0] cby_1__1__114_left_grid_pin_6_ ;
wire [0:0] cby_1__1__114_left_grid_pin_7_ ;
wire [0:0] cby_1__1__114_left_grid_pin_8_ ;
wire [0:0] cby_1__1__114_left_grid_pin_9_ ;
wire [0:0] cby_1__1__114_right_grid_pin_52_ ;
wire [0:0] cby_1__1__115_ccff_tail ;
wire [0:19] cby_1__1__115_chany_bottom_out ;
wire [0:19] cby_1__1__115_chany_top_out ;
wire [0:0] cby_1__1__115_left_grid_pin_0_ ;
wire [0:0] cby_1__1__115_left_grid_pin_10_ ;
wire [0:0] cby_1__1__115_left_grid_pin_11_ ;
wire [0:0] cby_1__1__115_left_grid_pin_12_ ;
wire [0:0] cby_1__1__115_left_grid_pin_13_ ;
wire [0:0] cby_1__1__115_left_grid_pin_14_ ;
wire [0:0] cby_1__1__115_left_grid_pin_15_ ;
wire [0:0] cby_1__1__115_left_grid_pin_1_ ;
wire [0:0] cby_1__1__115_left_grid_pin_2_ ;
wire [0:0] cby_1__1__115_left_grid_pin_3_ ;
wire [0:0] cby_1__1__115_left_grid_pin_4_ ;
wire [0:0] cby_1__1__115_left_grid_pin_5_ ;
wire [0:0] cby_1__1__115_left_grid_pin_6_ ;
wire [0:0] cby_1__1__115_left_grid_pin_7_ ;
wire [0:0] cby_1__1__115_left_grid_pin_8_ ;
wire [0:0] cby_1__1__115_left_grid_pin_9_ ;
wire [0:0] cby_1__1__115_right_grid_pin_52_ ;
wire [0:0] cby_1__1__116_ccff_tail ;
wire [0:19] cby_1__1__116_chany_bottom_out ;
wire [0:19] cby_1__1__116_chany_top_out ;
wire [0:0] cby_1__1__116_left_grid_pin_0_ ;
wire [0:0] cby_1__1__116_left_grid_pin_10_ ;
wire [0:0] cby_1__1__116_left_grid_pin_11_ ;
wire [0:0] cby_1__1__116_left_grid_pin_12_ ;
wire [0:0] cby_1__1__116_left_grid_pin_13_ ;
wire [0:0] cby_1__1__116_left_grid_pin_14_ ;
wire [0:0] cby_1__1__116_left_grid_pin_15_ ;
wire [0:0] cby_1__1__116_left_grid_pin_1_ ;
wire [0:0] cby_1__1__116_left_grid_pin_2_ ;
wire [0:0] cby_1__1__116_left_grid_pin_3_ ;
wire [0:0] cby_1__1__116_left_grid_pin_4_ ;
wire [0:0] cby_1__1__116_left_grid_pin_5_ ;
wire [0:0] cby_1__1__116_left_grid_pin_6_ ;
wire [0:0] cby_1__1__116_left_grid_pin_7_ ;
wire [0:0] cby_1__1__116_left_grid_pin_8_ ;
wire [0:0] cby_1__1__116_left_grid_pin_9_ ;
wire [0:0] cby_1__1__116_right_grid_pin_52_ ;
wire [0:0] cby_1__1__117_ccff_tail ;
wire [0:19] cby_1__1__117_chany_bottom_out ;
wire [0:19] cby_1__1__117_chany_top_out ;
wire [0:0] cby_1__1__117_left_grid_pin_0_ ;
wire [0:0] cby_1__1__117_left_grid_pin_10_ ;
wire [0:0] cby_1__1__117_left_grid_pin_11_ ;
wire [0:0] cby_1__1__117_left_grid_pin_12_ ;
wire [0:0] cby_1__1__117_left_grid_pin_13_ ;
wire [0:0] cby_1__1__117_left_grid_pin_14_ ;
wire [0:0] cby_1__1__117_left_grid_pin_15_ ;
wire [0:0] cby_1__1__117_left_grid_pin_1_ ;
wire [0:0] cby_1__1__117_left_grid_pin_2_ ;
wire [0:0] cby_1__1__117_left_grid_pin_3_ ;
wire [0:0] cby_1__1__117_left_grid_pin_4_ ;
wire [0:0] cby_1__1__117_left_grid_pin_5_ ;
wire [0:0] cby_1__1__117_left_grid_pin_6_ ;
wire [0:0] cby_1__1__117_left_grid_pin_7_ ;
wire [0:0] cby_1__1__117_left_grid_pin_8_ ;
wire [0:0] cby_1__1__117_left_grid_pin_9_ ;
wire [0:0] cby_1__1__117_right_grid_pin_52_ ;
wire [0:0] cby_1__1__118_ccff_tail ;
wire [0:19] cby_1__1__118_chany_bottom_out ;
wire [0:19] cby_1__1__118_chany_top_out ;
wire [0:0] cby_1__1__118_left_grid_pin_0_ ;
wire [0:0] cby_1__1__118_left_grid_pin_10_ ;
wire [0:0] cby_1__1__118_left_grid_pin_11_ ;
wire [0:0] cby_1__1__118_left_grid_pin_12_ ;
wire [0:0] cby_1__1__118_left_grid_pin_13_ ;
wire [0:0] cby_1__1__118_left_grid_pin_14_ ;
wire [0:0] cby_1__1__118_left_grid_pin_15_ ;
wire [0:0] cby_1__1__118_left_grid_pin_1_ ;
wire [0:0] cby_1__1__118_left_grid_pin_2_ ;
wire [0:0] cby_1__1__118_left_grid_pin_3_ ;
wire [0:0] cby_1__1__118_left_grid_pin_4_ ;
wire [0:0] cby_1__1__118_left_grid_pin_5_ ;
wire [0:0] cby_1__1__118_left_grid_pin_6_ ;
wire [0:0] cby_1__1__118_left_grid_pin_7_ ;
wire [0:0] cby_1__1__118_left_grid_pin_8_ ;
wire [0:0] cby_1__1__118_left_grid_pin_9_ ;
wire [0:0] cby_1__1__118_right_grid_pin_52_ ;
wire [0:0] cby_1__1__119_ccff_tail ;
wire [0:19] cby_1__1__119_chany_bottom_out ;
wire [0:19] cby_1__1__119_chany_top_out ;
wire [0:0] cby_1__1__119_left_grid_pin_0_ ;
wire [0:0] cby_1__1__119_left_grid_pin_10_ ;
wire [0:0] cby_1__1__119_left_grid_pin_11_ ;
wire [0:0] cby_1__1__119_left_grid_pin_12_ ;
wire [0:0] cby_1__1__119_left_grid_pin_13_ ;
wire [0:0] cby_1__1__119_left_grid_pin_14_ ;
wire [0:0] cby_1__1__119_left_grid_pin_15_ ;
wire [0:0] cby_1__1__119_left_grid_pin_1_ ;
wire [0:0] cby_1__1__119_left_grid_pin_2_ ;
wire [0:0] cby_1__1__119_left_grid_pin_3_ ;
wire [0:0] cby_1__1__119_left_grid_pin_4_ ;
wire [0:0] cby_1__1__119_left_grid_pin_5_ ;
wire [0:0] cby_1__1__119_left_grid_pin_6_ ;
wire [0:0] cby_1__1__119_left_grid_pin_7_ ;
wire [0:0] cby_1__1__119_left_grid_pin_8_ ;
wire [0:0] cby_1__1__119_left_grid_pin_9_ ;
wire [0:0] cby_1__1__119_right_grid_pin_52_ ;
wire [0:0] cby_1__1__11_ccff_tail ;
wire [0:19] cby_1__1__11_chany_bottom_out ;
wire [0:19] cby_1__1__11_chany_top_out ;
wire [0:0] cby_1__1__11_left_grid_pin_0_ ;
wire [0:0] cby_1__1__11_left_grid_pin_10_ ;
wire [0:0] cby_1__1__11_left_grid_pin_11_ ;
wire [0:0] cby_1__1__11_left_grid_pin_12_ ;
wire [0:0] cby_1__1__11_left_grid_pin_13_ ;
wire [0:0] cby_1__1__11_left_grid_pin_14_ ;
wire [0:0] cby_1__1__11_left_grid_pin_15_ ;
wire [0:0] cby_1__1__11_left_grid_pin_1_ ;
wire [0:0] cby_1__1__11_left_grid_pin_2_ ;
wire [0:0] cby_1__1__11_left_grid_pin_3_ ;
wire [0:0] cby_1__1__11_left_grid_pin_4_ ;
wire [0:0] cby_1__1__11_left_grid_pin_5_ ;
wire [0:0] cby_1__1__11_left_grid_pin_6_ ;
wire [0:0] cby_1__1__11_left_grid_pin_7_ ;
wire [0:0] cby_1__1__11_left_grid_pin_8_ ;
wire [0:0] cby_1__1__11_left_grid_pin_9_ ;
wire [0:0] cby_1__1__11_right_grid_pin_52_ ;
wire [0:0] cby_1__1__120_ccff_tail ;
wire [0:19] cby_1__1__120_chany_bottom_out ;
wire [0:19] cby_1__1__120_chany_top_out ;
wire [0:0] cby_1__1__120_left_grid_pin_0_ ;
wire [0:0] cby_1__1__120_left_grid_pin_10_ ;
wire [0:0] cby_1__1__120_left_grid_pin_11_ ;
wire [0:0] cby_1__1__120_left_grid_pin_12_ ;
wire [0:0] cby_1__1__120_left_grid_pin_13_ ;
wire [0:0] cby_1__1__120_left_grid_pin_14_ ;
wire [0:0] cby_1__1__120_left_grid_pin_15_ ;
wire [0:0] cby_1__1__120_left_grid_pin_1_ ;
wire [0:0] cby_1__1__120_left_grid_pin_2_ ;
wire [0:0] cby_1__1__120_left_grid_pin_3_ ;
wire [0:0] cby_1__1__120_left_grid_pin_4_ ;
wire [0:0] cby_1__1__120_left_grid_pin_5_ ;
wire [0:0] cby_1__1__120_left_grid_pin_6_ ;
wire [0:0] cby_1__1__120_left_grid_pin_7_ ;
wire [0:0] cby_1__1__120_left_grid_pin_8_ ;
wire [0:0] cby_1__1__120_left_grid_pin_9_ ;
wire [0:0] cby_1__1__120_right_grid_pin_52_ ;
wire [0:0] cby_1__1__121_ccff_tail ;
wire [0:19] cby_1__1__121_chany_bottom_out ;
wire [0:19] cby_1__1__121_chany_top_out ;
wire [0:0] cby_1__1__121_left_grid_pin_0_ ;
wire [0:0] cby_1__1__121_left_grid_pin_10_ ;
wire [0:0] cby_1__1__121_left_grid_pin_11_ ;
wire [0:0] cby_1__1__121_left_grid_pin_12_ ;
wire [0:0] cby_1__1__121_left_grid_pin_13_ ;
wire [0:0] cby_1__1__121_left_grid_pin_14_ ;
wire [0:0] cby_1__1__121_left_grid_pin_15_ ;
wire [0:0] cby_1__1__121_left_grid_pin_1_ ;
wire [0:0] cby_1__1__121_left_grid_pin_2_ ;
wire [0:0] cby_1__1__121_left_grid_pin_3_ ;
wire [0:0] cby_1__1__121_left_grid_pin_4_ ;
wire [0:0] cby_1__1__121_left_grid_pin_5_ ;
wire [0:0] cby_1__1__121_left_grid_pin_6_ ;
wire [0:0] cby_1__1__121_left_grid_pin_7_ ;
wire [0:0] cby_1__1__121_left_grid_pin_8_ ;
wire [0:0] cby_1__1__121_left_grid_pin_9_ ;
wire [0:0] cby_1__1__121_right_grid_pin_52_ ;
wire [0:0] cby_1__1__122_ccff_tail ;
wire [0:19] cby_1__1__122_chany_bottom_out ;
wire [0:19] cby_1__1__122_chany_top_out ;
wire [0:0] cby_1__1__122_left_grid_pin_0_ ;
wire [0:0] cby_1__1__122_left_grid_pin_10_ ;
wire [0:0] cby_1__1__122_left_grid_pin_11_ ;
wire [0:0] cby_1__1__122_left_grid_pin_12_ ;
wire [0:0] cby_1__1__122_left_grid_pin_13_ ;
wire [0:0] cby_1__1__122_left_grid_pin_14_ ;
wire [0:0] cby_1__1__122_left_grid_pin_15_ ;
wire [0:0] cby_1__1__122_left_grid_pin_1_ ;
wire [0:0] cby_1__1__122_left_grid_pin_2_ ;
wire [0:0] cby_1__1__122_left_grid_pin_3_ ;
wire [0:0] cby_1__1__122_left_grid_pin_4_ ;
wire [0:0] cby_1__1__122_left_grid_pin_5_ ;
wire [0:0] cby_1__1__122_left_grid_pin_6_ ;
wire [0:0] cby_1__1__122_left_grid_pin_7_ ;
wire [0:0] cby_1__1__122_left_grid_pin_8_ ;
wire [0:0] cby_1__1__122_left_grid_pin_9_ ;
wire [0:0] cby_1__1__122_right_grid_pin_52_ ;
wire [0:0] cby_1__1__123_ccff_tail ;
wire [0:19] cby_1__1__123_chany_bottom_out ;
wire [0:19] cby_1__1__123_chany_top_out ;
wire [0:0] cby_1__1__123_left_grid_pin_0_ ;
wire [0:0] cby_1__1__123_left_grid_pin_10_ ;
wire [0:0] cby_1__1__123_left_grid_pin_11_ ;
wire [0:0] cby_1__1__123_left_grid_pin_12_ ;
wire [0:0] cby_1__1__123_left_grid_pin_13_ ;
wire [0:0] cby_1__1__123_left_grid_pin_14_ ;
wire [0:0] cby_1__1__123_left_grid_pin_15_ ;
wire [0:0] cby_1__1__123_left_grid_pin_1_ ;
wire [0:0] cby_1__1__123_left_grid_pin_2_ ;
wire [0:0] cby_1__1__123_left_grid_pin_3_ ;
wire [0:0] cby_1__1__123_left_grid_pin_4_ ;
wire [0:0] cby_1__1__123_left_grid_pin_5_ ;
wire [0:0] cby_1__1__123_left_grid_pin_6_ ;
wire [0:0] cby_1__1__123_left_grid_pin_7_ ;
wire [0:0] cby_1__1__123_left_grid_pin_8_ ;
wire [0:0] cby_1__1__123_left_grid_pin_9_ ;
wire [0:0] cby_1__1__123_right_grid_pin_52_ ;
wire [0:0] cby_1__1__124_ccff_tail ;
wire [0:19] cby_1__1__124_chany_bottom_out ;
wire [0:19] cby_1__1__124_chany_top_out ;
wire [0:0] cby_1__1__124_left_grid_pin_0_ ;
wire [0:0] cby_1__1__124_left_grid_pin_10_ ;
wire [0:0] cby_1__1__124_left_grid_pin_11_ ;
wire [0:0] cby_1__1__124_left_grid_pin_12_ ;
wire [0:0] cby_1__1__124_left_grid_pin_13_ ;
wire [0:0] cby_1__1__124_left_grid_pin_14_ ;
wire [0:0] cby_1__1__124_left_grid_pin_15_ ;
wire [0:0] cby_1__1__124_left_grid_pin_1_ ;
wire [0:0] cby_1__1__124_left_grid_pin_2_ ;
wire [0:0] cby_1__1__124_left_grid_pin_3_ ;
wire [0:0] cby_1__1__124_left_grid_pin_4_ ;
wire [0:0] cby_1__1__124_left_grid_pin_5_ ;
wire [0:0] cby_1__1__124_left_grid_pin_6_ ;
wire [0:0] cby_1__1__124_left_grid_pin_7_ ;
wire [0:0] cby_1__1__124_left_grid_pin_8_ ;
wire [0:0] cby_1__1__124_left_grid_pin_9_ ;
wire [0:0] cby_1__1__124_right_grid_pin_52_ ;
wire [0:0] cby_1__1__125_ccff_tail ;
wire [0:19] cby_1__1__125_chany_bottom_out ;
wire [0:19] cby_1__1__125_chany_top_out ;
wire [0:0] cby_1__1__125_left_grid_pin_0_ ;
wire [0:0] cby_1__1__125_left_grid_pin_10_ ;
wire [0:0] cby_1__1__125_left_grid_pin_11_ ;
wire [0:0] cby_1__1__125_left_grid_pin_12_ ;
wire [0:0] cby_1__1__125_left_grid_pin_13_ ;
wire [0:0] cby_1__1__125_left_grid_pin_14_ ;
wire [0:0] cby_1__1__125_left_grid_pin_15_ ;
wire [0:0] cby_1__1__125_left_grid_pin_1_ ;
wire [0:0] cby_1__1__125_left_grid_pin_2_ ;
wire [0:0] cby_1__1__125_left_grid_pin_3_ ;
wire [0:0] cby_1__1__125_left_grid_pin_4_ ;
wire [0:0] cby_1__1__125_left_grid_pin_5_ ;
wire [0:0] cby_1__1__125_left_grid_pin_6_ ;
wire [0:0] cby_1__1__125_left_grid_pin_7_ ;
wire [0:0] cby_1__1__125_left_grid_pin_8_ ;
wire [0:0] cby_1__1__125_left_grid_pin_9_ ;
wire [0:0] cby_1__1__125_right_grid_pin_52_ ;
wire [0:0] cby_1__1__126_ccff_tail ;
wire [0:19] cby_1__1__126_chany_bottom_out ;
wire [0:19] cby_1__1__126_chany_top_out ;
wire [0:0] cby_1__1__126_left_grid_pin_0_ ;
wire [0:0] cby_1__1__126_left_grid_pin_10_ ;
wire [0:0] cby_1__1__126_left_grid_pin_11_ ;
wire [0:0] cby_1__1__126_left_grid_pin_12_ ;
wire [0:0] cby_1__1__126_left_grid_pin_13_ ;
wire [0:0] cby_1__1__126_left_grid_pin_14_ ;
wire [0:0] cby_1__1__126_left_grid_pin_15_ ;
wire [0:0] cby_1__1__126_left_grid_pin_1_ ;
wire [0:0] cby_1__1__126_left_grid_pin_2_ ;
wire [0:0] cby_1__1__126_left_grid_pin_3_ ;
wire [0:0] cby_1__1__126_left_grid_pin_4_ ;
wire [0:0] cby_1__1__126_left_grid_pin_5_ ;
wire [0:0] cby_1__1__126_left_grid_pin_6_ ;
wire [0:0] cby_1__1__126_left_grid_pin_7_ ;
wire [0:0] cby_1__1__126_left_grid_pin_8_ ;
wire [0:0] cby_1__1__126_left_grid_pin_9_ ;
wire [0:0] cby_1__1__126_right_grid_pin_52_ ;
wire [0:0] cby_1__1__127_ccff_tail ;
wire [0:19] cby_1__1__127_chany_bottom_out ;
wire [0:19] cby_1__1__127_chany_top_out ;
wire [0:0] cby_1__1__127_left_grid_pin_0_ ;
wire [0:0] cby_1__1__127_left_grid_pin_10_ ;
wire [0:0] cby_1__1__127_left_grid_pin_11_ ;
wire [0:0] cby_1__1__127_left_grid_pin_12_ ;
wire [0:0] cby_1__1__127_left_grid_pin_13_ ;
wire [0:0] cby_1__1__127_left_grid_pin_14_ ;
wire [0:0] cby_1__1__127_left_grid_pin_15_ ;
wire [0:0] cby_1__1__127_left_grid_pin_1_ ;
wire [0:0] cby_1__1__127_left_grid_pin_2_ ;
wire [0:0] cby_1__1__127_left_grid_pin_3_ ;
wire [0:0] cby_1__1__127_left_grid_pin_4_ ;
wire [0:0] cby_1__1__127_left_grid_pin_5_ ;
wire [0:0] cby_1__1__127_left_grid_pin_6_ ;
wire [0:0] cby_1__1__127_left_grid_pin_7_ ;
wire [0:0] cby_1__1__127_left_grid_pin_8_ ;
wire [0:0] cby_1__1__127_left_grid_pin_9_ ;
wire [0:0] cby_1__1__127_right_grid_pin_52_ ;
wire [0:0] cby_1__1__128_ccff_tail ;
wire [0:19] cby_1__1__128_chany_bottom_out ;
wire [0:19] cby_1__1__128_chany_top_out ;
wire [0:0] cby_1__1__128_left_grid_pin_0_ ;
wire [0:0] cby_1__1__128_left_grid_pin_10_ ;
wire [0:0] cby_1__1__128_left_grid_pin_11_ ;
wire [0:0] cby_1__1__128_left_grid_pin_12_ ;
wire [0:0] cby_1__1__128_left_grid_pin_13_ ;
wire [0:0] cby_1__1__128_left_grid_pin_14_ ;
wire [0:0] cby_1__1__128_left_grid_pin_15_ ;
wire [0:0] cby_1__1__128_left_grid_pin_1_ ;
wire [0:0] cby_1__1__128_left_grid_pin_2_ ;
wire [0:0] cby_1__1__128_left_grid_pin_3_ ;
wire [0:0] cby_1__1__128_left_grid_pin_4_ ;
wire [0:0] cby_1__1__128_left_grid_pin_5_ ;
wire [0:0] cby_1__1__128_left_grid_pin_6_ ;
wire [0:0] cby_1__1__128_left_grid_pin_7_ ;
wire [0:0] cby_1__1__128_left_grid_pin_8_ ;
wire [0:0] cby_1__1__128_left_grid_pin_9_ ;
wire [0:0] cby_1__1__128_right_grid_pin_52_ ;
wire [0:0] cby_1__1__129_ccff_tail ;
wire [0:19] cby_1__1__129_chany_bottom_out ;
wire [0:19] cby_1__1__129_chany_top_out ;
wire [0:0] cby_1__1__129_left_grid_pin_0_ ;
wire [0:0] cby_1__1__129_left_grid_pin_10_ ;
wire [0:0] cby_1__1__129_left_grid_pin_11_ ;
wire [0:0] cby_1__1__129_left_grid_pin_12_ ;
wire [0:0] cby_1__1__129_left_grid_pin_13_ ;
wire [0:0] cby_1__1__129_left_grid_pin_14_ ;
wire [0:0] cby_1__1__129_left_grid_pin_15_ ;
wire [0:0] cby_1__1__129_left_grid_pin_1_ ;
wire [0:0] cby_1__1__129_left_grid_pin_2_ ;
wire [0:0] cby_1__1__129_left_grid_pin_3_ ;
wire [0:0] cby_1__1__129_left_grid_pin_4_ ;
wire [0:0] cby_1__1__129_left_grid_pin_5_ ;
wire [0:0] cby_1__1__129_left_grid_pin_6_ ;
wire [0:0] cby_1__1__129_left_grid_pin_7_ ;
wire [0:0] cby_1__1__129_left_grid_pin_8_ ;
wire [0:0] cby_1__1__129_left_grid_pin_9_ ;
wire [0:0] cby_1__1__129_right_grid_pin_52_ ;
wire [0:0] cby_1__1__12_ccff_tail ;
wire [0:19] cby_1__1__12_chany_bottom_out ;
wire [0:19] cby_1__1__12_chany_top_out ;
wire [0:0] cby_1__1__12_left_grid_pin_0_ ;
wire [0:0] cby_1__1__12_left_grid_pin_10_ ;
wire [0:0] cby_1__1__12_left_grid_pin_11_ ;
wire [0:0] cby_1__1__12_left_grid_pin_12_ ;
wire [0:0] cby_1__1__12_left_grid_pin_13_ ;
wire [0:0] cby_1__1__12_left_grid_pin_14_ ;
wire [0:0] cby_1__1__12_left_grid_pin_15_ ;
wire [0:0] cby_1__1__12_left_grid_pin_1_ ;
wire [0:0] cby_1__1__12_left_grid_pin_2_ ;
wire [0:0] cby_1__1__12_left_grid_pin_3_ ;
wire [0:0] cby_1__1__12_left_grid_pin_4_ ;
wire [0:0] cby_1__1__12_left_grid_pin_5_ ;
wire [0:0] cby_1__1__12_left_grid_pin_6_ ;
wire [0:0] cby_1__1__12_left_grid_pin_7_ ;
wire [0:0] cby_1__1__12_left_grid_pin_8_ ;
wire [0:0] cby_1__1__12_left_grid_pin_9_ ;
wire [0:0] cby_1__1__12_right_grid_pin_52_ ;
wire [0:0] cby_1__1__130_ccff_tail ;
wire [0:19] cby_1__1__130_chany_bottom_out ;
wire [0:19] cby_1__1__130_chany_top_out ;
wire [0:0] cby_1__1__130_left_grid_pin_0_ ;
wire [0:0] cby_1__1__130_left_grid_pin_10_ ;
wire [0:0] cby_1__1__130_left_grid_pin_11_ ;
wire [0:0] cby_1__1__130_left_grid_pin_12_ ;
wire [0:0] cby_1__1__130_left_grid_pin_13_ ;
wire [0:0] cby_1__1__130_left_grid_pin_14_ ;
wire [0:0] cby_1__1__130_left_grid_pin_15_ ;
wire [0:0] cby_1__1__130_left_grid_pin_1_ ;
wire [0:0] cby_1__1__130_left_grid_pin_2_ ;
wire [0:0] cby_1__1__130_left_grid_pin_3_ ;
wire [0:0] cby_1__1__130_left_grid_pin_4_ ;
wire [0:0] cby_1__1__130_left_grid_pin_5_ ;
wire [0:0] cby_1__1__130_left_grid_pin_6_ ;
wire [0:0] cby_1__1__130_left_grid_pin_7_ ;
wire [0:0] cby_1__1__130_left_grid_pin_8_ ;
wire [0:0] cby_1__1__130_left_grid_pin_9_ ;
wire [0:0] cby_1__1__130_right_grid_pin_52_ ;
wire [0:0] cby_1__1__131_ccff_tail ;
wire [0:19] cby_1__1__131_chany_bottom_out ;
wire [0:19] cby_1__1__131_chany_top_out ;
wire [0:0] cby_1__1__131_left_grid_pin_0_ ;
wire [0:0] cby_1__1__131_left_grid_pin_10_ ;
wire [0:0] cby_1__1__131_left_grid_pin_11_ ;
wire [0:0] cby_1__1__131_left_grid_pin_12_ ;
wire [0:0] cby_1__1__131_left_grid_pin_13_ ;
wire [0:0] cby_1__1__131_left_grid_pin_14_ ;
wire [0:0] cby_1__1__131_left_grid_pin_15_ ;
wire [0:0] cby_1__1__131_left_grid_pin_1_ ;
wire [0:0] cby_1__1__131_left_grid_pin_2_ ;
wire [0:0] cby_1__1__131_left_grid_pin_3_ ;
wire [0:0] cby_1__1__131_left_grid_pin_4_ ;
wire [0:0] cby_1__1__131_left_grid_pin_5_ ;
wire [0:0] cby_1__1__131_left_grid_pin_6_ ;
wire [0:0] cby_1__1__131_left_grid_pin_7_ ;
wire [0:0] cby_1__1__131_left_grid_pin_8_ ;
wire [0:0] cby_1__1__131_left_grid_pin_9_ ;
wire [0:0] cby_1__1__131_right_grid_pin_52_ ;
wire [0:0] cby_1__1__132_ccff_tail ;
wire [0:19] cby_1__1__132_chany_bottom_out ;
wire [0:19] cby_1__1__132_chany_top_out ;
wire [0:0] cby_1__1__132_left_grid_pin_0_ ;
wire [0:0] cby_1__1__132_left_grid_pin_10_ ;
wire [0:0] cby_1__1__132_left_grid_pin_11_ ;
wire [0:0] cby_1__1__132_left_grid_pin_12_ ;
wire [0:0] cby_1__1__132_left_grid_pin_13_ ;
wire [0:0] cby_1__1__132_left_grid_pin_14_ ;
wire [0:0] cby_1__1__132_left_grid_pin_15_ ;
wire [0:0] cby_1__1__132_left_grid_pin_1_ ;
wire [0:0] cby_1__1__132_left_grid_pin_2_ ;
wire [0:0] cby_1__1__132_left_grid_pin_3_ ;
wire [0:0] cby_1__1__132_left_grid_pin_4_ ;
wire [0:0] cby_1__1__132_left_grid_pin_5_ ;
wire [0:0] cby_1__1__132_left_grid_pin_6_ ;
wire [0:0] cby_1__1__132_left_grid_pin_7_ ;
wire [0:0] cby_1__1__132_left_grid_pin_8_ ;
wire [0:0] cby_1__1__132_left_grid_pin_9_ ;
wire [0:0] cby_1__1__132_right_grid_pin_52_ ;
wire [0:0] cby_1__1__133_ccff_tail ;
wire [0:19] cby_1__1__133_chany_bottom_out ;
wire [0:19] cby_1__1__133_chany_top_out ;
wire [0:0] cby_1__1__133_left_grid_pin_0_ ;
wire [0:0] cby_1__1__133_left_grid_pin_10_ ;
wire [0:0] cby_1__1__133_left_grid_pin_11_ ;
wire [0:0] cby_1__1__133_left_grid_pin_12_ ;
wire [0:0] cby_1__1__133_left_grid_pin_13_ ;
wire [0:0] cby_1__1__133_left_grid_pin_14_ ;
wire [0:0] cby_1__1__133_left_grid_pin_15_ ;
wire [0:0] cby_1__1__133_left_grid_pin_1_ ;
wire [0:0] cby_1__1__133_left_grid_pin_2_ ;
wire [0:0] cby_1__1__133_left_grid_pin_3_ ;
wire [0:0] cby_1__1__133_left_grid_pin_4_ ;
wire [0:0] cby_1__1__133_left_grid_pin_5_ ;
wire [0:0] cby_1__1__133_left_grid_pin_6_ ;
wire [0:0] cby_1__1__133_left_grid_pin_7_ ;
wire [0:0] cby_1__1__133_left_grid_pin_8_ ;
wire [0:0] cby_1__1__133_left_grid_pin_9_ ;
wire [0:0] cby_1__1__133_right_grid_pin_52_ ;
wire [0:0] cby_1__1__134_ccff_tail ;
wire [0:19] cby_1__1__134_chany_bottom_out ;
wire [0:19] cby_1__1__134_chany_top_out ;
wire [0:0] cby_1__1__134_left_grid_pin_0_ ;
wire [0:0] cby_1__1__134_left_grid_pin_10_ ;
wire [0:0] cby_1__1__134_left_grid_pin_11_ ;
wire [0:0] cby_1__1__134_left_grid_pin_12_ ;
wire [0:0] cby_1__1__134_left_grid_pin_13_ ;
wire [0:0] cby_1__1__134_left_grid_pin_14_ ;
wire [0:0] cby_1__1__134_left_grid_pin_15_ ;
wire [0:0] cby_1__1__134_left_grid_pin_1_ ;
wire [0:0] cby_1__1__134_left_grid_pin_2_ ;
wire [0:0] cby_1__1__134_left_grid_pin_3_ ;
wire [0:0] cby_1__1__134_left_grid_pin_4_ ;
wire [0:0] cby_1__1__134_left_grid_pin_5_ ;
wire [0:0] cby_1__1__134_left_grid_pin_6_ ;
wire [0:0] cby_1__1__134_left_grid_pin_7_ ;
wire [0:0] cby_1__1__134_left_grid_pin_8_ ;
wire [0:0] cby_1__1__134_left_grid_pin_9_ ;
wire [0:0] cby_1__1__134_right_grid_pin_52_ ;
wire [0:0] cby_1__1__135_ccff_tail ;
wire [0:19] cby_1__1__135_chany_bottom_out ;
wire [0:19] cby_1__1__135_chany_top_out ;
wire [0:0] cby_1__1__135_left_grid_pin_0_ ;
wire [0:0] cby_1__1__135_left_grid_pin_10_ ;
wire [0:0] cby_1__1__135_left_grid_pin_11_ ;
wire [0:0] cby_1__1__135_left_grid_pin_12_ ;
wire [0:0] cby_1__1__135_left_grid_pin_13_ ;
wire [0:0] cby_1__1__135_left_grid_pin_14_ ;
wire [0:0] cby_1__1__135_left_grid_pin_15_ ;
wire [0:0] cby_1__1__135_left_grid_pin_1_ ;
wire [0:0] cby_1__1__135_left_grid_pin_2_ ;
wire [0:0] cby_1__1__135_left_grid_pin_3_ ;
wire [0:0] cby_1__1__135_left_grid_pin_4_ ;
wire [0:0] cby_1__1__135_left_grid_pin_5_ ;
wire [0:0] cby_1__1__135_left_grid_pin_6_ ;
wire [0:0] cby_1__1__135_left_grid_pin_7_ ;
wire [0:0] cby_1__1__135_left_grid_pin_8_ ;
wire [0:0] cby_1__1__135_left_grid_pin_9_ ;
wire [0:0] cby_1__1__135_right_grid_pin_52_ ;
wire [0:0] cby_1__1__136_ccff_tail ;
wire [0:19] cby_1__1__136_chany_bottom_out ;
wire [0:19] cby_1__1__136_chany_top_out ;
wire [0:0] cby_1__1__136_left_grid_pin_0_ ;
wire [0:0] cby_1__1__136_left_grid_pin_10_ ;
wire [0:0] cby_1__1__136_left_grid_pin_11_ ;
wire [0:0] cby_1__1__136_left_grid_pin_12_ ;
wire [0:0] cby_1__1__136_left_grid_pin_13_ ;
wire [0:0] cby_1__1__136_left_grid_pin_14_ ;
wire [0:0] cby_1__1__136_left_grid_pin_15_ ;
wire [0:0] cby_1__1__136_left_grid_pin_1_ ;
wire [0:0] cby_1__1__136_left_grid_pin_2_ ;
wire [0:0] cby_1__1__136_left_grid_pin_3_ ;
wire [0:0] cby_1__1__136_left_grid_pin_4_ ;
wire [0:0] cby_1__1__136_left_grid_pin_5_ ;
wire [0:0] cby_1__1__136_left_grid_pin_6_ ;
wire [0:0] cby_1__1__136_left_grid_pin_7_ ;
wire [0:0] cby_1__1__136_left_grid_pin_8_ ;
wire [0:0] cby_1__1__136_left_grid_pin_9_ ;
wire [0:0] cby_1__1__136_right_grid_pin_52_ ;
wire [0:0] cby_1__1__137_ccff_tail ;
wire [0:19] cby_1__1__137_chany_bottom_out ;
wire [0:19] cby_1__1__137_chany_top_out ;
wire [0:0] cby_1__1__137_left_grid_pin_0_ ;
wire [0:0] cby_1__1__137_left_grid_pin_10_ ;
wire [0:0] cby_1__1__137_left_grid_pin_11_ ;
wire [0:0] cby_1__1__137_left_grid_pin_12_ ;
wire [0:0] cby_1__1__137_left_grid_pin_13_ ;
wire [0:0] cby_1__1__137_left_grid_pin_14_ ;
wire [0:0] cby_1__1__137_left_grid_pin_15_ ;
wire [0:0] cby_1__1__137_left_grid_pin_1_ ;
wire [0:0] cby_1__1__137_left_grid_pin_2_ ;
wire [0:0] cby_1__1__137_left_grid_pin_3_ ;
wire [0:0] cby_1__1__137_left_grid_pin_4_ ;
wire [0:0] cby_1__1__137_left_grid_pin_5_ ;
wire [0:0] cby_1__1__137_left_grid_pin_6_ ;
wire [0:0] cby_1__1__137_left_grid_pin_7_ ;
wire [0:0] cby_1__1__137_left_grid_pin_8_ ;
wire [0:0] cby_1__1__137_left_grid_pin_9_ ;
wire [0:0] cby_1__1__137_right_grid_pin_52_ ;
wire [0:0] cby_1__1__138_ccff_tail ;
wire [0:19] cby_1__1__138_chany_bottom_out ;
wire [0:19] cby_1__1__138_chany_top_out ;
wire [0:0] cby_1__1__138_left_grid_pin_0_ ;
wire [0:0] cby_1__1__138_left_grid_pin_10_ ;
wire [0:0] cby_1__1__138_left_grid_pin_11_ ;
wire [0:0] cby_1__1__138_left_grid_pin_12_ ;
wire [0:0] cby_1__1__138_left_grid_pin_13_ ;
wire [0:0] cby_1__1__138_left_grid_pin_14_ ;
wire [0:0] cby_1__1__138_left_grid_pin_15_ ;
wire [0:0] cby_1__1__138_left_grid_pin_1_ ;
wire [0:0] cby_1__1__138_left_grid_pin_2_ ;
wire [0:0] cby_1__1__138_left_grid_pin_3_ ;
wire [0:0] cby_1__1__138_left_grid_pin_4_ ;
wire [0:0] cby_1__1__138_left_grid_pin_5_ ;
wire [0:0] cby_1__1__138_left_grid_pin_6_ ;
wire [0:0] cby_1__1__138_left_grid_pin_7_ ;
wire [0:0] cby_1__1__138_left_grid_pin_8_ ;
wire [0:0] cby_1__1__138_left_grid_pin_9_ ;
wire [0:0] cby_1__1__138_right_grid_pin_52_ ;
wire [0:0] cby_1__1__139_ccff_tail ;
wire [0:19] cby_1__1__139_chany_bottom_out ;
wire [0:19] cby_1__1__139_chany_top_out ;
wire [0:0] cby_1__1__139_left_grid_pin_0_ ;
wire [0:0] cby_1__1__139_left_grid_pin_10_ ;
wire [0:0] cby_1__1__139_left_grid_pin_11_ ;
wire [0:0] cby_1__1__139_left_grid_pin_12_ ;
wire [0:0] cby_1__1__139_left_grid_pin_13_ ;
wire [0:0] cby_1__1__139_left_grid_pin_14_ ;
wire [0:0] cby_1__1__139_left_grid_pin_15_ ;
wire [0:0] cby_1__1__139_left_grid_pin_1_ ;
wire [0:0] cby_1__1__139_left_grid_pin_2_ ;
wire [0:0] cby_1__1__139_left_grid_pin_3_ ;
wire [0:0] cby_1__1__139_left_grid_pin_4_ ;
wire [0:0] cby_1__1__139_left_grid_pin_5_ ;
wire [0:0] cby_1__1__139_left_grid_pin_6_ ;
wire [0:0] cby_1__1__139_left_grid_pin_7_ ;
wire [0:0] cby_1__1__139_left_grid_pin_8_ ;
wire [0:0] cby_1__1__139_left_grid_pin_9_ ;
wire [0:0] cby_1__1__139_right_grid_pin_52_ ;
wire [0:0] cby_1__1__13_ccff_tail ;
wire [0:19] cby_1__1__13_chany_bottom_out ;
wire [0:19] cby_1__1__13_chany_top_out ;
wire [0:0] cby_1__1__13_left_grid_pin_0_ ;
wire [0:0] cby_1__1__13_left_grid_pin_10_ ;
wire [0:0] cby_1__1__13_left_grid_pin_11_ ;
wire [0:0] cby_1__1__13_left_grid_pin_12_ ;
wire [0:0] cby_1__1__13_left_grid_pin_13_ ;
wire [0:0] cby_1__1__13_left_grid_pin_14_ ;
wire [0:0] cby_1__1__13_left_grid_pin_15_ ;
wire [0:0] cby_1__1__13_left_grid_pin_1_ ;
wire [0:0] cby_1__1__13_left_grid_pin_2_ ;
wire [0:0] cby_1__1__13_left_grid_pin_3_ ;
wire [0:0] cby_1__1__13_left_grid_pin_4_ ;
wire [0:0] cby_1__1__13_left_grid_pin_5_ ;
wire [0:0] cby_1__1__13_left_grid_pin_6_ ;
wire [0:0] cby_1__1__13_left_grid_pin_7_ ;
wire [0:0] cby_1__1__13_left_grid_pin_8_ ;
wire [0:0] cby_1__1__13_left_grid_pin_9_ ;
wire [0:0] cby_1__1__13_right_grid_pin_52_ ;
wire [0:0] cby_1__1__140_ccff_tail ;
wire [0:19] cby_1__1__140_chany_bottom_out ;
wire [0:19] cby_1__1__140_chany_top_out ;
wire [0:0] cby_1__1__140_left_grid_pin_0_ ;
wire [0:0] cby_1__1__140_left_grid_pin_10_ ;
wire [0:0] cby_1__1__140_left_grid_pin_11_ ;
wire [0:0] cby_1__1__140_left_grid_pin_12_ ;
wire [0:0] cby_1__1__140_left_grid_pin_13_ ;
wire [0:0] cby_1__1__140_left_grid_pin_14_ ;
wire [0:0] cby_1__1__140_left_grid_pin_15_ ;
wire [0:0] cby_1__1__140_left_grid_pin_1_ ;
wire [0:0] cby_1__1__140_left_grid_pin_2_ ;
wire [0:0] cby_1__1__140_left_grid_pin_3_ ;
wire [0:0] cby_1__1__140_left_grid_pin_4_ ;
wire [0:0] cby_1__1__140_left_grid_pin_5_ ;
wire [0:0] cby_1__1__140_left_grid_pin_6_ ;
wire [0:0] cby_1__1__140_left_grid_pin_7_ ;
wire [0:0] cby_1__1__140_left_grid_pin_8_ ;
wire [0:0] cby_1__1__140_left_grid_pin_9_ ;
wire [0:0] cby_1__1__140_right_grid_pin_52_ ;
wire [0:0] cby_1__1__141_ccff_tail ;
wire [0:19] cby_1__1__141_chany_bottom_out ;
wire [0:19] cby_1__1__141_chany_top_out ;
wire [0:0] cby_1__1__141_left_grid_pin_0_ ;
wire [0:0] cby_1__1__141_left_grid_pin_10_ ;
wire [0:0] cby_1__1__141_left_grid_pin_11_ ;
wire [0:0] cby_1__1__141_left_grid_pin_12_ ;
wire [0:0] cby_1__1__141_left_grid_pin_13_ ;
wire [0:0] cby_1__1__141_left_grid_pin_14_ ;
wire [0:0] cby_1__1__141_left_grid_pin_15_ ;
wire [0:0] cby_1__1__141_left_grid_pin_1_ ;
wire [0:0] cby_1__1__141_left_grid_pin_2_ ;
wire [0:0] cby_1__1__141_left_grid_pin_3_ ;
wire [0:0] cby_1__1__141_left_grid_pin_4_ ;
wire [0:0] cby_1__1__141_left_grid_pin_5_ ;
wire [0:0] cby_1__1__141_left_grid_pin_6_ ;
wire [0:0] cby_1__1__141_left_grid_pin_7_ ;
wire [0:0] cby_1__1__141_left_grid_pin_8_ ;
wire [0:0] cby_1__1__141_left_grid_pin_9_ ;
wire [0:0] cby_1__1__141_right_grid_pin_52_ ;
wire [0:0] cby_1__1__142_ccff_tail ;
wire [0:19] cby_1__1__142_chany_bottom_out ;
wire [0:19] cby_1__1__142_chany_top_out ;
wire [0:0] cby_1__1__142_left_grid_pin_0_ ;
wire [0:0] cby_1__1__142_left_grid_pin_10_ ;
wire [0:0] cby_1__1__142_left_grid_pin_11_ ;
wire [0:0] cby_1__1__142_left_grid_pin_12_ ;
wire [0:0] cby_1__1__142_left_grid_pin_13_ ;
wire [0:0] cby_1__1__142_left_grid_pin_14_ ;
wire [0:0] cby_1__1__142_left_grid_pin_15_ ;
wire [0:0] cby_1__1__142_left_grid_pin_1_ ;
wire [0:0] cby_1__1__142_left_grid_pin_2_ ;
wire [0:0] cby_1__1__142_left_grid_pin_3_ ;
wire [0:0] cby_1__1__142_left_grid_pin_4_ ;
wire [0:0] cby_1__1__142_left_grid_pin_5_ ;
wire [0:0] cby_1__1__142_left_grid_pin_6_ ;
wire [0:0] cby_1__1__142_left_grid_pin_7_ ;
wire [0:0] cby_1__1__142_left_grid_pin_8_ ;
wire [0:0] cby_1__1__142_left_grid_pin_9_ ;
wire [0:0] cby_1__1__142_right_grid_pin_52_ ;
wire [0:0] cby_1__1__143_ccff_tail ;
wire [0:19] cby_1__1__143_chany_bottom_out ;
wire [0:19] cby_1__1__143_chany_top_out ;
wire [0:0] cby_1__1__143_left_grid_pin_0_ ;
wire [0:0] cby_1__1__143_left_grid_pin_10_ ;
wire [0:0] cby_1__1__143_left_grid_pin_11_ ;
wire [0:0] cby_1__1__143_left_grid_pin_12_ ;
wire [0:0] cby_1__1__143_left_grid_pin_13_ ;
wire [0:0] cby_1__1__143_left_grid_pin_14_ ;
wire [0:0] cby_1__1__143_left_grid_pin_15_ ;
wire [0:0] cby_1__1__143_left_grid_pin_1_ ;
wire [0:0] cby_1__1__143_left_grid_pin_2_ ;
wire [0:0] cby_1__1__143_left_grid_pin_3_ ;
wire [0:0] cby_1__1__143_left_grid_pin_4_ ;
wire [0:0] cby_1__1__143_left_grid_pin_5_ ;
wire [0:0] cby_1__1__143_left_grid_pin_6_ ;
wire [0:0] cby_1__1__143_left_grid_pin_7_ ;
wire [0:0] cby_1__1__143_left_grid_pin_8_ ;
wire [0:0] cby_1__1__143_left_grid_pin_9_ ;
wire [0:0] cby_1__1__143_right_grid_pin_52_ ;
wire [0:0] cby_1__1__14_ccff_tail ;
wire [0:19] cby_1__1__14_chany_bottom_out ;
wire [0:19] cby_1__1__14_chany_top_out ;
wire [0:0] cby_1__1__14_left_grid_pin_0_ ;
wire [0:0] cby_1__1__14_left_grid_pin_10_ ;
wire [0:0] cby_1__1__14_left_grid_pin_11_ ;
wire [0:0] cby_1__1__14_left_grid_pin_12_ ;
wire [0:0] cby_1__1__14_left_grid_pin_13_ ;
wire [0:0] cby_1__1__14_left_grid_pin_14_ ;
wire [0:0] cby_1__1__14_left_grid_pin_15_ ;
wire [0:0] cby_1__1__14_left_grid_pin_1_ ;
wire [0:0] cby_1__1__14_left_grid_pin_2_ ;
wire [0:0] cby_1__1__14_left_grid_pin_3_ ;
wire [0:0] cby_1__1__14_left_grid_pin_4_ ;
wire [0:0] cby_1__1__14_left_grid_pin_5_ ;
wire [0:0] cby_1__1__14_left_grid_pin_6_ ;
wire [0:0] cby_1__1__14_left_grid_pin_7_ ;
wire [0:0] cby_1__1__14_left_grid_pin_8_ ;
wire [0:0] cby_1__1__14_left_grid_pin_9_ ;
wire [0:0] cby_1__1__14_right_grid_pin_52_ ;
wire [0:0] cby_1__1__15_ccff_tail ;
wire [0:19] cby_1__1__15_chany_bottom_out ;
wire [0:19] cby_1__1__15_chany_top_out ;
wire [0:0] cby_1__1__15_left_grid_pin_0_ ;
wire [0:0] cby_1__1__15_left_grid_pin_10_ ;
wire [0:0] cby_1__1__15_left_grid_pin_11_ ;
wire [0:0] cby_1__1__15_left_grid_pin_12_ ;
wire [0:0] cby_1__1__15_left_grid_pin_13_ ;
wire [0:0] cby_1__1__15_left_grid_pin_14_ ;
wire [0:0] cby_1__1__15_left_grid_pin_15_ ;
wire [0:0] cby_1__1__15_left_grid_pin_1_ ;
wire [0:0] cby_1__1__15_left_grid_pin_2_ ;
wire [0:0] cby_1__1__15_left_grid_pin_3_ ;
wire [0:0] cby_1__1__15_left_grid_pin_4_ ;
wire [0:0] cby_1__1__15_left_grid_pin_5_ ;
wire [0:0] cby_1__1__15_left_grid_pin_6_ ;
wire [0:0] cby_1__1__15_left_grid_pin_7_ ;
wire [0:0] cby_1__1__15_left_grid_pin_8_ ;
wire [0:0] cby_1__1__15_left_grid_pin_9_ ;
wire [0:0] cby_1__1__15_right_grid_pin_52_ ;
wire [0:0] cby_1__1__16_ccff_tail ;
wire [0:19] cby_1__1__16_chany_bottom_out ;
wire [0:19] cby_1__1__16_chany_top_out ;
wire [0:0] cby_1__1__16_left_grid_pin_0_ ;
wire [0:0] cby_1__1__16_left_grid_pin_10_ ;
wire [0:0] cby_1__1__16_left_grid_pin_11_ ;
wire [0:0] cby_1__1__16_left_grid_pin_12_ ;
wire [0:0] cby_1__1__16_left_grid_pin_13_ ;
wire [0:0] cby_1__1__16_left_grid_pin_14_ ;
wire [0:0] cby_1__1__16_left_grid_pin_15_ ;
wire [0:0] cby_1__1__16_left_grid_pin_1_ ;
wire [0:0] cby_1__1__16_left_grid_pin_2_ ;
wire [0:0] cby_1__1__16_left_grid_pin_3_ ;
wire [0:0] cby_1__1__16_left_grid_pin_4_ ;
wire [0:0] cby_1__1__16_left_grid_pin_5_ ;
wire [0:0] cby_1__1__16_left_grid_pin_6_ ;
wire [0:0] cby_1__1__16_left_grid_pin_7_ ;
wire [0:0] cby_1__1__16_left_grid_pin_8_ ;
wire [0:0] cby_1__1__16_left_grid_pin_9_ ;
wire [0:0] cby_1__1__16_right_grid_pin_52_ ;
wire [0:0] cby_1__1__17_ccff_tail ;
wire [0:19] cby_1__1__17_chany_bottom_out ;
wire [0:19] cby_1__1__17_chany_top_out ;
wire [0:0] cby_1__1__17_left_grid_pin_0_ ;
wire [0:0] cby_1__1__17_left_grid_pin_10_ ;
wire [0:0] cby_1__1__17_left_grid_pin_11_ ;
wire [0:0] cby_1__1__17_left_grid_pin_12_ ;
wire [0:0] cby_1__1__17_left_grid_pin_13_ ;
wire [0:0] cby_1__1__17_left_grid_pin_14_ ;
wire [0:0] cby_1__1__17_left_grid_pin_15_ ;
wire [0:0] cby_1__1__17_left_grid_pin_1_ ;
wire [0:0] cby_1__1__17_left_grid_pin_2_ ;
wire [0:0] cby_1__1__17_left_grid_pin_3_ ;
wire [0:0] cby_1__1__17_left_grid_pin_4_ ;
wire [0:0] cby_1__1__17_left_grid_pin_5_ ;
wire [0:0] cby_1__1__17_left_grid_pin_6_ ;
wire [0:0] cby_1__1__17_left_grid_pin_7_ ;
wire [0:0] cby_1__1__17_left_grid_pin_8_ ;
wire [0:0] cby_1__1__17_left_grid_pin_9_ ;
wire [0:0] cby_1__1__17_right_grid_pin_52_ ;
wire [0:0] cby_1__1__18_ccff_tail ;
wire [0:19] cby_1__1__18_chany_bottom_out ;
wire [0:19] cby_1__1__18_chany_top_out ;
wire [0:0] cby_1__1__18_left_grid_pin_0_ ;
wire [0:0] cby_1__1__18_left_grid_pin_10_ ;
wire [0:0] cby_1__1__18_left_grid_pin_11_ ;
wire [0:0] cby_1__1__18_left_grid_pin_12_ ;
wire [0:0] cby_1__1__18_left_grid_pin_13_ ;
wire [0:0] cby_1__1__18_left_grid_pin_14_ ;
wire [0:0] cby_1__1__18_left_grid_pin_15_ ;
wire [0:0] cby_1__1__18_left_grid_pin_1_ ;
wire [0:0] cby_1__1__18_left_grid_pin_2_ ;
wire [0:0] cby_1__1__18_left_grid_pin_3_ ;
wire [0:0] cby_1__1__18_left_grid_pin_4_ ;
wire [0:0] cby_1__1__18_left_grid_pin_5_ ;
wire [0:0] cby_1__1__18_left_grid_pin_6_ ;
wire [0:0] cby_1__1__18_left_grid_pin_7_ ;
wire [0:0] cby_1__1__18_left_grid_pin_8_ ;
wire [0:0] cby_1__1__18_left_grid_pin_9_ ;
wire [0:0] cby_1__1__18_right_grid_pin_52_ ;
wire [0:0] cby_1__1__19_ccff_tail ;
wire [0:19] cby_1__1__19_chany_bottom_out ;
wire [0:19] cby_1__1__19_chany_top_out ;
wire [0:0] cby_1__1__19_left_grid_pin_0_ ;
wire [0:0] cby_1__1__19_left_grid_pin_10_ ;
wire [0:0] cby_1__1__19_left_grid_pin_11_ ;
wire [0:0] cby_1__1__19_left_grid_pin_12_ ;
wire [0:0] cby_1__1__19_left_grid_pin_13_ ;
wire [0:0] cby_1__1__19_left_grid_pin_14_ ;
wire [0:0] cby_1__1__19_left_grid_pin_15_ ;
wire [0:0] cby_1__1__19_left_grid_pin_1_ ;
wire [0:0] cby_1__1__19_left_grid_pin_2_ ;
wire [0:0] cby_1__1__19_left_grid_pin_3_ ;
wire [0:0] cby_1__1__19_left_grid_pin_4_ ;
wire [0:0] cby_1__1__19_left_grid_pin_5_ ;
wire [0:0] cby_1__1__19_left_grid_pin_6_ ;
wire [0:0] cby_1__1__19_left_grid_pin_7_ ;
wire [0:0] cby_1__1__19_left_grid_pin_8_ ;
wire [0:0] cby_1__1__19_left_grid_pin_9_ ;
wire [0:0] cby_1__1__19_right_grid_pin_52_ ;
wire [0:0] cby_1__1__1_ccff_tail ;
wire [0:19] cby_1__1__1_chany_bottom_out ;
wire [0:19] cby_1__1__1_chany_top_out ;
wire [0:0] cby_1__1__1_left_grid_pin_0_ ;
wire [0:0] cby_1__1__1_left_grid_pin_10_ ;
wire [0:0] cby_1__1__1_left_grid_pin_11_ ;
wire [0:0] cby_1__1__1_left_grid_pin_12_ ;
wire [0:0] cby_1__1__1_left_grid_pin_13_ ;
wire [0:0] cby_1__1__1_left_grid_pin_14_ ;
wire [0:0] cby_1__1__1_left_grid_pin_15_ ;
wire [0:0] cby_1__1__1_left_grid_pin_1_ ;
wire [0:0] cby_1__1__1_left_grid_pin_2_ ;
wire [0:0] cby_1__1__1_left_grid_pin_3_ ;
wire [0:0] cby_1__1__1_left_grid_pin_4_ ;
wire [0:0] cby_1__1__1_left_grid_pin_5_ ;
wire [0:0] cby_1__1__1_left_grid_pin_6_ ;
wire [0:0] cby_1__1__1_left_grid_pin_7_ ;
wire [0:0] cby_1__1__1_left_grid_pin_8_ ;
wire [0:0] cby_1__1__1_left_grid_pin_9_ ;
wire [0:0] cby_1__1__1_right_grid_pin_52_ ;
wire [0:0] cby_1__1__20_ccff_tail ;
wire [0:19] cby_1__1__20_chany_bottom_out ;
wire [0:19] cby_1__1__20_chany_top_out ;
wire [0:0] cby_1__1__20_left_grid_pin_0_ ;
wire [0:0] cby_1__1__20_left_grid_pin_10_ ;
wire [0:0] cby_1__1__20_left_grid_pin_11_ ;
wire [0:0] cby_1__1__20_left_grid_pin_12_ ;
wire [0:0] cby_1__1__20_left_grid_pin_13_ ;
wire [0:0] cby_1__1__20_left_grid_pin_14_ ;
wire [0:0] cby_1__1__20_left_grid_pin_15_ ;
wire [0:0] cby_1__1__20_left_grid_pin_1_ ;
wire [0:0] cby_1__1__20_left_grid_pin_2_ ;
wire [0:0] cby_1__1__20_left_grid_pin_3_ ;
wire [0:0] cby_1__1__20_left_grid_pin_4_ ;
wire [0:0] cby_1__1__20_left_grid_pin_5_ ;
wire [0:0] cby_1__1__20_left_grid_pin_6_ ;
wire [0:0] cby_1__1__20_left_grid_pin_7_ ;
wire [0:0] cby_1__1__20_left_grid_pin_8_ ;
wire [0:0] cby_1__1__20_left_grid_pin_9_ ;
wire [0:0] cby_1__1__20_right_grid_pin_52_ ;
wire [0:0] cby_1__1__21_ccff_tail ;
wire [0:19] cby_1__1__21_chany_bottom_out ;
wire [0:19] cby_1__1__21_chany_top_out ;
wire [0:0] cby_1__1__21_left_grid_pin_0_ ;
wire [0:0] cby_1__1__21_left_grid_pin_10_ ;
wire [0:0] cby_1__1__21_left_grid_pin_11_ ;
wire [0:0] cby_1__1__21_left_grid_pin_12_ ;
wire [0:0] cby_1__1__21_left_grid_pin_13_ ;
wire [0:0] cby_1__1__21_left_grid_pin_14_ ;
wire [0:0] cby_1__1__21_left_grid_pin_15_ ;
wire [0:0] cby_1__1__21_left_grid_pin_1_ ;
wire [0:0] cby_1__1__21_left_grid_pin_2_ ;
wire [0:0] cby_1__1__21_left_grid_pin_3_ ;
wire [0:0] cby_1__1__21_left_grid_pin_4_ ;
wire [0:0] cby_1__1__21_left_grid_pin_5_ ;
wire [0:0] cby_1__1__21_left_grid_pin_6_ ;
wire [0:0] cby_1__1__21_left_grid_pin_7_ ;
wire [0:0] cby_1__1__21_left_grid_pin_8_ ;
wire [0:0] cby_1__1__21_left_grid_pin_9_ ;
wire [0:0] cby_1__1__21_right_grid_pin_52_ ;
wire [0:0] cby_1__1__22_ccff_tail ;
wire [0:19] cby_1__1__22_chany_bottom_out ;
wire [0:19] cby_1__1__22_chany_top_out ;
wire [0:0] cby_1__1__22_left_grid_pin_0_ ;
wire [0:0] cby_1__1__22_left_grid_pin_10_ ;
wire [0:0] cby_1__1__22_left_grid_pin_11_ ;
wire [0:0] cby_1__1__22_left_grid_pin_12_ ;
wire [0:0] cby_1__1__22_left_grid_pin_13_ ;
wire [0:0] cby_1__1__22_left_grid_pin_14_ ;
wire [0:0] cby_1__1__22_left_grid_pin_15_ ;
wire [0:0] cby_1__1__22_left_grid_pin_1_ ;
wire [0:0] cby_1__1__22_left_grid_pin_2_ ;
wire [0:0] cby_1__1__22_left_grid_pin_3_ ;
wire [0:0] cby_1__1__22_left_grid_pin_4_ ;
wire [0:0] cby_1__1__22_left_grid_pin_5_ ;
wire [0:0] cby_1__1__22_left_grid_pin_6_ ;
wire [0:0] cby_1__1__22_left_grid_pin_7_ ;
wire [0:0] cby_1__1__22_left_grid_pin_8_ ;
wire [0:0] cby_1__1__22_left_grid_pin_9_ ;
wire [0:0] cby_1__1__22_right_grid_pin_52_ ;
wire [0:0] cby_1__1__23_ccff_tail ;
wire [0:19] cby_1__1__23_chany_bottom_out ;
wire [0:19] cby_1__1__23_chany_top_out ;
wire [0:0] cby_1__1__23_left_grid_pin_0_ ;
wire [0:0] cby_1__1__23_left_grid_pin_10_ ;
wire [0:0] cby_1__1__23_left_grid_pin_11_ ;
wire [0:0] cby_1__1__23_left_grid_pin_12_ ;
wire [0:0] cby_1__1__23_left_grid_pin_13_ ;
wire [0:0] cby_1__1__23_left_grid_pin_14_ ;
wire [0:0] cby_1__1__23_left_grid_pin_15_ ;
wire [0:0] cby_1__1__23_left_grid_pin_1_ ;
wire [0:0] cby_1__1__23_left_grid_pin_2_ ;
wire [0:0] cby_1__1__23_left_grid_pin_3_ ;
wire [0:0] cby_1__1__23_left_grid_pin_4_ ;
wire [0:0] cby_1__1__23_left_grid_pin_5_ ;
wire [0:0] cby_1__1__23_left_grid_pin_6_ ;
wire [0:0] cby_1__1__23_left_grid_pin_7_ ;
wire [0:0] cby_1__1__23_left_grid_pin_8_ ;
wire [0:0] cby_1__1__23_left_grid_pin_9_ ;
wire [0:0] cby_1__1__23_right_grid_pin_52_ ;
wire [0:0] cby_1__1__24_ccff_tail ;
wire [0:19] cby_1__1__24_chany_bottom_out ;
wire [0:19] cby_1__1__24_chany_top_out ;
wire [0:0] cby_1__1__24_left_grid_pin_0_ ;
wire [0:0] cby_1__1__24_left_grid_pin_10_ ;
wire [0:0] cby_1__1__24_left_grid_pin_11_ ;
wire [0:0] cby_1__1__24_left_grid_pin_12_ ;
wire [0:0] cby_1__1__24_left_grid_pin_13_ ;
wire [0:0] cby_1__1__24_left_grid_pin_14_ ;
wire [0:0] cby_1__1__24_left_grid_pin_15_ ;
wire [0:0] cby_1__1__24_left_grid_pin_1_ ;
wire [0:0] cby_1__1__24_left_grid_pin_2_ ;
wire [0:0] cby_1__1__24_left_grid_pin_3_ ;
wire [0:0] cby_1__1__24_left_grid_pin_4_ ;
wire [0:0] cby_1__1__24_left_grid_pin_5_ ;
wire [0:0] cby_1__1__24_left_grid_pin_6_ ;
wire [0:0] cby_1__1__24_left_grid_pin_7_ ;
wire [0:0] cby_1__1__24_left_grid_pin_8_ ;
wire [0:0] cby_1__1__24_left_grid_pin_9_ ;
wire [0:0] cby_1__1__24_right_grid_pin_52_ ;
wire [0:0] cby_1__1__25_ccff_tail ;
wire [0:19] cby_1__1__25_chany_bottom_out ;
wire [0:19] cby_1__1__25_chany_top_out ;
wire [0:0] cby_1__1__25_left_grid_pin_0_ ;
wire [0:0] cby_1__1__25_left_grid_pin_10_ ;
wire [0:0] cby_1__1__25_left_grid_pin_11_ ;
wire [0:0] cby_1__1__25_left_grid_pin_12_ ;
wire [0:0] cby_1__1__25_left_grid_pin_13_ ;
wire [0:0] cby_1__1__25_left_grid_pin_14_ ;
wire [0:0] cby_1__1__25_left_grid_pin_15_ ;
wire [0:0] cby_1__1__25_left_grid_pin_1_ ;
wire [0:0] cby_1__1__25_left_grid_pin_2_ ;
wire [0:0] cby_1__1__25_left_grid_pin_3_ ;
wire [0:0] cby_1__1__25_left_grid_pin_4_ ;
wire [0:0] cby_1__1__25_left_grid_pin_5_ ;
wire [0:0] cby_1__1__25_left_grid_pin_6_ ;
wire [0:0] cby_1__1__25_left_grid_pin_7_ ;
wire [0:0] cby_1__1__25_left_grid_pin_8_ ;
wire [0:0] cby_1__1__25_left_grid_pin_9_ ;
wire [0:0] cby_1__1__25_right_grid_pin_52_ ;
wire [0:0] cby_1__1__26_ccff_tail ;
wire [0:19] cby_1__1__26_chany_bottom_out ;
wire [0:19] cby_1__1__26_chany_top_out ;
wire [0:0] cby_1__1__26_left_grid_pin_0_ ;
wire [0:0] cby_1__1__26_left_grid_pin_10_ ;
wire [0:0] cby_1__1__26_left_grid_pin_11_ ;
wire [0:0] cby_1__1__26_left_grid_pin_12_ ;
wire [0:0] cby_1__1__26_left_grid_pin_13_ ;
wire [0:0] cby_1__1__26_left_grid_pin_14_ ;
wire [0:0] cby_1__1__26_left_grid_pin_15_ ;
wire [0:0] cby_1__1__26_left_grid_pin_1_ ;
wire [0:0] cby_1__1__26_left_grid_pin_2_ ;
wire [0:0] cby_1__1__26_left_grid_pin_3_ ;
wire [0:0] cby_1__1__26_left_grid_pin_4_ ;
wire [0:0] cby_1__1__26_left_grid_pin_5_ ;
wire [0:0] cby_1__1__26_left_grid_pin_6_ ;
wire [0:0] cby_1__1__26_left_grid_pin_7_ ;
wire [0:0] cby_1__1__26_left_grid_pin_8_ ;
wire [0:0] cby_1__1__26_left_grid_pin_9_ ;
wire [0:0] cby_1__1__26_right_grid_pin_52_ ;
wire [0:0] cby_1__1__27_ccff_tail ;
wire [0:19] cby_1__1__27_chany_bottom_out ;
wire [0:19] cby_1__1__27_chany_top_out ;
wire [0:0] cby_1__1__27_left_grid_pin_0_ ;
wire [0:0] cby_1__1__27_left_grid_pin_10_ ;
wire [0:0] cby_1__1__27_left_grid_pin_11_ ;
wire [0:0] cby_1__1__27_left_grid_pin_12_ ;
wire [0:0] cby_1__1__27_left_grid_pin_13_ ;
wire [0:0] cby_1__1__27_left_grid_pin_14_ ;
wire [0:0] cby_1__1__27_left_grid_pin_15_ ;
wire [0:0] cby_1__1__27_left_grid_pin_1_ ;
wire [0:0] cby_1__1__27_left_grid_pin_2_ ;
wire [0:0] cby_1__1__27_left_grid_pin_3_ ;
wire [0:0] cby_1__1__27_left_grid_pin_4_ ;
wire [0:0] cby_1__1__27_left_grid_pin_5_ ;
wire [0:0] cby_1__1__27_left_grid_pin_6_ ;
wire [0:0] cby_1__1__27_left_grid_pin_7_ ;
wire [0:0] cby_1__1__27_left_grid_pin_8_ ;
wire [0:0] cby_1__1__27_left_grid_pin_9_ ;
wire [0:0] cby_1__1__27_right_grid_pin_52_ ;
wire [0:0] cby_1__1__28_ccff_tail ;
wire [0:19] cby_1__1__28_chany_bottom_out ;
wire [0:19] cby_1__1__28_chany_top_out ;
wire [0:0] cby_1__1__28_left_grid_pin_0_ ;
wire [0:0] cby_1__1__28_left_grid_pin_10_ ;
wire [0:0] cby_1__1__28_left_grid_pin_11_ ;
wire [0:0] cby_1__1__28_left_grid_pin_12_ ;
wire [0:0] cby_1__1__28_left_grid_pin_13_ ;
wire [0:0] cby_1__1__28_left_grid_pin_14_ ;
wire [0:0] cby_1__1__28_left_grid_pin_15_ ;
wire [0:0] cby_1__1__28_left_grid_pin_1_ ;
wire [0:0] cby_1__1__28_left_grid_pin_2_ ;
wire [0:0] cby_1__1__28_left_grid_pin_3_ ;
wire [0:0] cby_1__1__28_left_grid_pin_4_ ;
wire [0:0] cby_1__1__28_left_grid_pin_5_ ;
wire [0:0] cby_1__1__28_left_grid_pin_6_ ;
wire [0:0] cby_1__1__28_left_grid_pin_7_ ;
wire [0:0] cby_1__1__28_left_grid_pin_8_ ;
wire [0:0] cby_1__1__28_left_grid_pin_9_ ;
wire [0:0] cby_1__1__28_right_grid_pin_52_ ;
wire [0:0] cby_1__1__29_ccff_tail ;
wire [0:19] cby_1__1__29_chany_bottom_out ;
wire [0:19] cby_1__1__29_chany_top_out ;
wire [0:0] cby_1__1__29_left_grid_pin_0_ ;
wire [0:0] cby_1__1__29_left_grid_pin_10_ ;
wire [0:0] cby_1__1__29_left_grid_pin_11_ ;
wire [0:0] cby_1__1__29_left_grid_pin_12_ ;
wire [0:0] cby_1__1__29_left_grid_pin_13_ ;
wire [0:0] cby_1__1__29_left_grid_pin_14_ ;
wire [0:0] cby_1__1__29_left_grid_pin_15_ ;
wire [0:0] cby_1__1__29_left_grid_pin_1_ ;
wire [0:0] cby_1__1__29_left_grid_pin_2_ ;
wire [0:0] cby_1__1__29_left_grid_pin_3_ ;
wire [0:0] cby_1__1__29_left_grid_pin_4_ ;
wire [0:0] cby_1__1__29_left_grid_pin_5_ ;
wire [0:0] cby_1__1__29_left_grid_pin_6_ ;
wire [0:0] cby_1__1__29_left_grid_pin_7_ ;
wire [0:0] cby_1__1__29_left_grid_pin_8_ ;
wire [0:0] cby_1__1__29_left_grid_pin_9_ ;
wire [0:0] cby_1__1__29_right_grid_pin_52_ ;
wire [0:0] cby_1__1__2_ccff_tail ;
wire [0:19] cby_1__1__2_chany_bottom_out ;
wire [0:19] cby_1__1__2_chany_top_out ;
wire [0:0] cby_1__1__2_left_grid_pin_0_ ;
wire [0:0] cby_1__1__2_left_grid_pin_10_ ;
wire [0:0] cby_1__1__2_left_grid_pin_11_ ;
wire [0:0] cby_1__1__2_left_grid_pin_12_ ;
wire [0:0] cby_1__1__2_left_grid_pin_13_ ;
wire [0:0] cby_1__1__2_left_grid_pin_14_ ;
wire [0:0] cby_1__1__2_left_grid_pin_15_ ;
wire [0:0] cby_1__1__2_left_grid_pin_1_ ;
wire [0:0] cby_1__1__2_left_grid_pin_2_ ;
wire [0:0] cby_1__1__2_left_grid_pin_3_ ;
wire [0:0] cby_1__1__2_left_grid_pin_4_ ;
wire [0:0] cby_1__1__2_left_grid_pin_5_ ;
wire [0:0] cby_1__1__2_left_grid_pin_6_ ;
wire [0:0] cby_1__1__2_left_grid_pin_7_ ;
wire [0:0] cby_1__1__2_left_grid_pin_8_ ;
wire [0:0] cby_1__1__2_left_grid_pin_9_ ;
wire [0:0] cby_1__1__2_right_grid_pin_52_ ;
wire [0:0] cby_1__1__30_ccff_tail ;
wire [0:19] cby_1__1__30_chany_bottom_out ;
wire [0:19] cby_1__1__30_chany_top_out ;
wire [0:0] cby_1__1__30_left_grid_pin_0_ ;
wire [0:0] cby_1__1__30_left_grid_pin_10_ ;
wire [0:0] cby_1__1__30_left_grid_pin_11_ ;
wire [0:0] cby_1__1__30_left_grid_pin_12_ ;
wire [0:0] cby_1__1__30_left_grid_pin_13_ ;
wire [0:0] cby_1__1__30_left_grid_pin_14_ ;
wire [0:0] cby_1__1__30_left_grid_pin_15_ ;
wire [0:0] cby_1__1__30_left_grid_pin_1_ ;
wire [0:0] cby_1__1__30_left_grid_pin_2_ ;
wire [0:0] cby_1__1__30_left_grid_pin_3_ ;
wire [0:0] cby_1__1__30_left_grid_pin_4_ ;
wire [0:0] cby_1__1__30_left_grid_pin_5_ ;
wire [0:0] cby_1__1__30_left_grid_pin_6_ ;
wire [0:0] cby_1__1__30_left_grid_pin_7_ ;
wire [0:0] cby_1__1__30_left_grid_pin_8_ ;
wire [0:0] cby_1__1__30_left_grid_pin_9_ ;
wire [0:0] cby_1__1__30_right_grid_pin_52_ ;
wire [0:0] cby_1__1__31_ccff_tail ;
wire [0:19] cby_1__1__31_chany_bottom_out ;
wire [0:19] cby_1__1__31_chany_top_out ;
wire [0:0] cby_1__1__31_left_grid_pin_0_ ;
wire [0:0] cby_1__1__31_left_grid_pin_10_ ;
wire [0:0] cby_1__1__31_left_grid_pin_11_ ;
wire [0:0] cby_1__1__31_left_grid_pin_12_ ;
wire [0:0] cby_1__1__31_left_grid_pin_13_ ;
wire [0:0] cby_1__1__31_left_grid_pin_14_ ;
wire [0:0] cby_1__1__31_left_grid_pin_15_ ;
wire [0:0] cby_1__1__31_left_grid_pin_1_ ;
wire [0:0] cby_1__1__31_left_grid_pin_2_ ;
wire [0:0] cby_1__1__31_left_grid_pin_3_ ;
wire [0:0] cby_1__1__31_left_grid_pin_4_ ;
wire [0:0] cby_1__1__31_left_grid_pin_5_ ;
wire [0:0] cby_1__1__31_left_grid_pin_6_ ;
wire [0:0] cby_1__1__31_left_grid_pin_7_ ;
wire [0:0] cby_1__1__31_left_grid_pin_8_ ;
wire [0:0] cby_1__1__31_left_grid_pin_9_ ;
wire [0:0] cby_1__1__31_right_grid_pin_52_ ;
wire [0:0] cby_1__1__32_ccff_tail ;
wire [0:19] cby_1__1__32_chany_bottom_out ;
wire [0:19] cby_1__1__32_chany_top_out ;
wire [0:0] cby_1__1__32_left_grid_pin_0_ ;
wire [0:0] cby_1__1__32_left_grid_pin_10_ ;
wire [0:0] cby_1__1__32_left_grid_pin_11_ ;
wire [0:0] cby_1__1__32_left_grid_pin_12_ ;
wire [0:0] cby_1__1__32_left_grid_pin_13_ ;
wire [0:0] cby_1__1__32_left_grid_pin_14_ ;
wire [0:0] cby_1__1__32_left_grid_pin_15_ ;
wire [0:0] cby_1__1__32_left_grid_pin_1_ ;
wire [0:0] cby_1__1__32_left_grid_pin_2_ ;
wire [0:0] cby_1__1__32_left_grid_pin_3_ ;
wire [0:0] cby_1__1__32_left_grid_pin_4_ ;
wire [0:0] cby_1__1__32_left_grid_pin_5_ ;
wire [0:0] cby_1__1__32_left_grid_pin_6_ ;
wire [0:0] cby_1__1__32_left_grid_pin_7_ ;
wire [0:0] cby_1__1__32_left_grid_pin_8_ ;
wire [0:0] cby_1__1__32_left_grid_pin_9_ ;
wire [0:0] cby_1__1__32_right_grid_pin_52_ ;
wire [0:0] cby_1__1__33_ccff_tail ;
wire [0:19] cby_1__1__33_chany_bottom_out ;
wire [0:19] cby_1__1__33_chany_top_out ;
wire [0:0] cby_1__1__33_left_grid_pin_0_ ;
wire [0:0] cby_1__1__33_left_grid_pin_10_ ;
wire [0:0] cby_1__1__33_left_grid_pin_11_ ;
wire [0:0] cby_1__1__33_left_grid_pin_12_ ;
wire [0:0] cby_1__1__33_left_grid_pin_13_ ;
wire [0:0] cby_1__1__33_left_grid_pin_14_ ;
wire [0:0] cby_1__1__33_left_grid_pin_15_ ;
wire [0:0] cby_1__1__33_left_grid_pin_1_ ;
wire [0:0] cby_1__1__33_left_grid_pin_2_ ;
wire [0:0] cby_1__1__33_left_grid_pin_3_ ;
wire [0:0] cby_1__1__33_left_grid_pin_4_ ;
wire [0:0] cby_1__1__33_left_grid_pin_5_ ;
wire [0:0] cby_1__1__33_left_grid_pin_6_ ;
wire [0:0] cby_1__1__33_left_grid_pin_7_ ;
wire [0:0] cby_1__1__33_left_grid_pin_8_ ;
wire [0:0] cby_1__1__33_left_grid_pin_9_ ;
wire [0:0] cby_1__1__33_right_grid_pin_52_ ;
wire [0:0] cby_1__1__34_ccff_tail ;
wire [0:19] cby_1__1__34_chany_bottom_out ;
wire [0:19] cby_1__1__34_chany_top_out ;
wire [0:0] cby_1__1__34_left_grid_pin_0_ ;
wire [0:0] cby_1__1__34_left_grid_pin_10_ ;
wire [0:0] cby_1__1__34_left_grid_pin_11_ ;
wire [0:0] cby_1__1__34_left_grid_pin_12_ ;
wire [0:0] cby_1__1__34_left_grid_pin_13_ ;
wire [0:0] cby_1__1__34_left_grid_pin_14_ ;
wire [0:0] cby_1__1__34_left_grid_pin_15_ ;
wire [0:0] cby_1__1__34_left_grid_pin_1_ ;
wire [0:0] cby_1__1__34_left_grid_pin_2_ ;
wire [0:0] cby_1__1__34_left_grid_pin_3_ ;
wire [0:0] cby_1__1__34_left_grid_pin_4_ ;
wire [0:0] cby_1__1__34_left_grid_pin_5_ ;
wire [0:0] cby_1__1__34_left_grid_pin_6_ ;
wire [0:0] cby_1__1__34_left_grid_pin_7_ ;
wire [0:0] cby_1__1__34_left_grid_pin_8_ ;
wire [0:0] cby_1__1__34_left_grid_pin_9_ ;
wire [0:0] cby_1__1__34_right_grid_pin_52_ ;
wire [0:0] cby_1__1__35_ccff_tail ;
wire [0:19] cby_1__1__35_chany_bottom_out ;
wire [0:19] cby_1__1__35_chany_top_out ;
wire [0:0] cby_1__1__35_left_grid_pin_0_ ;
wire [0:0] cby_1__1__35_left_grid_pin_10_ ;
wire [0:0] cby_1__1__35_left_grid_pin_11_ ;
wire [0:0] cby_1__1__35_left_grid_pin_12_ ;
wire [0:0] cby_1__1__35_left_grid_pin_13_ ;
wire [0:0] cby_1__1__35_left_grid_pin_14_ ;
wire [0:0] cby_1__1__35_left_grid_pin_15_ ;
wire [0:0] cby_1__1__35_left_grid_pin_1_ ;
wire [0:0] cby_1__1__35_left_grid_pin_2_ ;
wire [0:0] cby_1__1__35_left_grid_pin_3_ ;
wire [0:0] cby_1__1__35_left_grid_pin_4_ ;
wire [0:0] cby_1__1__35_left_grid_pin_5_ ;
wire [0:0] cby_1__1__35_left_grid_pin_6_ ;
wire [0:0] cby_1__1__35_left_grid_pin_7_ ;
wire [0:0] cby_1__1__35_left_grid_pin_8_ ;
wire [0:0] cby_1__1__35_left_grid_pin_9_ ;
wire [0:0] cby_1__1__35_right_grid_pin_52_ ;
wire [0:0] cby_1__1__36_ccff_tail ;
wire [0:19] cby_1__1__36_chany_bottom_out ;
wire [0:19] cby_1__1__36_chany_top_out ;
wire [0:0] cby_1__1__36_left_grid_pin_0_ ;
wire [0:0] cby_1__1__36_left_grid_pin_10_ ;
wire [0:0] cby_1__1__36_left_grid_pin_11_ ;
wire [0:0] cby_1__1__36_left_grid_pin_12_ ;
wire [0:0] cby_1__1__36_left_grid_pin_13_ ;
wire [0:0] cby_1__1__36_left_grid_pin_14_ ;
wire [0:0] cby_1__1__36_left_grid_pin_15_ ;
wire [0:0] cby_1__1__36_left_grid_pin_1_ ;
wire [0:0] cby_1__1__36_left_grid_pin_2_ ;
wire [0:0] cby_1__1__36_left_grid_pin_3_ ;
wire [0:0] cby_1__1__36_left_grid_pin_4_ ;
wire [0:0] cby_1__1__36_left_grid_pin_5_ ;
wire [0:0] cby_1__1__36_left_grid_pin_6_ ;
wire [0:0] cby_1__1__36_left_grid_pin_7_ ;
wire [0:0] cby_1__1__36_left_grid_pin_8_ ;
wire [0:0] cby_1__1__36_left_grid_pin_9_ ;
wire [0:0] cby_1__1__36_right_grid_pin_52_ ;
wire [0:0] cby_1__1__37_ccff_tail ;
wire [0:19] cby_1__1__37_chany_bottom_out ;
wire [0:19] cby_1__1__37_chany_top_out ;
wire [0:0] cby_1__1__37_left_grid_pin_0_ ;
wire [0:0] cby_1__1__37_left_grid_pin_10_ ;
wire [0:0] cby_1__1__37_left_grid_pin_11_ ;
wire [0:0] cby_1__1__37_left_grid_pin_12_ ;
wire [0:0] cby_1__1__37_left_grid_pin_13_ ;
wire [0:0] cby_1__1__37_left_grid_pin_14_ ;
wire [0:0] cby_1__1__37_left_grid_pin_15_ ;
wire [0:0] cby_1__1__37_left_grid_pin_1_ ;
wire [0:0] cby_1__1__37_left_grid_pin_2_ ;
wire [0:0] cby_1__1__37_left_grid_pin_3_ ;
wire [0:0] cby_1__1__37_left_grid_pin_4_ ;
wire [0:0] cby_1__1__37_left_grid_pin_5_ ;
wire [0:0] cby_1__1__37_left_grid_pin_6_ ;
wire [0:0] cby_1__1__37_left_grid_pin_7_ ;
wire [0:0] cby_1__1__37_left_grid_pin_8_ ;
wire [0:0] cby_1__1__37_left_grid_pin_9_ ;
wire [0:0] cby_1__1__37_right_grid_pin_52_ ;
wire [0:0] cby_1__1__38_ccff_tail ;
wire [0:19] cby_1__1__38_chany_bottom_out ;
wire [0:19] cby_1__1__38_chany_top_out ;
wire [0:0] cby_1__1__38_left_grid_pin_0_ ;
wire [0:0] cby_1__1__38_left_grid_pin_10_ ;
wire [0:0] cby_1__1__38_left_grid_pin_11_ ;
wire [0:0] cby_1__1__38_left_grid_pin_12_ ;
wire [0:0] cby_1__1__38_left_grid_pin_13_ ;
wire [0:0] cby_1__1__38_left_grid_pin_14_ ;
wire [0:0] cby_1__1__38_left_grid_pin_15_ ;
wire [0:0] cby_1__1__38_left_grid_pin_1_ ;
wire [0:0] cby_1__1__38_left_grid_pin_2_ ;
wire [0:0] cby_1__1__38_left_grid_pin_3_ ;
wire [0:0] cby_1__1__38_left_grid_pin_4_ ;
wire [0:0] cby_1__1__38_left_grid_pin_5_ ;
wire [0:0] cby_1__1__38_left_grid_pin_6_ ;
wire [0:0] cby_1__1__38_left_grid_pin_7_ ;
wire [0:0] cby_1__1__38_left_grid_pin_8_ ;
wire [0:0] cby_1__1__38_left_grid_pin_9_ ;
wire [0:0] cby_1__1__38_right_grid_pin_52_ ;
wire [0:0] cby_1__1__39_ccff_tail ;
wire [0:19] cby_1__1__39_chany_bottom_out ;
wire [0:19] cby_1__1__39_chany_top_out ;
wire [0:0] cby_1__1__39_left_grid_pin_0_ ;
wire [0:0] cby_1__1__39_left_grid_pin_10_ ;
wire [0:0] cby_1__1__39_left_grid_pin_11_ ;
wire [0:0] cby_1__1__39_left_grid_pin_12_ ;
wire [0:0] cby_1__1__39_left_grid_pin_13_ ;
wire [0:0] cby_1__1__39_left_grid_pin_14_ ;
wire [0:0] cby_1__1__39_left_grid_pin_15_ ;
wire [0:0] cby_1__1__39_left_grid_pin_1_ ;
wire [0:0] cby_1__1__39_left_grid_pin_2_ ;
wire [0:0] cby_1__1__39_left_grid_pin_3_ ;
wire [0:0] cby_1__1__39_left_grid_pin_4_ ;
wire [0:0] cby_1__1__39_left_grid_pin_5_ ;
wire [0:0] cby_1__1__39_left_grid_pin_6_ ;
wire [0:0] cby_1__1__39_left_grid_pin_7_ ;
wire [0:0] cby_1__1__39_left_grid_pin_8_ ;
wire [0:0] cby_1__1__39_left_grid_pin_9_ ;
wire [0:0] cby_1__1__39_right_grid_pin_52_ ;
wire [0:0] cby_1__1__3_ccff_tail ;
wire [0:19] cby_1__1__3_chany_bottom_out ;
wire [0:19] cby_1__1__3_chany_top_out ;
wire [0:0] cby_1__1__3_left_grid_pin_0_ ;
wire [0:0] cby_1__1__3_left_grid_pin_10_ ;
wire [0:0] cby_1__1__3_left_grid_pin_11_ ;
wire [0:0] cby_1__1__3_left_grid_pin_12_ ;
wire [0:0] cby_1__1__3_left_grid_pin_13_ ;
wire [0:0] cby_1__1__3_left_grid_pin_14_ ;
wire [0:0] cby_1__1__3_left_grid_pin_15_ ;
wire [0:0] cby_1__1__3_left_grid_pin_1_ ;
wire [0:0] cby_1__1__3_left_grid_pin_2_ ;
wire [0:0] cby_1__1__3_left_grid_pin_3_ ;
wire [0:0] cby_1__1__3_left_grid_pin_4_ ;
wire [0:0] cby_1__1__3_left_grid_pin_5_ ;
wire [0:0] cby_1__1__3_left_grid_pin_6_ ;
wire [0:0] cby_1__1__3_left_grid_pin_7_ ;
wire [0:0] cby_1__1__3_left_grid_pin_8_ ;
wire [0:0] cby_1__1__3_left_grid_pin_9_ ;
wire [0:0] cby_1__1__3_right_grid_pin_52_ ;
wire [0:0] cby_1__1__40_ccff_tail ;
wire [0:19] cby_1__1__40_chany_bottom_out ;
wire [0:19] cby_1__1__40_chany_top_out ;
wire [0:0] cby_1__1__40_left_grid_pin_0_ ;
wire [0:0] cby_1__1__40_left_grid_pin_10_ ;
wire [0:0] cby_1__1__40_left_grid_pin_11_ ;
wire [0:0] cby_1__1__40_left_grid_pin_12_ ;
wire [0:0] cby_1__1__40_left_grid_pin_13_ ;
wire [0:0] cby_1__1__40_left_grid_pin_14_ ;
wire [0:0] cby_1__1__40_left_grid_pin_15_ ;
wire [0:0] cby_1__1__40_left_grid_pin_1_ ;
wire [0:0] cby_1__1__40_left_grid_pin_2_ ;
wire [0:0] cby_1__1__40_left_grid_pin_3_ ;
wire [0:0] cby_1__1__40_left_grid_pin_4_ ;
wire [0:0] cby_1__1__40_left_grid_pin_5_ ;
wire [0:0] cby_1__1__40_left_grid_pin_6_ ;
wire [0:0] cby_1__1__40_left_grid_pin_7_ ;
wire [0:0] cby_1__1__40_left_grid_pin_8_ ;
wire [0:0] cby_1__1__40_left_grid_pin_9_ ;
wire [0:0] cby_1__1__40_right_grid_pin_52_ ;
wire [0:0] cby_1__1__41_ccff_tail ;
wire [0:19] cby_1__1__41_chany_bottom_out ;
wire [0:19] cby_1__1__41_chany_top_out ;
wire [0:0] cby_1__1__41_left_grid_pin_0_ ;
wire [0:0] cby_1__1__41_left_grid_pin_10_ ;
wire [0:0] cby_1__1__41_left_grid_pin_11_ ;
wire [0:0] cby_1__1__41_left_grid_pin_12_ ;
wire [0:0] cby_1__1__41_left_grid_pin_13_ ;
wire [0:0] cby_1__1__41_left_grid_pin_14_ ;
wire [0:0] cby_1__1__41_left_grid_pin_15_ ;
wire [0:0] cby_1__1__41_left_grid_pin_1_ ;
wire [0:0] cby_1__1__41_left_grid_pin_2_ ;
wire [0:0] cby_1__1__41_left_grid_pin_3_ ;
wire [0:0] cby_1__1__41_left_grid_pin_4_ ;
wire [0:0] cby_1__1__41_left_grid_pin_5_ ;
wire [0:0] cby_1__1__41_left_grid_pin_6_ ;
wire [0:0] cby_1__1__41_left_grid_pin_7_ ;
wire [0:0] cby_1__1__41_left_grid_pin_8_ ;
wire [0:0] cby_1__1__41_left_grid_pin_9_ ;
wire [0:0] cby_1__1__41_right_grid_pin_52_ ;
wire [0:0] cby_1__1__42_ccff_tail ;
wire [0:19] cby_1__1__42_chany_bottom_out ;
wire [0:19] cby_1__1__42_chany_top_out ;
wire [0:0] cby_1__1__42_left_grid_pin_0_ ;
wire [0:0] cby_1__1__42_left_grid_pin_10_ ;
wire [0:0] cby_1__1__42_left_grid_pin_11_ ;
wire [0:0] cby_1__1__42_left_grid_pin_12_ ;
wire [0:0] cby_1__1__42_left_grid_pin_13_ ;
wire [0:0] cby_1__1__42_left_grid_pin_14_ ;
wire [0:0] cby_1__1__42_left_grid_pin_15_ ;
wire [0:0] cby_1__1__42_left_grid_pin_1_ ;
wire [0:0] cby_1__1__42_left_grid_pin_2_ ;
wire [0:0] cby_1__1__42_left_grid_pin_3_ ;
wire [0:0] cby_1__1__42_left_grid_pin_4_ ;
wire [0:0] cby_1__1__42_left_grid_pin_5_ ;
wire [0:0] cby_1__1__42_left_grid_pin_6_ ;
wire [0:0] cby_1__1__42_left_grid_pin_7_ ;
wire [0:0] cby_1__1__42_left_grid_pin_8_ ;
wire [0:0] cby_1__1__42_left_grid_pin_9_ ;
wire [0:0] cby_1__1__42_right_grid_pin_52_ ;
wire [0:0] cby_1__1__43_ccff_tail ;
wire [0:19] cby_1__1__43_chany_bottom_out ;
wire [0:19] cby_1__1__43_chany_top_out ;
wire [0:0] cby_1__1__43_left_grid_pin_0_ ;
wire [0:0] cby_1__1__43_left_grid_pin_10_ ;
wire [0:0] cby_1__1__43_left_grid_pin_11_ ;
wire [0:0] cby_1__1__43_left_grid_pin_12_ ;
wire [0:0] cby_1__1__43_left_grid_pin_13_ ;
wire [0:0] cby_1__1__43_left_grid_pin_14_ ;
wire [0:0] cby_1__1__43_left_grid_pin_15_ ;
wire [0:0] cby_1__1__43_left_grid_pin_1_ ;
wire [0:0] cby_1__1__43_left_grid_pin_2_ ;
wire [0:0] cby_1__1__43_left_grid_pin_3_ ;
wire [0:0] cby_1__1__43_left_grid_pin_4_ ;
wire [0:0] cby_1__1__43_left_grid_pin_5_ ;
wire [0:0] cby_1__1__43_left_grid_pin_6_ ;
wire [0:0] cby_1__1__43_left_grid_pin_7_ ;
wire [0:0] cby_1__1__43_left_grid_pin_8_ ;
wire [0:0] cby_1__1__43_left_grid_pin_9_ ;
wire [0:0] cby_1__1__43_right_grid_pin_52_ ;
wire [0:0] cby_1__1__44_ccff_tail ;
wire [0:19] cby_1__1__44_chany_bottom_out ;
wire [0:19] cby_1__1__44_chany_top_out ;
wire [0:0] cby_1__1__44_left_grid_pin_0_ ;
wire [0:0] cby_1__1__44_left_grid_pin_10_ ;
wire [0:0] cby_1__1__44_left_grid_pin_11_ ;
wire [0:0] cby_1__1__44_left_grid_pin_12_ ;
wire [0:0] cby_1__1__44_left_grid_pin_13_ ;
wire [0:0] cby_1__1__44_left_grid_pin_14_ ;
wire [0:0] cby_1__1__44_left_grid_pin_15_ ;
wire [0:0] cby_1__1__44_left_grid_pin_1_ ;
wire [0:0] cby_1__1__44_left_grid_pin_2_ ;
wire [0:0] cby_1__1__44_left_grid_pin_3_ ;
wire [0:0] cby_1__1__44_left_grid_pin_4_ ;
wire [0:0] cby_1__1__44_left_grid_pin_5_ ;
wire [0:0] cby_1__1__44_left_grid_pin_6_ ;
wire [0:0] cby_1__1__44_left_grid_pin_7_ ;
wire [0:0] cby_1__1__44_left_grid_pin_8_ ;
wire [0:0] cby_1__1__44_left_grid_pin_9_ ;
wire [0:0] cby_1__1__44_right_grid_pin_52_ ;
wire [0:0] cby_1__1__45_ccff_tail ;
wire [0:19] cby_1__1__45_chany_bottom_out ;
wire [0:19] cby_1__1__45_chany_top_out ;
wire [0:0] cby_1__1__45_left_grid_pin_0_ ;
wire [0:0] cby_1__1__45_left_grid_pin_10_ ;
wire [0:0] cby_1__1__45_left_grid_pin_11_ ;
wire [0:0] cby_1__1__45_left_grid_pin_12_ ;
wire [0:0] cby_1__1__45_left_grid_pin_13_ ;
wire [0:0] cby_1__1__45_left_grid_pin_14_ ;
wire [0:0] cby_1__1__45_left_grid_pin_15_ ;
wire [0:0] cby_1__1__45_left_grid_pin_1_ ;
wire [0:0] cby_1__1__45_left_grid_pin_2_ ;
wire [0:0] cby_1__1__45_left_grid_pin_3_ ;
wire [0:0] cby_1__1__45_left_grid_pin_4_ ;
wire [0:0] cby_1__1__45_left_grid_pin_5_ ;
wire [0:0] cby_1__1__45_left_grid_pin_6_ ;
wire [0:0] cby_1__1__45_left_grid_pin_7_ ;
wire [0:0] cby_1__1__45_left_grid_pin_8_ ;
wire [0:0] cby_1__1__45_left_grid_pin_9_ ;
wire [0:0] cby_1__1__45_right_grid_pin_52_ ;
wire [0:0] cby_1__1__46_ccff_tail ;
wire [0:19] cby_1__1__46_chany_bottom_out ;
wire [0:19] cby_1__1__46_chany_top_out ;
wire [0:0] cby_1__1__46_left_grid_pin_0_ ;
wire [0:0] cby_1__1__46_left_grid_pin_10_ ;
wire [0:0] cby_1__1__46_left_grid_pin_11_ ;
wire [0:0] cby_1__1__46_left_grid_pin_12_ ;
wire [0:0] cby_1__1__46_left_grid_pin_13_ ;
wire [0:0] cby_1__1__46_left_grid_pin_14_ ;
wire [0:0] cby_1__1__46_left_grid_pin_15_ ;
wire [0:0] cby_1__1__46_left_grid_pin_1_ ;
wire [0:0] cby_1__1__46_left_grid_pin_2_ ;
wire [0:0] cby_1__1__46_left_grid_pin_3_ ;
wire [0:0] cby_1__1__46_left_grid_pin_4_ ;
wire [0:0] cby_1__1__46_left_grid_pin_5_ ;
wire [0:0] cby_1__1__46_left_grid_pin_6_ ;
wire [0:0] cby_1__1__46_left_grid_pin_7_ ;
wire [0:0] cby_1__1__46_left_grid_pin_8_ ;
wire [0:0] cby_1__1__46_left_grid_pin_9_ ;
wire [0:0] cby_1__1__46_right_grid_pin_52_ ;
wire [0:0] cby_1__1__47_ccff_tail ;
wire [0:19] cby_1__1__47_chany_bottom_out ;
wire [0:19] cby_1__1__47_chany_top_out ;
wire [0:0] cby_1__1__47_left_grid_pin_0_ ;
wire [0:0] cby_1__1__47_left_grid_pin_10_ ;
wire [0:0] cby_1__1__47_left_grid_pin_11_ ;
wire [0:0] cby_1__1__47_left_grid_pin_12_ ;
wire [0:0] cby_1__1__47_left_grid_pin_13_ ;
wire [0:0] cby_1__1__47_left_grid_pin_14_ ;
wire [0:0] cby_1__1__47_left_grid_pin_15_ ;
wire [0:0] cby_1__1__47_left_grid_pin_1_ ;
wire [0:0] cby_1__1__47_left_grid_pin_2_ ;
wire [0:0] cby_1__1__47_left_grid_pin_3_ ;
wire [0:0] cby_1__1__47_left_grid_pin_4_ ;
wire [0:0] cby_1__1__47_left_grid_pin_5_ ;
wire [0:0] cby_1__1__47_left_grid_pin_6_ ;
wire [0:0] cby_1__1__47_left_grid_pin_7_ ;
wire [0:0] cby_1__1__47_left_grid_pin_8_ ;
wire [0:0] cby_1__1__47_left_grid_pin_9_ ;
wire [0:0] cby_1__1__47_right_grid_pin_52_ ;
wire [0:0] cby_1__1__48_ccff_tail ;
wire [0:19] cby_1__1__48_chany_bottom_out ;
wire [0:19] cby_1__1__48_chany_top_out ;
wire [0:0] cby_1__1__48_left_grid_pin_0_ ;
wire [0:0] cby_1__1__48_left_grid_pin_10_ ;
wire [0:0] cby_1__1__48_left_grid_pin_11_ ;
wire [0:0] cby_1__1__48_left_grid_pin_12_ ;
wire [0:0] cby_1__1__48_left_grid_pin_13_ ;
wire [0:0] cby_1__1__48_left_grid_pin_14_ ;
wire [0:0] cby_1__1__48_left_grid_pin_15_ ;
wire [0:0] cby_1__1__48_left_grid_pin_1_ ;
wire [0:0] cby_1__1__48_left_grid_pin_2_ ;
wire [0:0] cby_1__1__48_left_grid_pin_3_ ;
wire [0:0] cby_1__1__48_left_grid_pin_4_ ;
wire [0:0] cby_1__1__48_left_grid_pin_5_ ;
wire [0:0] cby_1__1__48_left_grid_pin_6_ ;
wire [0:0] cby_1__1__48_left_grid_pin_7_ ;
wire [0:0] cby_1__1__48_left_grid_pin_8_ ;
wire [0:0] cby_1__1__48_left_grid_pin_9_ ;
wire [0:0] cby_1__1__48_right_grid_pin_52_ ;
wire [0:0] cby_1__1__49_ccff_tail ;
wire [0:19] cby_1__1__49_chany_bottom_out ;
wire [0:19] cby_1__1__49_chany_top_out ;
wire [0:0] cby_1__1__49_left_grid_pin_0_ ;
wire [0:0] cby_1__1__49_left_grid_pin_10_ ;
wire [0:0] cby_1__1__49_left_grid_pin_11_ ;
wire [0:0] cby_1__1__49_left_grid_pin_12_ ;
wire [0:0] cby_1__1__49_left_grid_pin_13_ ;
wire [0:0] cby_1__1__49_left_grid_pin_14_ ;
wire [0:0] cby_1__1__49_left_grid_pin_15_ ;
wire [0:0] cby_1__1__49_left_grid_pin_1_ ;
wire [0:0] cby_1__1__49_left_grid_pin_2_ ;
wire [0:0] cby_1__1__49_left_grid_pin_3_ ;
wire [0:0] cby_1__1__49_left_grid_pin_4_ ;
wire [0:0] cby_1__1__49_left_grid_pin_5_ ;
wire [0:0] cby_1__1__49_left_grid_pin_6_ ;
wire [0:0] cby_1__1__49_left_grid_pin_7_ ;
wire [0:0] cby_1__1__49_left_grid_pin_8_ ;
wire [0:0] cby_1__1__49_left_grid_pin_9_ ;
wire [0:0] cby_1__1__49_right_grid_pin_52_ ;
wire [0:0] cby_1__1__4_ccff_tail ;
wire [0:19] cby_1__1__4_chany_bottom_out ;
wire [0:19] cby_1__1__4_chany_top_out ;
wire [0:0] cby_1__1__4_left_grid_pin_0_ ;
wire [0:0] cby_1__1__4_left_grid_pin_10_ ;
wire [0:0] cby_1__1__4_left_grid_pin_11_ ;
wire [0:0] cby_1__1__4_left_grid_pin_12_ ;
wire [0:0] cby_1__1__4_left_grid_pin_13_ ;
wire [0:0] cby_1__1__4_left_grid_pin_14_ ;
wire [0:0] cby_1__1__4_left_grid_pin_15_ ;
wire [0:0] cby_1__1__4_left_grid_pin_1_ ;
wire [0:0] cby_1__1__4_left_grid_pin_2_ ;
wire [0:0] cby_1__1__4_left_grid_pin_3_ ;
wire [0:0] cby_1__1__4_left_grid_pin_4_ ;
wire [0:0] cby_1__1__4_left_grid_pin_5_ ;
wire [0:0] cby_1__1__4_left_grid_pin_6_ ;
wire [0:0] cby_1__1__4_left_grid_pin_7_ ;
wire [0:0] cby_1__1__4_left_grid_pin_8_ ;
wire [0:0] cby_1__1__4_left_grid_pin_9_ ;
wire [0:0] cby_1__1__4_right_grid_pin_52_ ;
wire [0:0] cby_1__1__50_ccff_tail ;
wire [0:19] cby_1__1__50_chany_bottom_out ;
wire [0:19] cby_1__1__50_chany_top_out ;
wire [0:0] cby_1__1__50_left_grid_pin_0_ ;
wire [0:0] cby_1__1__50_left_grid_pin_10_ ;
wire [0:0] cby_1__1__50_left_grid_pin_11_ ;
wire [0:0] cby_1__1__50_left_grid_pin_12_ ;
wire [0:0] cby_1__1__50_left_grid_pin_13_ ;
wire [0:0] cby_1__1__50_left_grid_pin_14_ ;
wire [0:0] cby_1__1__50_left_grid_pin_15_ ;
wire [0:0] cby_1__1__50_left_grid_pin_1_ ;
wire [0:0] cby_1__1__50_left_grid_pin_2_ ;
wire [0:0] cby_1__1__50_left_grid_pin_3_ ;
wire [0:0] cby_1__1__50_left_grid_pin_4_ ;
wire [0:0] cby_1__1__50_left_grid_pin_5_ ;
wire [0:0] cby_1__1__50_left_grid_pin_6_ ;
wire [0:0] cby_1__1__50_left_grid_pin_7_ ;
wire [0:0] cby_1__1__50_left_grid_pin_8_ ;
wire [0:0] cby_1__1__50_left_grid_pin_9_ ;
wire [0:0] cby_1__1__50_right_grid_pin_52_ ;
wire [0:0] cby_1__1__51_ccff_tail ;
wire [0:19] cby_1__1__51_chany_bottom_out ;
wire [0:19] cby_1__1__51_chany_top_out ;
wire [0:0] cby_1__1__51_left_grid_pin_0_ ;
wire [0:0] cby_1__1__51_left_grid_pin_10_ ;
wire [0:0] cby_1__1__51_left_grid_pin_11_ ;
wire [0:0] cby_1__1__51_left_grid_pin_12_ ;
wire [0:0] cby_1__1__51_left_grid_pin_13_ ;
wire [0:0] cby_1__1__51_left_grid_pin_14_ ;
wire [0:0] cby_1__1__51_left_grid_pin_15_ ;
wire [0:0] cby_1__1__51_left_grid_pin_1_ ;
wire [0:0] cby_1__1__51_left_grid_pin_2_ ;
wire [0:0] cby_1__1__51_left_grid_pin_3_ ;
wire [0:0] cby_1__1__51_left_grid_pin_4_ ;
wire [0:0] cby_1__1__51_left_grid_pin_5_ ;
wire [0:0] cby_1__1__51_left_grid_pin_6_ ;
wire [0:0] cby_1__1__51_left_grid_pin_7_ ;
wire [0:0] cby_1__1__51_left_grid_pin_8_ ;
wire [0:0] cby_1__1__51_left_grid_pin_9_ ;
wire [0:0] cby_1__1__51_right_grid_pin_52_ ;
wire [0:0] cby_1__1__52_ccff_tail ;
wire [0:19] cby_1__1__52_chany_bottom_out ;
wire [0:19] cby_1__1__52_chany_top_out ;
wire [0:0] cby_1__1__52_left_grid_pin_0_ ;
wire [0:0] cby_1__1__52_left_grid_pin_10_ ;
wire [0:0] cby_1__1__52_left_grid_pin_11_ ;
wire [0:0] cby_1__1__52_left_grid_pin_12_ ;
wire [0:0] cby_1__1__52_left_grid_pin_13_ ;
wire [0:0] cby_1__1__52_left_grid_pin_14_ ;
wire [0:0] cby_1__1__52_left_grid_pin_15_ ;
wire [0:0] cby_1__1__52_left_grid_pin_1_ ;
wire [0:0] cby_1__1__52_left_grid_pin_2_ ;
wire [0:0] cby_1__1__52_left_grid_pin_3_ ;
wire [0:0] cby_1__1__52_left_grid_pin_4_ ;
wire [0:0] cby_1__1__52_left_grid_pin_5_ ;
wire [0:0] cby_1__1__52_left_grid_pin_6_ ;
wire [0:0] cby_1__1__52_left_grid_pin_7_ ;
wire [0:0] cby_1__1__52_left_grid_pin_8_ ;
wire [0:0] cby_1__1__52_left_grid_pin_9_ ;
wire [0:0] cby_1__1__52_right_grid_pin_52_ ;
wire [0:0] cby_1__1__53_ccff_tail ;
wire [0:19] cby_1__1__53_chany_bottom_out ;
wire [0:19] cby_1__1__53_chany_top_out ;
wire [0:0] cby_1__1__53_left_grid_pin_0_ ;
wire [0:0] cby_1__1__53_left_grid_pin_10_ ;
wire [0:0] cby_1__1__53_left_grid_pin_11_ ;
wire [0:0] cby_1__1__53_left_grid_pin_12_ ;
wire [0:0] cby_1__1__53_left_grid_pin_13_ ;
wire [0:0] cby_1__1__53_left_grid_pin_14_ ;
wire [0:0] cby_1__1__53_left_grid_pin_15_ ;
wire [0:0] cby_1__1__53_left_grid_pin_1_ ;
wire [0:0] cby_1__1__53_left_grid_pin_2_ ;
wire [0:0] cby_1__1__53_left_grid_pin_3_ ;
wire [0:0] cby_1__1__53_left_grid_pin_4_ ;
wire [0:0] cby_1__1__53_left_grid_pin_5_ ;
wire [0:0] cby_1__1__53_left_grid_pin_6_ ;
wire [0:0] cby_1__1__53_left_grid_pin_7_ ;
wire [0:0] cby_1__1__53_left_grid_pin_8_ ;
wire [0:0] cby_1__1__53_left_grid_pin_9_ ;
wire [0:0] cby_1__1__53_right_grid_pin_52_ ;
wire [0:0] cby_1__1__54_ccff_tail ;
wire [0:19] cby_1__1__54_chany_bottom_out ;
wire [0:19] cby_1__1__54_chany_top_out ;
wire [0:0] cby_1__1__54_left_grid_pin_0_ ;
wire [0:0] cby_1__1__54_left_grid_pin_10_ ;
wire [0:0] cby_1__1__54_left_grid_pin_11_ ;
wire [0:0] cby_1__1__54_left_grid_pin_12_ ;
wire [0:0] cby_1__1__54_left_grid_pin_13_ ;
wire [0:0] cby_1__1__54_left_grid_pin_14_ ;
wire [0:0] cby_1__1__54_left_grid_pin_15_ ;
wire [0:0] cby_1__1__54_left_grid_pin_1_ ;
wire [0:0] cby_1__1__54_left_grid_pin_2_ ;
wire [0:0] cby_1__1__54_left_grid_pin_3_ ;
wire [0:0] cby_1__1__54_left_grid_pin_4_ ;
wire [0:0] cby_1__1__54_left_grid_pin_5_ ;
wire [0:0] cby_1__1__54_left_grid_pin_6_ ;
wire [0:0] cby_1__1__54_left_grid_pin_7_ ;
wire [0:0] cby_1__1__54_left_grid_pin_8_ ;
wire [0:0] cby_1__1__54_left_grid_pin_9_ ;
wire [0:0] cby_1__1__54_right_grid_pin_52_ ;
wire [0:0] cby_1__1__55_ccff_tail ;
wire [0:19] cby_1__1__55_chany_bottom_out ;
wire [0:19] cby_1__1__55_chany_top_out ;
wire [0:0] cby_1__1__55_left_grid_pin_0_ ;
wire [0:0] cby_1__1__55_left_grid_pin_10_ ;
wire [0:0] cby_1__1__55_left_grid_pin_11_ ;
wire [0:0] cby_1__1__55_left_grid_pin_12_ ;
wire [0:0] cby_1__1__55_left_grid_pin_13_ ;
wire [0:0] cby_1__1__55_left_grid_pin_14_ ;
wire [0:0] cby_1__1__55_left_grid_pin_15_ ;
wire [0:0] cby_1__1__55_left_grid_pin_1_ ;
wire [0:0] cby_1__1__55_left_grid_pin_2_ ;
wire [0:0] cby_1__1__55_left_grid_pin_3_ ;
wire [0:0] cby_1__1__55_left_grid_pin_4_ ;
wire [0:0] cby_1__1__55_left_grid_pin_5_ ;
wire [0:0] cby_1__1__55_left_grid_pin_6_ ;
wire [0:0] cby_1__1__55_left_grid_pin_7_ ;
wire [0:0] cby_1__1__55_left_grid_pin_8_ ;
wire [0:0] cby_1__1__55_left_grid_pin_9_ ;
wire [0:0] cby_1__1__55_right_grid_pin_52_ ;
wire [0:0] cby_1__1__56_ccff_tail ;
wire [0:19] cby_1__1__56_chany_bottom_out ;
wire [0:19] cby_1__1__56_chany_top_out ;
wire [0:0] cby_1__1__56_left_grid_pin_0_ ;
wire [0:0] cby_1__1__56_left_grid_pin_10_ ;
wire [0:0] cby_1__1__56_left_grid_pin_11_ ;
wire [0:0] cby_1__1__56_left_grid_pin_12_ ;
wire [0:0] cby_1__1__56_left_grid_pin_13_ ;
wire [0:0] cby_1__1__56_left_grid_pin_14_ ;
wire [0:0] cby_1__1__56_left_grid_pin_15_ ;
wire [0:0] cby_1__1__56_left_grid_pin_1_ ;
wire [0:0] cby_1__1__56_left_grid_pin_2_ ;
wire [0:0] cby_1__1__56_left_grid_pin_3_ ;
wire [0:0] cby_1__1__56_left_grid_pin_4_ ;
wire [0:0] cby_1__1__56_left_grid_pin_5_ ;
wire [0:0] cby_1__1__56_left_grid_pin_6_ ;
wire [0:0] cby_1__1__56_left_grid_pin_7_ ;
wire [0:0] cby_1__1__56_left_grid_pin_8_ ;
wire [0:0] cby_1__1__56_left_grid_pin_9_ ;
wire [0:0] cby_1__1__56_right_grid_pin_52_ ;
wire [0:0] cby_1__1__57_ccff_tail ;
wire [0:19] cby_1__1__57_chany_bottom_out ;
wire [0:19] cby_1__1__57_chany_top_out ;
wire [0:0] cby_1__1__57_left_grid_pin_0_ ;
wire [0:0] cby_1__1__57_left_grid_pin_10_ ;
wire [0:0] cby_1__1__57_left_grid_pin_11_ ;
wire [0:0] cby_1__1__57_left_grid_pin_12_ ;
wire [0:0] cby_1__1__57_left_grid_pin_13_ ;
wire [0:0] cby_1__1__57_left_grid_pin_14_ ;
wire [0:0] cby_1__1__57_left_grid_pin_15_ ;
wire [0:0] cby_1__1__57_left_grid_pin_1_ ;
wire [0:0] cby_1__1__57_left_grid_pin_2_ ;
wire [0:0] cby_1__1__57_left_grid_pin_3_ ;
wire [0:0] cby_1__1__57_left_grid_pin_4_ ;
wire [0:0] cby_1__1__57_left_grid_pin_5_ ;
wire [0:0] cby_1__1__57_left_grid_pin_6_ ;
wire [0:0] cby_1__1__57_left_grid_pin_7_ ;
wire [0:0] cby_1__1__57_left_grid_pin_8_ ;
wire [0:0] cby_1__1__57_left_grid_pin_9_ ;
wire [0:0] cby_1__1__57_right_grid_pin_52_ ;
wire [0:0] cby_1__1__58_ccff_tail ;
wire [0:19] cby_1__1__58_chany_bottom_out ;
wire [0:19] cby_1__1__58_chany_top_out ;
wire [0:0] cby_1__1__58_left_grid_pin_0_ ;
wire [0:0] cby_1__1__58_left_grid_pin_10_ ;
wire [0:0] cby_1__1__58_left_grid_pin_11_ ;
wire [0:0] cby_1__1__58_left_grid_pin_12_ ;
wire [0:0] cby_1__1__58_left_grid_pin_13_ ;
wire [0:0] cby_1__1__58_left_grid_pin_14_ ;
wire [0:0] cby_1__1__58_left_grid_pin_15_ ;
wire [0:0] cby_1__1__58_left_grid_pin_1_ ;
wire [0:0] cby_1__1__58_left_grid_pin_2_ ;
wire [0:0] cby_1__1__58_left_grid_pin_3_ ;
wire [0:0] cby_1__1__58_left_grid_pin_4_ ;
wire [0:0] cby_1__1__58_left_grid_pin_5_ ;
wire [0:0] cby_1__1__58_left_grid_pin_6_ ;
wire [0:0] cby_1__1__58_left_grid_pin_7_ ;
wire [0:0] cby_1__1__58_left_grid_pin_8_ ;
wire [0:0] cby_1__1__58_left_grid_pin_9_ ;
wire [0:0] cby_1__1__58_right_grid_pin_52_ ;
wire [0:0] cby_1__1__59_ccff_tail ;
wire [0:19] cby_1__1__59_chany_bottom_out ;
wire [0:19] cby_1__1__59_chany_top_out ;
wire [0:0] cby_1__1__59_left_grid_pin_0_ ;
wire [0:0] cby_1__1__59_left_grid_pin_10_ ;
wire [0:0] cby_1__1__59_left_grid_pin_11_ ;
wire [0:0] cby_1__1__59_left_grid_pin_12_ ;
wire [0:0] cby_1__1__59_left_grid_pin_13_ ;
wire [0:0] cby_1__1__59_left_grid_pin_14_ ;
wire [0:0] cby_1__1__59_left_grid_pin_15_ ;
wire [0:0] cby_1__1__59_left_grid_pin_1_ ;
wire [0:0] cby_1__1__59_left_grid_pin_2_ ;
wire [0:0] cby_1__1__59_left_grid_pin_3_ ;
wire [0:0] cby_1__1__59_left_grid_pin_4_ ;
wire [0:0] cby_1__1__59_left_grid_pin_5_ ;
wire [0:0] cby_1__1__59_left_grid_pin_6_ ;
wire [0:0] cby_1__1__59_left_grid_pin_7_ ;
wire [0:0] cby_1__1__59_left_grid_pin_8_ ;
wire [0:0] cby_1__1__59_left_grid_pin_9_ ;
wire [0:0] cby_1__1__59_right_grid_pin_52_ ;
wire [0:0] cby_1__1__5_ccff_tail ;
wire [0:19] cby_1__1__5_chany_bottom_out ;
wire [0:19] cby_1__1__5_chany_top_out ;
wire [0:0] cby_1__1__5_left_grid_pin_0_ ;
wire [0:0] cby_1__1__5_left_grid_pin_10_ ;
wire [0:0] cby_1__1__5_left_grid_pin_11_ ;
wire [0:0] cby_1__1__5_left_grid_pin_12_ ;
wire [0:0] cby_1__1__5_left_grid_pin_13_ ;
wire [0:0] cby_1__1__5_left_grid_pin_14_ ;
wire [0:0] cby_1__1__5_left_grid_pin_15_ ;
wire [0:0] cby_1__1__5_left_grid_pin_1_ ;
wire [0:0] cby_1__1__5_left_grid_pin_2_ ;
wire [0:0] cby_1__1__5_left_grid_pin_3_ ;
wire [0:0] cby_1__1__5_left_grid_pin_4_ ;
wire [0:0] cby_1__1__5_left_grid_pin_5_ ;
wire [0:0] cby_1__1__5_left_grid_pin_6_ ;
wire [0:0] cby_1__1__5_left_grid_pin_7_ ;
wire [0:0] cby_1__1__5_left_grid_pin_8_ ;
wire [0:0] cby_1__1__5_left_grid_pin_9_ ;
wire [0:0] cby_1__1__5_right_grid_pin_52_ ;
wire [0:0] cby_1__1__60_ccff_tail ;
wire [0:19] cby_1__1__60_chany_bottom_out ;
wire [0:19] cby_1__1__60_chany_top_out ;
wire [0:0] cby_1__1__60_left_grid_pin_0_ ;
wire [0:0] cby_1__1__60_left_grid_pin_10_ ;
wire [0:0] cby_1__1__60_left_grid_pin_11_ ;
wire [0:0] cby_1__1__60_left_grid_pin_12_ ;
wire [0:0] cby_1__1__60_left_grid_pin_13_ ;
wire [0:0] cby_1__1__60_left_grid_pin_14_ ;
wire [0:0] cby_1__1__60_left_grid_pin_15_ ;
wire [0:0] cby_1__1__60_left_grid_pin_1_ ;
wire [0:0] cby_1__1__60_left_grid_pin_2_ ;
wire [0:0] cby_1__1__60_left_grid_pin_3_ ;
wire [0:0] cby_1__1__60_left_grid_pin_4_ ;
wire [0:0] cby_1__1__60_left_grid_pin_5_ ;
wire [0:0] cby_1__1__60_left_grid_pin_6_ ;
wire [0:0] cby_1__1__60_left_grid_pin_7_ ;
wire [0:0] cby_1__1__60_left_grid_pin_8_ ;
wire [0:0] cby_1__1__60_left_grid_pin_9_ ;
wire [0:0] cby_1__1__60_right_grid_pin_52_ ;
wire [0:0] cby_1__1__61_ccff_tail ;
wire [0:19] cby_1__1__61_chany_bottom_out ;
wire [0:19] cby_1__1__61_chany_top_out ;
wire [0:0] cby_1__1__61_left_grid_pin_0_ ;
wire [0:0] cby_1__1__61_left_grid_pin_10_ ;
wire [0:0] cby_1__1__61_left_grid_pin_11_ ;
wire [0:0] cby_1__1__61_left_grid_pin_12_ ;
wire [0:0] cby_1__1__61_left_grid_pin_13_ ;
wire [0:0] cby_1__1__61_left_grid_pin_14_ ;
wire [0:0] cby_1__1__61_left_grid_pin_15_ ;
wire [0:0] cby_1__1__61_left_grid_pin_1_ ;
wire [0:0] cby_1__1__61_left_grid_pin_2_ ;
wire [0:0] cby_1__1__61_left_grid_pin_3_ ;
wire [0:0] cby_1__1__61_left_grid_pin_4_ ;
wire [0:0] cby_1__1__61_left_grid_pin_5_ ;
wire [0:0] cby_1__1__61_left_grid_pin_6_ ;
wire [0:0] cby_1__1__61_left_grid_pin_7_ ;
wire [0:0] cby_1__1__61_left_grid_pin_8_ ;
wire [0:0] cby_1__1__61_left_grid_pin_9_ ;
wire [0:0] cby_1__1__61_right_grid_pin_52_ ;
wire [0:0] cby_1__1__62_ccff_tail ;
wire [0:19] cby_1__1__62_chany_bottom_out ;
wire [0:19] cby_1__1__62_chany_top_out ;
wire [0:0] cby_1__1__62_left_grid_pin_0_ ;
wire [0:0] cby_1__1__62_left_grid_pin_10_ ;
wire [0:0] cby_1__1__62_left_grid_pin_11_ ;
wire [0:0] cby_1__1__62_left_grid_pin_12_ ;
wire [0:0] cby_1__1__62_left_grid_pin_13_ ;
wire [0:0] cby_1__1__62_left_grid_pin_14_ ;
wire [0:0] cby_1__1__62_left_grid_pin_15_ ;
wire [0:0] cby_1__1__62_left_grid_pin_1_ ;
wire [0:0] cby_1__1__62_left_grid_pin_2_ ;
wire [0:0] cby_1__1__62_left_grid_pin_3_ ;
wire [0:0] cby_1__1__62_left_grid_pin_4_ ;
wire [0:0] cby_1__1__62_left_grid_pin_5_ ;
wire [0:0] cby_1__1__62_left_grid_pin_6_ ;
wire [0:0] cby_1__1__62_left_grid_pin_7_ ;
wire [0:0] cby_1__1__62_left_grid_pin_8_ ;
wire [0:0] cby_1__1__62_left_grid_pin_9_ ;
wire [0:0] cby_1__1__62_right_grid_pin_52_ ;
wire [0:0] cby_1__1__63_ccff_tail ;
wire [0:19] cby_1__1__63_chany_bottom_out ;
wire [0:19] cby_1__1__63_chany_top_out ;
wire [0:0] cby_1__1__63_left_grid_pin_0_ ;
wire [0:0] cby_1__1__63_left_grid_pin_10_ ;
wire [0:0] cby_1__1__63_left_grid_pin_11_ ;
wire [0:0] cby_1__1__63_left_grid_pin_12_ ;
wire [0:0] cby_1__1__63_left_grid_pin_13_ ;
wire [0:0] cby_1__1__63_left_grid_pin_14_ ;
wire [0:0] cby_1__1__63_left_grid_pin_15_ ;
wire [0:0] cby_1__1__63_left_grid_pin_1_ ;
wire [0:0] cby_1__1__63_left_grid_pin_2_ ;
wire [0:0] cby_1__1__63_left_grid_pin_3_ ;
wire [0:0] cby_1__1__63_left_grid_pin_4_ ;
wire [0:0] cby_1__1__63_left_grid_pin_5_ ;
wire [0:0] cby_1__1__63_left_grid_pin_6_ ;
wire [0:0] cby_1__1__63_left_grid_pin_7_ ;
wire [0:0] cby_1__1__63_left_grid_pin_8_ ;
wire [0:0] cby_1__1__63_left_grid_pin_9_ ;
wire [0:0] cby_1__1__63_right_grid_pin_52_ ;
wire [0:0] cby_1__1__64_ccff_tail ;
wire [0:19] cby_1__1__64_chany_bottom_out ;
wire [0:19] cby_1__1__64_chany_top_out ;
wire [0:0] cby_1__1__64_left_grid_pin_0_ ;
wire [0:0] cby_1__1__64_left_grid_pin_10_ ;
wire [0:0] cby_1__1__64_left_grid_pin_11_ ;
wire [0:0] cby_1__1__64_left_grid_pin_12_ ;
wire [0:0] cby_1__1__64_left_grid_pin_13_ ;
wire [0:0] cby_1__1__64_left_grid_pin_14_ ;
wire [0:0] cby_1__1__64_left_grid_pin_15_ ;
wire [0:0] cby_1__1__64_left_grid_pin_1_ ;
wire [0:0] cby_1__1__64_left_grid_pin_2_ ;
wire [0:0] cby_1__1__64_left_grid_pin_3_ ;
wire [0:0] cby_1__1__64_left_grid_pin_4_ ;
wire [0:0] cby_1__1__64_left_grid_pin_5_ ;
wire [0:0] cby_1__1__64_left_grid_pin_6_ ;
wire [0:0] cby_1__1__64_left_grid_pin_7_ ;
wire [0:0] cby_1__1__64_left_grid_pin_8_ ;
wire [0:0] cby_1__1__64_left_grid_pin_9_ ;
wire [0:0] cby_1__1__64_right_grid_pin_52_ ;
wire [0:0] cby_1__1__65_ccff_tail ;
wire [0:19] cby_1__1__65_chany_bottom_out ;
wire [0:19] cby_1__1__65_chany_top_out ;
wire [0:0] cby_1__1__65_left_grid_pin_0_ ;
wire [0:0] cby_1__1__65_left_grid_pin_10_ ;
wire [0:0] cby_1__1__65_left_grid_pin_11_ ;
wire [0:0] cby_1__1__65_left_grid_pin_12_ ;
wire [0:0] cby_1__1__65_left_grid_pin_13_ ;
wire [0:0] cby_1__1__65_left_grid_pin_14_ ;
wire [0:0] cby_1__1__65_left_grid_pin_15_ ;
wire [0:0] cby_1__1__65_left_grid_pin_1_ ;
wire [0:0] cby_1__1__65_left_grid_pin_2_ ;
wire [0:0] cby_1__1__65_left_grid_pin_3_ ;
wire [0:0] cby_1__1__65_left_grid_pin_4_ ;
wire [0:0] cby_1__1__65_left_grid_pin_5_ ;
wire [0:0] cby_1__1__65_left_grid_pin_6_ ;
wire [0:0] cby_1__1__65_left_grid_pin_7_ ;
wire [0:0] cby_1__1__65_left_grid_pin_8_ ;
wire [0:0] cby_1__1__65_left_grid_pin_9_ ;
wire [0:0] cby_1__1__65_right_grid_pin_52_ ;
wire [0:0] cby_1__1__66_ccff_tail ;
wire [0:19] cby_1__1__66_chany_bottom_out ;
wire [0:19] cby_1__1__66_chany_top_out ;
wire [0:0] cby_1__1__66_left_grid_pin_0_ ;
wire [0:0] cby_1__1__66_left_grid_pin_10_ ;
wire [0:0] cby_1__1__66_left_grid_pin_11_ ;
wire [0:0] cby_1__1__66_left_grid_pin_12_ ;
wire [0:0] cby_1__1__66_left_grid_pin_13_ ;
wire [0:0] cby_1__1__66_left_grid_pin_14_ ;
wire [0:0] cby_1__1__66_left_grid_pin_15_ ;
wire [0:0] cby_1__1__66_left_grid_pin_1_ ;
wire [0:0] cby_1__1__66_left_grid_pin_2_ ;
wire [0:0] cby_1__1__66_left_grid_pin_3_ ;
wire [0:0] cby_1__1__66_left_grid_pin_4_ ;
wire [0:0] cby_1__1__66_left_grid_pin_5_ ;
wire [0:0] cby_1__1__66_left_grid_pin_6_ ;
wire [0:0] cby_1__1__66_left_grid_pin_7_ ;
wire [0:0] cby_1__1__66_left_grid_pin_8_ ;
wire [0:0] cby_1__1__66_left_grid_pin_9_ ;
wire [0:0] cby_1__1__66_right_grid_pin_52_ ;
wire [0:0] cby_1__1__67_ccff_tail ;
wire [0:19] cby_1__1__67_chany_bottom_out ;
wire [0:19] cby_1__1__67_chany_top_out ;
wire [0:0] cby_1__1__67_left_grid_pin_0_ ;
wire [0:0] cby_1__1__67_left_grid_pin_10_ ;
wire [0:0] cby_1__1__67_left_grid_pin_11_ ;
wire [0:0] cby_1__1__67_left_grid_pin_12_ ;
wire [0:0] cby_1__1__67_left_grid_pin_13_ ;
wire [0:0] cby_1__1__67_left_grid_pin_14_ ;
wire [0:0] cby_1__1__67_left_grid_pin_15_ ;
wire [0:0] cby_1__1__67_left_grid_pin_1_ ;
wire [0:0] cby_1__1__67_left_grid_pin_2_ ;
wire [0:0] cby_1__1__67_left_grid_pin_3_ ;
wire [0:0] cby_1__1__67_left_grid_pin_4_ ;
wire [0:0] cby_1__1__67_left_grid_pin_5_ ;
wire [0:0] cby_1__1__67_left_grid_pin_6_ ;
wire [0:0] cby_1__1__67_left_grid_pin_7_ ;
wire [0:0] cby_1__1__67_left_grid_pin_8_ ;
wire [0:0] cby_1__1__67_left_grid_pin_9_ ;
wire [0:0] cby_1__1__67_right_grid_pin_52_ ;
wire [0:0] cby_1__1__68_ccff_tail ;
wire [0:19] cby_1__1__68_chany_bottom_out ;
wire [0:19] cby_1__1__68_chany_top_out ;
wire [0:0] cby_1__1__68_left_grid_pin_0_ ;
wire [0:0] cby_1__1__68_left_grid_pin_10_ ;
wire [0:0] cby_1__1__68_left_grid_pin_11_ ;
wire [0:0] cby_1__1__68_left_grid_pin_12_ ;
wire [0:0] cby_1__1__68_left_grid_pin_13_ ;
wire [0:0] cby_1__1__68_left_grid_pin_14_ ;
wire [0:0] cby_1__1__68_left_grid_pin_15_ ;
wire [0:0] cby_1__1__68_left_grid_pin_1_ ;
wire [0:0] cby_1__1__68_left_grid_pin_2_ ;
wire [0:0] cby_1__1__68_left_grid_pin_3_ ;
wire [0:0] cby_1__1__68_left_grid_pin_4_ ;
wire [0:0] cby_1__1__68_left_grid_pin_5_ ;
wire [0:0] cby_1__1__68_left_grid_pin_6_ ;
wire [0:0] cby_1__1__68_left_grid_pin_7_ ;
wire [0:0] cby_1__1__68_left_grid_pin_8_ ;
wire [0:0] cby_1__1__68_left_grid_pin_9_ ;
wire [0:0] cby_1__1__68_right_grid_pin_52_ ;
wire [0:0] cby_1__1__69_ccff_tail ;
wire [0:19] cby_1__1__69_chany_bottom_out ;
wire [0:19] cby_1__1__69_chany_top_out ;
wire [0:0] cby_1__1__69_left_grid_pin_0_ ;
wire [0:0] cby_1__1__69_left_grid_pin_10_ ;
wire [0:0] cby_1__1__69_left_grid_pin_11_ ;
wire [0:0] cby_1__1__69_left_grid_pin_12_ ;
wire [0:0] cby_1__1__69_left_grid_pin_13_ ;
wire [0:0] cby_1__1__69_left_grid_pin_14_ ;
wire [0:0] cby_1__1__69_left_grid_pin_15_ ;
wire [0:0] cby_1__1__69_left_grid_pin_1_ ;
wire [0:0] cby_1__1__69_left_grid_pin_2_ ;
wire [0:0] cby_1__1__69_left_grid_pin_3_ ;
wire [0:0] cby_1__1__69_left_grid_pin_4_ ;
wire [0:0] cby_1__1__69_left_grid_pin_5_ ;
wire [0:0] cby_1__1__69_left_grid_pin_6_ ;
wire [0:0] cby_1__1__69_left_grid_pin_7_ ;
wire [0:0] cby_1__1__69_left_grid_pin_8_ ;
wire [0:0] cby_1__1__69_left_grid_pin_9_ ;
wire [0:0] cby_1__1__69_right_grid_pin_52_ ;
wire [0:0] cby_1__1__6_ccff_tail ;
wire [0:19] cby_1__1__6_chany_bottom_out ;
wire [0:19] cby_1__1__6_chany_top_out ;
wire [0:0] cby_1__1__6_left_grid_pin_0_ ;
wire [0:0] cby_1__1__6_left_grid_pin_10_ ;
wire [0:0] cby_1__1__6_left_grid_pin_11_ ;
wire [0:0] cby_1__1__6_left_grid_pin_12_ ;
wire [0:0] cby_1__1__6_left_grid_pin_13_ ;
wire [0:0] cby_1__1__6_left_grid_pin_14_ ;
wire [0:0] cby_1__1__6_left_grid_pin_15_ ;
wire [0:0] cby_1__1__6_left_grid_pin_1_ ;
wire [0:0] cby_1__1__6_left_grid_pin_2_ ;
wire [0:0] cby_1__1__6_left_grid_pin_3_ ;
wire [0:0] cby_1__1__6_left_grid_pin_4_ ;
wire [0:0] cby_1__1__6_left_grid_pin_5_ ;
wire [0:0] cby_1__1__6_left_grid_pin_6_ ;
wire [0:0] cby_1__1__6_left_grid_pin_7_ ;
wire [0:0] cby_1__1__6_left_grid_pin_8_ ;
wire [0:0] cby_1__1__6_left_grid_pin_9_ ;
wire [0:0] cby_1__1__6_right_grid_pin_52_ ;
wire [0:0] cby_1__1__70_ccff_tail ;
wire [0:19] cby_1__1__70_chany_bottom_out ;
wire [0:19] cby_1__1__70_chany_top_out ;
wire [0:0] cby_1__1__70_left_grid_pin_0_ ;
wire [0:0] cby_1__1__70_left_grid_pin_10_ ;
wire [0:0] cby_1__1__70_left_grid_pin_11_ ;
wire [0:0] cby_1__1__70_left_grid_pin_12_ ;
wire [0:0] cby_1__1__70_left_grid_pin_13_ ;
wire [0:0] cby_1__1__70_left_grid_pin_14_ ;
wire [0:0] cby_1__1__70_left_grid_pin_15_ ;
wire [0:0] cby_1__1__70_left_grid_pin_1_ ;
wire [0:0] cby_1__1__70_left_grid_pin_2_ ;
wire [0:0] cby_1__1__70_left_grid_pin_3_ ;
wire [0:0] cby_1__1__70_left_grid_pin_4_ ;
wire [0:0] cby_1__1__70_left_grid_pin_5_ ;
wire [0:0] cby_1__1__70_left_grid_pin_6_ ;
wire [0:0] cby_1__1__70_left_grid_pin_7_ ;
wire [0:0] cby_1__1__70_left_grid_pin_8_ ;
wire [0:0] cby_1__1__70_left_grid_pin_9_ ;
wire [0:0] cby_1__1__70_right_grid_pin_52_ ;
wire [0:0] cby_1__1__71_ccff_tail ;
wire [0:19] cby_1__1__71_chany_bottom_out ;
wire [0:19] cby_1__1__71_chany_top_out ;
wire [0:0] cby_1__1__71_left_grid_pin_0_ ;
wire [0:0] cby_1__1__71_left_grid_pin_10_ ;
wire [0:0] cby_1__1__71_left_grid_pin_11_ ;
wire [0:0] cby_1__1__71_left_grid_pin_12_ ;
wire [0:0] cby_1__1__71_left_grid_pin_13_ ;
wire [0:0] cby_1__1__71_left_grid_pin_14_ ;
wire [0:0] cby_1__1__71_left_grid_pin_15_ ;
wire [0:0] cby_1__1__71_left_grid_pin_1_ ;
wire [0:0] cby_1__1__71_left_grid_pin_2_ ;
wire [0:0] cby_1__1__71_left_grid_pin_3_ ;
wire [0:0] cby_1__1__71_left_grid_pin_4_ ;
wire [0:0] cby_1__1__71_left_grid_pin_5_ ;
wire [0:0] cby_1__1__71_left_grid_pin_6_ ;
wire [0:0] cby_1__1__71_left_grid_pin_7_ ;
wire [0:0] cby_1__1__71_left_grid_pin_8_ ;
wire [0:0] cby_1__1__71_left_grid_pin_9_ ;
wire [0:0] cby_1__1__71_right_grid_pin_52_ ;
wire [0:0] cby_1__1__72_ccff_tail ;
wire [0:19] cby_1__1__72_chany_bottom_out ;
wire [0:19] cby_1__1__72_chany_top_out ;
wire [0:0] cby_1__1__72_left_grid_pin_0_ ;
wire [0:0] cby_1__1__72_left_grid_pin_10_ ;
wire [0:0] cby_1__1__72_left_grid_pin_11_ ;
wire [0:0] cby_1__1__72_left_grid_pin_12_ ;
wire [0:0] cby_1__1__72_left_grid_pin_13_ ;
wire [0:0] cby_1__1__72_left_grid_pin_14_ ;
wire [0:0] cby_1__1__72_left_grid_pin_15_ ;
wire [0:0] cby_1__1__72_left_grid_pin_1_ ;
wire [0:0] cby_1__1__72_left_grid_pin_2_ ;
wire [0:0] cby_1__1__72_left_grid_pin_3_ ;
wire [0:0] cby_1__1__72_left_grid_pin_4_ ;
wire [0:0] cby_1__1__72_left_grid_pin_5_ ;
wire [0:0] cby_1__1__72_left_grid_pin_6_ ;
wire [0:0] cby_1__1__72_left_grid_pin_7_ ;
wire [0:0] cby_1__1__72_left_grid_pin_8_ ;
wire [0:0] cby_1__1__72_left_grid_pin_9_ ;
wire [0:0] cby_1__1__72_right_grid_pin_52_ ;
wire [0:0] cby_1__1__73_ccff_tail ;
wire [0:19] cby_1__1__73_chany_bottom_out ;
wire [0:19] cby_1__1__73_chany_top_out ;
wire [0:0] cby_1__1__73_left_grid_pin_0_ ;
wire [0:0] cby_1__1__73_left_grid_pin_10_ ;
wire [0:0] cby_1__1__73_left_grid_pin_11_ ;
wire [0:0] cby_1__1__73_left_grid_pin_12_ ;
wire [0:0] cby_1__1__73_left_grid_pin_13_ ;
wire [0:0] cby_1__1__73_left_grid_pin_14_ ;
wire [0:0] cby_1__1__73_left_grid_pin_15_ ;
wire [0:0] cby_1__1__73_left_grid_pin_1_ ;
wire [0:0] cby_1__1__73_left_grid_pin_2_ ;
wire [0:0] cby_1__1__73_left_grid_pin_3_ ;
wire [0:0] cby_1__1__73_left_grid_pin_4_ ;
wire [0:0] cby_1__1__73_left_grid_pin_5_ ;
wire [0:0] cby_1__1__73_left_grid_pin_6_ ;
wire [0:0] cby_1__1__73_left_grid_pin_7_ ;
wire [0:0] cby_1__1__73_left_grid_pin_8_ ;
wire [0:0] cby_1__1__73_left_grid_pin_9_ ;
wire [0:0] cby_1__1__73_right_grid_pin_52_ ;
wire [0:0] cby_1__1__74_ccff_tail ;
wire [0:19] cby_1__1__74_chany_bottom_out ;
wire [0:19] cby_1__1__74_chany_top_out ;
wire [0:0] cby_1__1__74_left_grid_pin_0_ ;
wire [0:0] cby_1__1__74_left_grid_pin_10_ ;
wire [0:0] cby_1__1__74_left_grid_pin_11_ ;
wire [0:0] cby_1__1__74_left_grid_pin_12_ ;
wire [0:0] cby_1__1__74_left_grid_pin_13_ ;
wire [0:0] cby_1__1__74_left_grid_pin_14_ ;
wire [0:0] cby_1__1__74_left_grid_pin_15_ ;
wire [0:0] cby_1__1__74_left_grid_pin_1_ ;
wire [0:0] cby_1__1__74_left_grid_pin_2_ ;
wire [0:0] cby_1__1__74_left_grid_pin_3_ ;
wire [0:0] cby_1__1__74_left_grid_pin_4_ ;
wire [0:0] cby_1__1__74_left_grid_pin_5_ ;
wire [0:0] cby_1__1__74_left_grid_pin_6_ ;
wire [0:0] cby_1__1__74_left_grid_pin_7_ ;
wire [0:0] cby_1__1__74_left_grid_pin_8_ ;
wire [0:0] cby_1__1__74_left_grid_pin_9_ ;
wire [0:0] cby_1__1__74_right_grid_pin_52_ ;
wire [0:0] cby_1__1__75_ccff_tail ;
wire [0:19] cby_1__1__75_chany_bottom_out ;
wire [0:19] cby_1__1__75_chany_top_out ;
wire [0:0] cby_1__1__75_left_grid_pin_0_ ;
wire [0:0] cby_1__1__75_left_grid_pin_10_ ;
wire [0:0] cby_1__1__75_left_grid_pin_11_ ;
wire [0:0] cby_1__1__75_left_grid_pin_12_ ;
wire [0:0] cby_1__1__75_left_grid_pin_13_ ;
wire [0:0] cby_1__1__75_left_grid_pin_14_ ;
wire [0:0] cby_1__1__75_left_grid_pin_15_ ;
wire [0:0] cby_1__1__75_left_grid_pin_1_ ;
wire [0:0] cby_1__1__75_left_grid_pin_2_ ;
wire [0:0] cby_1__1__75_left_grid_pin_3_ ;
wire [0:0] cby_1__1__75_left_grid_pin_4_ ;
wire [0:0] cby_1__1__75_left_grid_pin_5_ ;
wire [0:0] cby_1__1__75_left_grid_pin_6_ ;
wire [0:0] cby_1__1__75_left_grid_pin_7_ ;
wire [0:0] cby_1__1__75_left_grid_pin_8_ ;
wire [0:0] cby_1__1__75_left_grid_pin_9_ ;
wire [0:0] cby_1__1__75_right_grid_pin_52_ ;
wire [0:0] cby_1__1__76_ccff_tail ;
wire [0:19] cby_1__1__76_chany_bottom_out ;
wire [0:19] cby_1__1__76_chany_top_out ;
wire [0:0] cby_1__1__76_left_grid_pin_0_ ;
wire [0:0] cby_1__1__76_left_grid_pin_10_ ;
wire [0:0] cby_1__1__76_left_grid_pin_11_ ;
wire [0:0] cby_1__1__76_left_grid_pin_12_ ;
wire [0:0] cby_1__1__76_left_grid_pin_13_ ;
wire [0:0] cby_1__1__76_left_grid_pin_14_ ;
wire [0:0] cby_1__1__76_left_grid_pin_15_ ;
wire [0:0] cby_1__1__76_left_grid_pin_1_ ;
wire [0:0] cby_1__1__76_left_grid_pin_2_ ;
wire [0:0] cby_1__1__76_left_grid_pin_3_ ;
wire [0:0] cby_1__1__76_left_grid_pin_4_ ;
wire [0:0] cby_1__1__76_left_grid_pin_5_ ;
wire [0:0] cby_1__1__76_left_grid_pin_6_ ;
wire [0:0] cby_1__1__76_left_grid_pin_7_ ;
wire [0:0] cby_1__1__76_left_grid_pin_8_ ;
wire [0:0] cby_1__1__76_left_grid_pin_9_ ;
wire [0:0] cby_1__1__76_right_grid_pin_52_ ;
wire [0:0] cby_1__1__77_ccff_tail ;
wire [0:19] cby_1__1__77_chany_bottom_out ;
wire [0:19] cby_1__1__77_chany_top_out ;
wire [0:0] cby_1__1__77_left_grid_pin_0_ ;
wire [0:0] cby_1__1__77_left_grid_pin_10_ ;
wire [0:0] cby_1__1__77_left_grid_pin_11_ ;
wire [0:0] cby_1__1__77_left_grid_pin_12_ ;
wire [0:0] cby_1__1__77_left_grid_pin_13_ ;
wire [0:0] cby_1__1__77_left_grid_pin_14_ ;
wire [0:0] cby_1__1__77_left_grid_pin_15_ ;
wire [0:0] cby_1__1__77_left_grid_pin_1_ ;
wire [0:0] cby_1__1__77_left_grid_pin_2_ ;
wire [0:0] cby_1__1__77_left_grid_pin_3_ ;
wire [0:0] cby_1__1__77_left_grid_pin_4_ ;
wire [0:0] cby_1__1__77_left_grid_pin_5_ ;
wire [0:0] cby_1__1__77_left_grid_pin_6_ ;
wire [0:0] cby_1__1__77_left_grid_pin_7_ ;
wire [0:0] cby_1__1__77_left_grid_pin_8_ ;
wire [0:0] cby_1__1__77_left_grid_pin_9_ ;
wire [0:0] cby_1__1__77_right_grid_pin_52_ ;
wire [0:0] cby_1__1__78_ccff_tail ;
wire [0:19] cby_1__1__78_chany_bottom_out ;
wire [0:19] cby_1__1__78_chany_top_out ;
wire [0:0] cby_1__1__78_left_grid_pin_0_ ;
wire [0:0] cby_1__1__78_left_grid_pin_10_ ;
wire [0:0] cby_1__1__78_left_grid_pin_11_ ;
wire [0:0] cby_1__1__78_left_grid_pin_12_ ;
wire [0:0] cby_1__1__78_left_grid_pin_13_ ;
wire [0:0] cby_1__1__78_left_grid_pin_14_ ;
wire [0:0] cby_1__1__78_left_grid_pin_15_ ;
wire [0:0] cby_1__1__78_left_grid_pin_1_ ;
wire [0:0] cby_1__1__78_left_grid_pin_2_ ;
wire [0:0] cby_1__1__78_left_grid_pin_3_ ;
wire [0:0] cby_1__1__78_left_grid_pin_4_ ;
wire [0:0] cby_1__1__78_left_grid_pin_5_ ;
wire [0:0] cby_1__1__78_left_grid_pin_6_ ;
wire [0:0] cby_1__1__78_left_grid_pin_7_ ;
wire [0:0] cby_1__1__78_left_grid_pin_8_ ;
wire [0:0] cby_1__1__78_left_grid_pin_9_ ;
wire [0:0] cby_1__1__78_right_grid_pin_52_ ;
wire [0:0] cby_1__1__79_ccff_tail ;
wire [0:19] cby_1__1__79_chany_bottom_out ;
wire [0:19] cby_1__1__79_chany_top_out ;
wire [0:0] cby_1__1__79_left_grid_pin_0_ ;
wire [0:0] cby_1__1__79_left_grid_pin_10_ ;
wire [0:0] cby_1__1__79_left_grid_pin_11_ ;
wire [0:0] cby_1__1__79_left_grid_pin_12_ ;
wire [0:0] cby_1__1__79_left_grid_pin_13_ ;
wire [0:0] cby_1__1__79_left_grid_pin_14_ ;
wire [0:0] cby_1__1__79_left_grid_pin_15_ ;
wire [0:0] cby_1__1__79_left_grid_pin_1_ ;
wire [0:0] cby_1__1__79_left_grid_pin_2_ ;
wire [0:0] cby_1__1__79_left_grid_pin_3_ ;
wire [0:0] cby_1__1__79_left_grid_pin_4_ ;
wire [0:0] cby_1__1__79_left_grid_pin_5_ ;
wire [0:0] cby_1__1__79_left_grid_pin_6_ ;
wire [0:0] cby_1__1__79_left_grid_pin_7_ ;
wire [0:0] cby_1__1__79_left_grid_pin_8_ ;
wire [0:0] cby_1__1__79_left_grid_pin_9_ ;
wire [0:0] cby_1__1__79_right_grid_pin_52_ ;
wire [0:0] cby_1__1__7_ccff_tail ;
wire [0:19] cby_1__1__7_chany_bottom_out ;
wire [0:19] cby_1__1__7_chany_top_out ;
wire [0:0] cby_1__1__7_left_grid_pin_0_ ;
wire [0:0] cby_1__1__7_left_grid_pin_10_ ;
wire [0:0] cby_1__1__7_left_grid_pin_11_ ;
wire [0:0] cby_1__1__7_left_grid_pin_12_ ;
wire [0:0] cby_1__1__7_left_grid_pin_13_ ;
wire [0:0] cby_1__1__7_left_grid_pin_14_ ;
wire [0:0] cby_1__1__7_left_grid_pin_15_ ;
wire [0:0] cby_1__1__7_left_grid_pin_1_ ;
wire [0:0] cby_1__1__7_left_grid_pin_2_ ;
wire [0:0] cby_1__1__7_left_grid_pin_3_ ;
wire [0:0] cby_1__1__7_left_grid_pin_4_ ;
wire [0:0] cby_1__1__7_left_grid_pin_5_ ;
wire [0:0] cby_1__1__7_left_grid_pin_6_ ;
wire [0:0] cby_1__1__7_left_grid_pin_7_ ;
wire [0:0] cby_1__1__7_left_grid_pin_8_ ;
wire [0:0] cby_1__1__7_left_grid_pin_9_ ;
wire [0:0] cby_1__1__7_right_grid_pin_52_ ;
wire [0:0] cby_1__1__80_ccff_tail ;
wire [0:19] cby_1__1__80_chany_bottom_out ;
wire [0:19] cby_1__1__80_chany_top_out ;
wire [0:0] cby_1__1__80_left_grid_pin_0_ ;
wire [0:0] cby_1__1__80_left_grid_pin_10_ ;
wire [0:0] cby_1__1__80_left_grid_pin_11_ ;
wire [0:0] cby_1__1__80_left_grid_pin_12_ ;
wire [0:0] cby_1__1__80_left_grid_pin_13_ ;
wire [0:0] cby_1__1__80_left_grid_pin_14_ ;
wire [0:0] cby_1__1__80_left_grid_pin_15_ ;
wire [0:0] cby_1__1__80_left_grid_pin_1_ ;
wire [0:0] cby_1__1__80_left_grid_pin_2_ ;
wire [0:0] cby_1__1__80_left_grid_pin_3_ ;
wire [0:0] cby_1__1__80_left_grid_pin_4_ ;
wire [0:0] cby_1__1__80_left_grid_pin_5_ ;
wire [0:0] cby_1__1__80_left_grid_pin_6_ ;
wire [0:0] cby_1__1__80_left_grid_pin_7_ ;
wire [0:0] cby_1__1__80_left_grid_pin_8_ ;
wire [0:0] cby_1__1__80_left_grid_pin_9_ ;
wire [0:0] cby_1__1__80_right_grid_pin_52_ ;
wire [0:0] cby_1__1__81_ccff_tail ;
wire [0:19] cby_1__1__81_chany_bottom_out ;
wire [0:19] cby_1__1__81_chany_top_out ;
wire [0:0] cby_1__1__81_left_grid_pin_0_ ;
wire [0:0] cby_1__1__81_left_grid_pin_10_ ;
wire [0:0] cby_1__1__81_left_grid_pin_11_ ;
wire [0:0] cby_1__1__81_left_grid_pin_12_ ;
wire [0:0] cby_1__1__81_left_grid_pin_13_ ;
wire [0:0] cby_1__1__81_left_grid_pin_14_ ;
wire [0:0] cby_1__1__81_left_grid_pin_15_ ;
wire [0:0] cby_1__1__81_left_grid_pin_1_ ;
wire [0:0] cby_1__1__81_left_grid_pin_2_ ;
wire [0:0] cby_1__1__81_left_grid_pin_3_ ;
wire [0:0] cby_1__1__81_left_grid_pin_4_ ;
wire [0:0] cby_1__1__81_left_grid_pin_5_ ;
wire [0:0] cby_1__1__81_left_grid_pin_6_ ;
wire [0:0] cby_1__1__81_left_grid_pin_7_ ;
wire [0:0] cby_1__1__81_left_grid_pin_8_ ;
wire [0:0] cby_1__1__81_left_grid_pin_9_ ;
wire [0:0] cby_1__1__81_right_grid_pin_52_ ;
wire [0:0] cby_1__1__82_ccff_tail ;
wire [0:19] cby_1__1__82_chany_bottom_out ;
wire [0:19] cby_1__1__82_chany_top_out ;
wire [0:0] cby_1__1__82_left_grid_pin_0_ ;
wire [0:0] cby_1__1__82_left_grid_pin_10_ ;
wire [0:0] cby_1__1__82_left_grid_pin_11_ ;
wire [0:0] cby_1__1__82_left_grid_pin_12_ ;
wire [0:0] cby_1__1__82_left_grid_pin_13_ ;
wire [0:0] cby_1__1__82_left_grid_pin_14_ ;
wire [0:0] cby_1__1__82_left_grid_pin_15_ ;
wire [0:0] cby_1__1__82_left_grid_pin_1_ ;
wire [0:0] cby_1__1__82_left_grid_pin_2_ ;
wire [0:0] cby_1__1__82_left_grid_pin_3_ ;
wire [0:0] cby_1__1__82_left_grid_pin_4_ ;
wire [0:0] cby_1__1__82_left_grid_pin_5_ ;
wire [0:0] cby_1__1__82_left_grid_pin_6_ ;
wire [0:0] cby_1__1__82_left_grid_pin_7_ ;
wire [0:0] cby_1__1__82_left_grid_pin_8_ ;
wire [0:0] cby_1__1__82_left_grid_pin_9_ ;
wire [0:0] cby_1__1__82_right_grid_pin_52_ ;
wire [0:0] cby_1__1__83_ccff_tail ;
wire [0:19] cby_1__1__83_chany_bottom_out ;
wire [0:19] cby_1__1__83_chany_top_out ;
wire [0:0] cby_1__1__83_left_grid_pin_0_ ;
wire [0:0] cby_1__1__83_left_grid_pin_10_ ;
wire [0:0] cby_1__1__83_left_grid_pin_11_ ;
wire [0:0] cby_1__1__83_left_grid_pin_12_ ;
wire [0:0] cby_1__1__83_left_grid_pin_13_ ;
wire [0:0] cby_1__1__83_left_grid_pin_14_ ;
wire [0:0] cby_1__1__83_left_grid_pin_15_ ;
wire [0:0] cby_1__1__83_left_grid_pin_1_ ;
wire [0:0] cby_1__1__83_left_grid_pin_2_ ;
wire [0:0] cby_1__1__83_left_grid_pin_3_ ;
wire [0:0] cby_1__1__83_left_grid_pin_4_ ;
wire [0:0] cby_1__1__83_left_grid_pin_5_ ;
wire [0:0] cby_1__1__83_left_grid_pin_6_ ;
wire [0:0] cby_1__1__83_left_grid_pin_7_ ;
wire [0:0] cby_1__1__83_left_grid_pin_8_ ;
wire [0:0] cby_1__1__83_left_grid_pin_9_ ;
wire [0:0] cby_1__1__83_right_grid_pin_52_ ;
wire [0:0] cby_1__1__84_ccff_tail ;
wire [0:19] cby_1__1__84_chany_bottom_out ;
wire [0:19] cby_1__1__84_chany_top_out ;
wire [0:0] cby_1__1__84_left_grid_pin_0_ ;
wire [0:0] cby_1__1__84_left_grid_pin_10_ ;
wire [0:0] cby_1__1__84_left_grid_pin_11_ ;
wire [0:0] cby_1__1__84_left_grid_pin_12_ ;
wire [0:0] cby_1__1__84_left_grid_pin_13_ ;
wire [0:0] cby_1__1__84_left_grid_pin_14_ ;
wire [0:0] cby_1__1__84_left_grid_pin_15_ ;
wire [0:0] cby_1__1__84_left_grid_pin_1_ ;
wire [0:0] cby_1__1__84_left_grid_pin_2_ ;
wire [0:0] cby_1__1__84_left_grid_pin_3_ ;
wire [0:0] cby_1__1__84_left_grid_pin_4_ ;
wire [0:0] cby_1__1__84_left_grid_pin_5_ ;
wire [0:0] cby_1__1__84_left_grid_pin_6_ ;
wire [0:0] cby_1__1__84_left_grid_pin_7_ ;
wire [0:0] cby_1__1__84_left_grid_pin_8_ ;
wire [0:0] cby_1__1__84_left_grid_pin_9_ ;
wire [0:0] cby_1__1__84_right_grid_pin_52_ ;
wire [0:0] cby_1__1__85_ccff_tail ;
wire [0:19] cby_1__1__85_chany_bottom_out ;
wire [0:19] cby_1__1__85_chany_top_out ;
wire [0:0] cby_1__1__85_left_grid_pin_0_ ;
wire [0:0] cby_1__1__85_left_grid_pin_10_ ;
wire [0:0] cby_1__1__85_left_grid_pin_11_ ;
wire [0:0] cby_1__1__85_left_grid_pin_12_ ;
wire [0:0] cby_1__1__85_left_grid_pin_13_ ;
wire [0:0] cby_1__1__85_left_grid_pin_14_ ;
wire [0:0] cby_1__1__85_left_grid_pin_15_ ;
wire [0:0] cby_1__1__85_left_grid_pin_1_ ;
wire [0:0] cby_1__1__85_left_grid_pin_2_ ;
wire [0:0] cby_1__1__85_left_grid_pin_3_ ;
wire [0:0] cby_1__1__85_left_grid_pin_4_ ;
wire [0:0] cby_1__1__85_left_grid_pin_5_ ;
wire [0:0] cby_1__1__85_left_grid_pin_6_ ;
wire [0:0] cby_1__1__85_left_grid_pin_7_ ;
wire [0:0] cby_1__1__85_left_grid_pin_8_ ;
wire [0:0] cby_1__1__85_left_grid_pin_9_ ;
wire [0:0] cby_1__1__85_right_grid_pin_52_ ;
wire [0:0] cby_1__1__86_ccff_tail ;
wire [0:19] cby_1__1__86_chany_bottom_out ;
wire [0:19] cby_1__1__86_chany_top_out ;
wire [0:0] cby_1__1__86_left_grid_pin_0_ ;
wire [0:0] cby_1__1__86_left_grid_pin_10_ ;
wire [0:0] cby_1__1__86_left_grid_pin_11_ ;
wire [0:0] cby_1__1__86_left_grid_pin_12_ ;
wire [0:0] cby_1__1__86_left_grid_pin_13_ ;
wire [0:0] cby_1__1__86_left_grid_pin_14_ ;
wire [0:0] cby_1__1__86_left_grid_pin_15_ ;
wire [0:0] cby_1__1__86_left_grid_pin_1_ ;
wire [0:0] cby_1__1__86_left_grid_pin_2_ ;
wire [0:0] cby_1__1__86_left_grid_pin_3_ ;
wire [0:0] cby_1__1__86_left_grid_pin_4_ ;
wire [0:0] cby_1__1__86_left_grid_pin_5_ ;
wire [0:0] cby_1__1__86_left_grid_pin_6_ ;
wire [0:0] cby_1__1__86_left_grid_pin_7_ ;
wire [0:0] cby_1__1__86_left_grid_pin_8_ ;
wire [0:0] cby_1__1__86_left_grid_pin_9_ ;
wire [0:0] cby_1__1__86_right_grid_pin_52_ ;
wire [0:0] cby_1__1__87_ccff_tail ;
wire [0:19] cby_1__1__87_chany_bottom_out ;
wire [0:19] cby_1__1__87_chany_top_out ;
wire [0:0] cby_1__1__87_left_grid_pin_0_ ;
wire [0:0] cby_1__1__87_left_grid_pin_10_ ;
wire [0:0] cby_1__1__87_left_grid_pin_11_ ;
wire [0:0] cby_1__1__87_left_grid_pin_12_ ;
wire [0:0] cby_1__1__87_left_grid_pin_13_ ;
wire [0:0] cby_1__1__87_left_grid_pin_14_ ;
wire [0:0] cby_1__1__87_left_grid_pin_15_ ;
wire [0:0] cby_1__1__87_left_grid_pin_1_ ;
wire [0:0] cby_1__1__87_left_grid_pin_2_ ;
wire [0:0] cby_1__1__87_left_grid_pin_3_ ;
wire [0:0] cby_1__1__87_left_grid_pin_4_ ;
wire [0:0] cby_1__1__87_left_grid_pin_5_ ;
wire [0:0] cby_1__1__87_left_grid_pin_6_ ;
wire [0:0] cby_1__1__87_left_grid_pin_7_ ;
wire [0:0] cby_1__1__87_left_grid_pin_8_ ;
wire [0:0] cby_1__1__87_left_grid_pin_9_ ;
wire [0:0] cby_1__1__87_right_grid_pin_52_ ;
wire [0:0] cby_1__1__88_ccff_tail ;
wire [0:19] cby_1__1__88_chany_bottom_out ;
wire [0:19] cby_1__1__88_chany_top_out ;
wire [0:0] cby_1__1__88_left_grid_pin_0_ ;
wire [0:0] cby_1__1__88_left_grid_pin_10_ ;
wire [0:0] cby_1__1__88_left_grid_pin_11_ ;
wire [0:0] cby_1__1__88_left_grid_pin_12_ ;
wire [0:0] cby_1__1__88_left_grid_pin_13_ ;
wire [0:0] cby_1__1__88_left_grid_pin_14_ ;
wire [0:0] cby_1__1__88_left_grid_pin_15_ ;
wire [0:0] cby_1__1__88_left_grid_pin_1_ ;
wire [0:0] cby_1__1__88_left_grid_pin_2_ ;
wire [0:0] cby_1__1__88_left_grid_pin_3_ ;
wire [0:0] cby_1__1__88_left_grid_pin_4_ ;
wire [0:0] cby_1__1__88_left_grid_pin_5_ ;
wire [0:0] cby_1__1__88_left_grid_pin_6_ ;
wire [0:0] cby_1__1__88_left_grid_pin_7_ ;
wire [0:0] cby_1__1__88_left_grid_pin_8_ ;
wire [0:0] cby_1__1__88_left_grid_pin_9_ ;
wire [0:0] cby_1__1__88_right_grid_pin_52_ ;
wire [0:0] cby_1__1__89_ccff_tail ;
wire [0:19] cby_1__1__89_chany_bottom_out ;
wire [0:19] cby_1__1__89_chany_top_out ;
wire [0:0] cby_1__1__89_left_grid_pin_0_ ;
wire [0:0] cby_1__1__89_left_grid_pin_10_ ;
wire [0:0] cby_1__1__89_left_grid_pin_11_ ;
wire [0:0] cby_1__1__89_left_grid_pin_12_ ;
wire [0:0] cby_1__1__89_left_grid_pin_13_ ;
wire [0:0] cby_1__1__89_left_grid_pin_14_ ;
wire [0:0] cby_1__1__89_left_grid_pin_15_ ;
wire [0:0] cby_1__1__89_left_grid_pin_1_ ;
wire [0:0] cby_1__1__89_left_grid_pin_2_ ;
wire [0:0] cby_1__1__89_left_grid_pin_3_ ;
wire [0:0] cby_1__1__89_left_grid_pin_4_ ;
wire [0:0] cby_1__1__89_left_grid_pin_5_ ;
wire [0:0] cby_1__1__89_left_grid_pin_6_ ;
wire [0:0] cby_1__1__89_left_grid_pin_7_ ;
wire [0:0] cby_1__1__89_left_grid_pin_8_ ;
wire [0:0] cby_1__1__89_left_grid_pin_9_ ;
wire [0:0] cby_1__1__89_right_grid_pin_52_ ;
wire [0:0] cby_1__1__8_ccff_tail ;
wire [0:19] cby_1__1__8_chany_bottom_out ;
wire [0:19] cby_1__1__8_chany_top_out ;
wire [0:0] cby_1__1__8_left_grid_pin_0_ ;
wire [0:0] cby_1__1__8_left_grid_pin_10_ ;
wire [0:0] cby_1__1__8_left_grid_pin_11_ ;
wire [0:0] cby_1__1__8_left_grid_pin_12_ ;
wire [0:0] cby_1__1__8_left_grid_pin_13_ ;
wire [0:0] cby_1__1__8_left_grid_pin_14_ ;
wire [0:0] cby_1__1__8_left_grid_pin_15_ ;
wire [0:0] cby_1__1__8_left_grid_pin_1_ ;
wire [0:0] cby_1__1__8_left_grid_pin_2_ ;
wire [0:0] cby_1__1__8_left_grid_pin_3_ ;
wire [0:0] cby_1__1__8_left_grid_pin_4_ ;
wire [0:0] cby_1__1__8_left_grid_pin_5_ ;
wire [0:0] cby_1__1__8_left_grid_pin_6_ ;
wire [0:0] cby_1__1__8_left_grid_pin_7_ ;
wire [0:0] cby_1__1__8_left_grid_pin_8_ ;
wire [0:0] cby_1__1__8_left_grid_pin_9_ ;
wire [0:0] cby_1__1__8_right_grid_pin_52_ ;
wire [0:0] cby_1__1__90_ccff_tail ;
wire [0:19] cby_1__1__90_chany_bottom_out ;
wire [0:19] cby_1__1__90_chany_top_out ;
wire [0:0] cby_1__1__90_left_grid_pin_0_ ;
wire [0:0] cby_1__1__90_left_grid_pin_10_ ;
wire [0:0] cby_1__1__90_left_grid_pin_11_ ;
wire [0:0] cby_1__1__90_left_grid_pin_12_ ;
wire [0:0] cby_1__1__90_left_grid_pin_13_ ;
wire [0:0] cby_1__1__90_left_grid_pin_14_ ;
wire [0:0] cby_1__1__90_left_grid_pin_15_ ;
wire [0:0] cby_1__1__90_left_grid_pin_1_ ;
wire [0:0] cby_1__1__90_left_grid_pin_2_ ;
wire [0:0] cby_1__1__90_left_grid_pin_3_ ;
wire [0:0] cby_1__1__90_left_grid_pin_4_ ;
wire [0:0] cby_1__1__90_left_grid_pin_5_ ;
wire [0:0] cby_1__1__90_left_grid_pin_6_ ;
wire [0:0] cby_1__1__90_left_grid_pin_7_ ;
wire [0:0] cby_1__1__90_left_grid_pin_8_ ;
wire [0:0] cby_1__1__90_left_grid_pin_9_ ;
wire [0:0] cby_1__1__90_right_grid_pin_52_ ;
wire [0:0] cby_1__1__91_ccff_tail ;
wire [0:19] cby_1__1__91_chany_bottom_out ;
wire [0:19] cby_1__1__91_chany_top_out ;
wire [0:0] cby_1__1__91_left_grid_pin_0_ ;
wire [0:0] cby_1__1__91_left_grid_pin_10_ ;
wire [0:0] cby_1__1__91_left_grid_pin_11_ ;
wire [0:0] cby_1__1__91_left_grid_pin_12_ ;
wire [0:0] cby_1__1__91_left_grid_pin_13_ ;
wire [0:0] cby_1__1__91_left_grid_pin_14_ ;
wire [0:0] cby_1__1__91_left_grid_pin_15_ ;
wire [0:0] cby_1__1__91_left_grid_pin_1_ ;
wire [0:0] cby_1__1__91_left_grid_pin_2_ ;
wire [0:0] cby_1__1__91_left_grid_pin_3_ ;
wire [0:0] cby_1__1__91_left_grid_pin_4_ ;
wire [0:0] cby_1__1__91_left_grid_pin_5_ ;
wire [0:0] cby_1__1__91_left_grid_pin_6_ ;
wire [0:0] cby_1__1__91_left_grid_pin_7_ ;
wire [0:0] cby_1__1__91_left_grid_pin_8_ ;
wire [0:0] cby_1__1__91_left_grid_pin_9_ ;
wire [0:0] cby_1__1__91_right_grid_pin_52_ ;
wire [0:0] cby_1__1__92_ccff_tail ;
wire [0:19] cby_1__1__92_chany_bottom_out ;
wire [0:19] cby_1__1__92_chany_top_out ;
wire [0:0] cby_1__1__92_left_grid_pin_0_ ;
wire [0:0] cby_1__1__92_left_grid_pin_10_ ;
wire [0:0] cby_1__1__92_left_grid_pin_11_ ;
wire [0:0] cby_1__1__92_left_grid_pin_12_ ;
wire [0:0] cby_1__1__92_left_grid_pin_13_ ;
wire [0:0] cby_1__1__92_left_grid_pin_14_ ;
wire [0:0] cby_1__1__92_left_grid_pin_15_ ;
wire [0:0] cby_1__1__92_left_grid_pin_1_ ;
wire [0:0] cby_1__1__92_left_grid_pin_2_ ;
wire [0:0] cby_1__1__92_left_grid_pin_3_ ;
wire [0:0] cby_1__1__92_left_grid_pin_4_ ;
wire [0:0] cby_1__1__92_left_grid_pin_5_ ;
wire [0:0] cby_1__1__92_left_grid_pin_6_ ;
wire [0:0] cby_1__1__92_left_grid_pin_7_ ;
wire [0:0] cby_1__1__92_left_grid_pin_8_ ;
wire [0:0] cby_1__1__92_left_grid_pin_9_ ;
wire [0:0] cby_1__1__92_right_grid_pin_52_ ;
wire [0:0] cby_1__1__93_ccff_tail ;
wire [0:19] cby_1__1__93_chany_bottom_out ;
wire [0:19] cby_1__1__93_chany_top_out ;
wire [0:0] cby_1__1__93_left_grid_pin_0_ ;
wire [0:0] cby_1__1__93_left_grid_pin_10_ ;
wire [0:0] cby_1__1__93_left_grid_pin_11_ ;
wire [0:0] cby_1__1__93_left_grid_pin_12_ ;
wire [0:0] cby_1__1__93_left_grid_pin_13_ ;
wire [0:0] cby_1__1__93_left_grid_pin_14_ ;
wire [0:0] cby_1__1__93_left_grid_pin_15_ ;
wire [0:0] cby_1__1__93_left_grid_pin_1_ ;
wire [0:0] cby_1__1__93_left_grid_pin_2_ ;
wire [0:0] cby_1__1__93_left_grid_pin_3_ ;
wire [0:0] cby_1__1__93_left_grid_pin_4_ ;
wire [0:0] cby_1__1__93_left_grid_pin_5_ ;
wire [0:0] cby_1__1__93_left_grid_pin_6_ ;
wire [0:0] cby_1__1__93_left_grid_pin_7_ ;
wire [0:0] cby_1__1__93_left_grid_pin_8_ ;
wire [0:0] cby_1__1__93_left_grid_pin_9_ ;
wire [0:0] cby_1__1__93_right_grid_pin_52_ ;
wire [0:0] cby_1__1__94_ccff_tail ;
wire [0:19] cby_1__1__94_chany_bottom_out ;
wire [0:19] cby_1__1__94_chany_top_out ;
wire [0:0] cby_1__1__94_left_grid_pin_0_ ;
wire [0:0] cby_1__1__94_left_grid_pin_10_ ;
wire [0:0] cby_1__1__94_left_grid_pin_11_ ;
wire [0:0] cby_1__1__94_left_grid_pin_12_ ;
wire [0:0] cby_1__1__94_left_grid_pin_13_ ;
wire [0:0] cby_1__1__94_left_grid_pin_14_ ;
wire [0:0] cby_1__1__94_left_grid_pin_15_ ;
wire [0:0] cby_1__1__94_left_grid_pin_1_ ;
wire [0:0] cby_1__1__94_left_grid_pin_2_ ;
wire [0:0] cby_1__1__94_left_grid_pin_3_ ;
wire [0:0] cby_1__1__94_left_grid_pin_4_ ;
wire [0:0] cby_1__1__94_left_grid_pin_5_ ;
wire [0:0] cby_1__1__94_left_grid_pin_6_ ;
wire [0:0] cby_1__1__94_left_grid_pin_7_ ;
wire [0:0] cby_1__1__94_left_grid_pin_8_ ;
wire [0:0] cby_1__1__94_left_grid_pin_9_ ;
wire [0:0] cby_1__1__94_right_grid_pin_52_ ;
wire [0:0] cby_1__1__95_ccff_tail ;
wire [0:19] cby_1__1__95_chany_bottom_out ;
wire [0:19] cby_1__1__95_chany_top_out ;
wire [0:0] cby_1__1__95_left_grid_pin_0_ ;
wire [0:0] cby_1__1__95_left_grid_pin_10_ ;
wire [0:0] cby_1__1__95_left_grid_pin_11_ ;
wire [0:0] cby_1__1__95_left_grid_pin_12_ ;
wire [0:0] cby_1__1__95_left_grid_pin_13_ ;
wire [0:0] cby_1__1__95_left_grid_pin_14_ ;
wire [0:0] cby_1__1__95_left_grid_pin_15_ ;
wire [0:0] cby_1__1__95_left_grid_pin_1_ ;
wire [0:0] cby_1__1__95_left_grid_pin_2_ ;
wire [0:0] cby_1__1__95_left_grid_pin_3_ ;
wire [0:0] cby_1__1__95_left_grid_pin_4_ ;
wire [0:0] cby_1__1__95_left_grid_pin_5_ ;
wire [0:0] cby_1__1__95_left_grid_pin_6_ ;
wire [0:0] cby_1__1__95_left_grid_pin_7_ ;
wire [0:0] cby_1__1__95_left_grid_pin_8_ ;
wire [0:0] cby_1__1__95_left_grid_pin_9_ ;
wire [0:0] cby_1__1__95_right_grid_pin_52_ ;
wire [0:0] cby_1__1__96_ccff_tail ;
wire [0:19] cby_1__1__96_chany_bottom_out ;
wire [0:19] cby_1__1__96_chany_top_out ;
wire [0:0] cby_1__1__96_left_grid_pin_0_ ;
wire [0:0] cby_1__1__96_left_grid_pin_10_ ;
wire [0:0] cby_1__1__96_left_grid_pin_11_ ;
wire [0:0] cby_1__1__96_left_grid_pin_12_ ;
wire [0:0] cby_1__1__96_left_grid_pin_13_ ;
wire [0:0] cby_1__1__96_left_grid_pin_14_ ;
wire [0:0] cby_1__1__96_left_grid_pin_15_ ;
wire [0:0] cby_1__1__96_left_grid_pin_1_ ;
wire [0:0] cby_1__1__96_left_grid_pin_2_ ;
wire [0:0] cby_1__1__96_left_grid_pin_3_ ;
wire [0:0] cby_1__1__96_left_grid_pin_4_ ;
wire [0:0] cby_1__1__96_left_grid_pin_5_ ;
wire [0:0] cby_1__1__96_left_grid_pin_6_ ;
wire [0:0] cby_1__1__96_left_grid_pin_7_ ;
wire [0:0] cby_1__1__96_left_grid_pin_8_ ;
wire [0:0] cby_1__1__96_left_grid_pin_9_ ;
wire [0:0] cby_1__1__96_right_grid_pin_52_ ;
wire [0:0] cby_1__1__97_ccff_tail ;
wire [0:19] cby_1__1__97_chany_bottom_out ;
wire [0:19] cby_1__1__97_chany_top_out ;
wire [0:0] cby_1__1__97_left_grid_pin_0_ ;
wire [0:0] cby_1__1__97_left_grid_pin_10_ ;
wire [0:0] cby_1__1__97_left_grid_pin_11_ ;
wire [0:0] cby_1__1__97_left_grid_pin_12_ ;
wire [0:0] cby_1__1__97_left_grid_pin_13_ ;
wire [0:0] cby_1__1__97_left_grid_pin_14_ ;
wire [0:0] cby_1__1__97_left_grid_pin_15_ ;
wire [0:0] cby_1__1__97_left_grid_pin_1_ ;
wire [0:0] cby_1__1__97_left_grid_pin_2_ ;
wire [0:0] cby_1__1__97_left_grid_pin_3_ ;
wire [0:0] cby_1__1__97_left_grid_pin_4_ ;
wire [0:0] cby_1__1__97_left_grid_pin_5_ ;
wire [0:0] cby_1__1__97_left_grid_pin_6_ ;
wire [0:0] cby_1__1__97_left_grid_pin_7_ ;
wire [0:0] cby_1__1__97_left_grid_pin_8_ ;
wire [0:0] cby_1__1__97_left_grid_pin_9_ ;
wire [0:0] cby_1__1__97_right_grid_pin_52_ ;
wire [0:0] cby_1__1__98_ccff_tail ;
wire [0:19] cby_1__1__98_chany_bottom_out ;
wire [0:19] cby_1__1__98_chany_top_out ;
wire [0:0] cby_1__1__98_left_grid_pin_0_ ;
wire [0:0] cby_1__1__98_left_grid_pin_10_ ;
wire [0:0] cby_1__1__98_left_grid_pin_11_ ;
wire [0:0] cby_1__1__98_left_grid_pin_12_ ;
wire [0:0] cby_1__1__98_left_grid_pin_13_ ;
wire [0:0] cby_1__1__98_left_grid_pin_14_ ;
wire [0:0] cby_1__1__98_left_grid_pin_15_ ;
wire [0:0] cby_1__1__98_left_grid_pin_1_ ;
wire [0:0] cby_1__1__98_left_grid_pin_2_ ;
wire [0:0] cby_1__1__98_left_grid_pin_3_ ;
wire [0:0] cby_1__1__98_left_grid_pin_4_ ;
wire [0:0] cby_1__1__98_left_grid_pin_5_ ;
wire [0:0] cby_1__1__98_left_grid_pin_6_ ;
wire [0:0] cby_1__1__98_left_grid_pin_7_ ;
wire [0:0] cby_1__1__98_left_grid_pin_8_ ;
wire [0:0] cby_1__1__98_left_grid_pin_9_ ;
wire [0:0] cby_1__1__98_right_grid_pin_52_ ;
wire [0:0] cby_1__1__99_ccff_tail ;
wire [0:19] cby_1__1__99_chany_bottom_out ;
wire [0:19] cby_1__1__99_chany_top_out ;
wire [0:0] cby_1__1__99_left_grid_pin_0_ ;
wire [0:0] cby_1__1__99_left_grid_pin_10_ ;
wire [0:0] cby_1__1__99_left_grid_pin_11_ ;
wire [0:0] cby_1__1__99_left_grid_pin_12_ ;
wire [0:0] cby_1__1__99_left_grid_pin_13_ ;
wire [0:0] cby_1__1__99_left_grid_pin_14_ ;
wire [0:0] cby_1__1__99_left_grid_pin_15_ ;
wire [0:0] cby_1__1__99_left_grid_pin_1_ ;
wire [0:0] cby_1__1__99_left_grid_pin_2_ ;
wire [0:0] cby_1__1__99_left_grid_pin_3_ ;
wire [0:0] cby_1__1__99_left_grid_pin_4_ ;
wire [0:0] cby_1__1__99_left_grid_pin_5_ ;
wire [0:0] cby_1__1__99_left_grid_pin_6_ ;
wire [0:0] cby_1__1__99_left_grid_pin_7_ ;
wire [0:0] cby_1__1__99_left_grid_pin_8_ ;
wire [0:0] cby_1__1__99_left_grid_pin_9_ ;
wire [0:0] cby_1__1__99_right_grid_pin_52_ ;
wire [0:0] cby_1__1__9_ccff_tail ;
wire [0:19] cby_1__1__9_chany_bottom_out ;
wire [0:19] cby_1__1__9_chany_top_out ;
wire [0:0] cby_1__1__9_left_grid_pin_0_ ;
wire [0:0] cby_1__1__9_left_grid_pin_10_ ;
wire [0:0] cby_1__1__9_left_grid_pin_11_ ;
wire [0:0] cby_1__1__9_left_grid_pin_12_ ;
wire [0:0] cby_1__1__9_left_grid_pin_13_ ;
wire [0:0] cby_1__1__9_left_grid_pin_14_ ;
wire [0:0] cby_1__1__9_left_grid_pin_15_ ;
wire [0:0] cby_1__1__9_left_grid_pin_1_ ;
wire [0:0] cby_1__1__9_left_grid_pin_2_ ;
wire [0:0] cby_1__1__9_left_grid_pin_3_ ;
wire [0:0] cby_1__1__9_left_grid_pin_4_ ;
wire [0:0] cby_1__1__9_left_grid_pin_5_ ;
wire [0:0] cby_1__1__9_left_grid_pin_6_ ;
wire [0:0] cby_1__1__9_left_grid_pin_7_ ;
wire [0:0] cby_1__1__9_left_grid_pin_8_ ;
wire [0:0] cby_1__1__9_left_grid_pin_9_ ;
wire [0:0] cby_1__1__9_right_grid_pin_52_ ;
wire [0:0] direct_interc_0_out ;
wire [0:0] direct_interc_100_out ;
wire [0:0] direct_interc_101_out ;
wire [0:0] direct_interc_102_out ;
wire [0:0] direct_interc_103_out ;
wire [0:0] direct_interc_104_out ;
wire [0:0] direct_interc_105_out ;
wire [0:0] direct_interc_106_out ;
wire [0:0] direct_interc_107_out ;
wire [0:0] direct_interc_108_out ;
wire [0:0] direct_interc_109_out ;
wire [0:0] direct_interc_10_out ;
wire [0:0] direct_interc_110_out ;
wire [0:0] direct_interc_111_out ;
wire [0:0] direct_interc_112_out ;
wire [0:0] direct_interc_113_out ;
wire [0:0] direct_interc_114_out ;
wire [0:0] direct_interc_115_out ;
wire [0:0] direct_interc_116_out ;
wire [0:0] direct_interc_117_out ;
wire [0:0] direct_interc_118_out ;
wire [0:0] direct_interc_119_out ;
wire [0:0] direct_interc_11_out ;
wire [0:0] direct_interc_120_out ;
wire [0:0] direct_interc_121_out ;
wire [0:0] direct_interc_122_out ;
wire [0:0] direct_interc_123_out ;
wire [0:0] direct_interc_124_out ;
wire [0:0] direct_interc_125_out ;
wire [0:0] direct_interc_126_out ;
wire [0:0] direct_interc_127_out ;
wire [0:0] direct_interc_128_out ;
wire [0:0] direct_interc_129_out ;
wire [0:0] direct_interc_12_out ;
wire [0:0] direct_interc_130_out ;
wire [0:0] direct_interc_131_out ;
wire [0:0] direct_interc_132_out ;
wire [0:0] direct_interc_133_out ;
wire [0:0] direct_interc_134_out ;
wire [0:0] direct_interc_135_out ;
wire [0:0] direct_interc_136_out ;
wire [0:0] direct_interc_137_out ;
wire [0:0] direct_interc_138_out ;
wire [0:0] direct_interc_139_out ;
wire [0:0] direct_interc_13_out ;
wire [0:0] direct_interc_140_out ;
wire [0:0] direct_interc_141_out ;
wire [0:0] direct_interc_142_out ;
wire [0:0] direct_interc_143_out ;
wire [0:0] direct_interc_144_out ;
wire [0:0] direct_interc_145_out ;
wire [0:0] direct_interc_146_out ;
wire [0:0] direct_interc_147_out ;
wire [0:0] direct_interc_148_out ;
wire [0:0] direct_interc_149_out ;
wire [0:0] direct_interc_14_out ;
wire [0:0] direct_interc_150_out ;
wire [0:0] direct_interc_151_out ;
wire [0:0] direct_interc_152_out ;
wire [0:0] direct_interc_153_out ;
wire [0:0] direct_interc_154_out ;
wire [0:0] direct_interc_155_out ;
wire [0:0] direct_interc_156_out ;
wire [0:0] direct_interc_157_out ;
wire [0:0] direct_interc_158_out ;
wire [0:0] direct_interc_159_out ;
wire [0:0] direct_interc_15_out ;
wire [0:0] direct_interc_160_out ;
wire [0:0] direct_interc_161_out ;
wire [0:0] direct_interc_162_out ;
wire [0:0] direct_interc_163_out ;
wire [0:0] direct_interc_164_out ;
wire [0:0] direct_interc_165_out ;
wire [0:0] direct_interc_166_out ;
wire [0:0] direct_interc_167_out ;
wire [0:0] direct_interc_168_out ;
wire [0:0] direct_interc_169_out ;
wire [0:0] direct_interc_16_out ;
wire [0:0] direct_interc_170_out ;
wire [0:0] direct_interc_171_out ;
wire [0:0] direct_interc_172_out ;
wire [0:0] direct_interc_173_out ;
wire [0:0] direct_interc_174_out ;
wire [0:0] direct_interc_175_out ;
wire [0:0] direct_interc_176_out ;
wire [0:0] direct_interc_177_out ;
wire [0:0] direct_interc_178_out ;
wire [0:0] direct_interc_179_out ;
wire [0:0] direct_interc_17_out ;
wire [0:0] direct_interc_180_out ;
wire [0:0] direct_interc_181_out ;
wire [0:0] direct_interc_182_out ;
wire [0:0] direct_interc_183_out ;
wire [0:0] direct_interc_184_out ;
wire [0:0] direct_interc_185_out ;
wire [0:0] direct_interc_186_out ;
wire [0:0] direct_interc_187_out ;
wire [0:0] direct_interc_188_out ;
wire [0:0] direct_interc_189_out ;
wire [0:0] direct_interc_18_out ;
wire [0:0] direct_interc_190_out ;
wire [0:0] direct_interc_191_out ;
wire [0:0] direct_interc_192_out ;
wire [0:0] direct_interc_193_out ;
wire [0:0] direct_interc_194_out ;
wire [0:0] direct_interc_195_out ;
wire [0:0] direct_interc_196_out ;
wire [0:0] direct_interc_197_out ;
wire [0:0] direct_interc_198_out ;
wire [0:0] direct_interc_199_out ;
wire [0:0] direct_interc_19_out ;
wire [0:0] direct_interc_1_out ;
wire [0:0] direct_interc_200_out ;
wire [0:0] direct_interc_201_out ;
wire [0:0] direct_interc_202_out ;
wire [0:0] direct_interc_203_out ;
wire [0:0] direct_interc_204_out ;
wire [0:0] direct_interc_205_out ;
wire [0:0] direct_interc_206_out ;
wire [0:0] direct_interc_207_out ;
wire [0:0] direct_interc_208_out ;
wire [0:0] direct_interc_209_out ;
wire [0:0] direct_interc_20_out ;
wire [0:0] direct_interc_210_out ;
wire [0:0] direct_interc_211_out ;
wire [0:0] direct_interc_212_out ;
wire [0:0] direct_interc_213_out ;
wire [0:0] direct_interc_214_out ;
wire [0:0] direct_interc_215_out ;
wire [0:0] direct_interc_216_out ;
wire [0:0] direct_interc_217_out ;
wire [0:0] direct_interc_218_out ;
wire [0:0] direct_interc_219_out ;
wire [0:0] direct_interc_21_out ;
wire [0:0] direct_interc_220_out ;
wire [0:0] direct_interc_221_out ;
wire [0:0] direct_interc_222_out ;
wire [0:0] direct_interc_223_out ;
wire [0:0] direct_interc_224_out ;
wire [0:0] direct_interc_225_out ;
wire [0:0] direct_interc_226_out ;
wire [0:0] direct_interc_227_out ;
wire [0:0] direct_interc_228_out ;
wire [0:0] direct_interc_229_out ;
wire [0:0] direct_interc_22_out ;
wire [0:0] direct_interc_230_out ;
wire [0:0] direct_interc_231_out ;
wire [0:0] direct_interc_232_out ;
wire [0:0] direct_interc_233_out ;
wire [0:0] direct_interc_234_out ;
wire [0:0] direct_interc_235_out ;
wire [0:0] direct_interc_236_out ;
wire [0:0] direct_interc_237_out ;
wire [0:0] direct_interc_238_out ;
wire [0:0] direct_interc_239_out ;
wire [0:0] direct_interc_23_out ;
wire [0:0] direct_interc_240_out ;
wire [0:0] direct_interc_241_out ;
wire [0:0] direct_interc_242_out ;
wire [0:0] direct_interc_243_out ;
wire [0:0] direct_interc_244_out ;
wire [0:0] direct_interc_245_out ;
wire [0:0] direct_interc_246_out ;
wire [0:0] direct_interc_247_out ;
wire [0:0] direct_interc_248_out ;
wire [0:0] direct_interc_249_out ;
wire [0:0] direct_interc_24_out ;
wire [0:0] direct_interc_250_out ;
wire [0:0] direct_interc_251_out ;
wire [0:0] direct_interc_252_out ;
wire [0:0] direct_interc_253_out ;
wire [0:0] direct_interc_254_out ;
wire [0:0] direct_interc_255_out ;
wire [0:0] direct_interc_256_out ;
wire [0:0] direct_interc_257_out ;
wire [0:0] direct_interc_258_out ;
wire [0:0] direct_interc_259_out ;
wire [0:0] direct_interc_25_out ;
wire [0:0] direct_interc_260_out ;
wire [0:0] direct_interc_261_out ;
wire [0:0] direct_interc_262_out ;
wire [0:0] direct_interc_263_out ;
wire [0:0] direct_interc_264_out ;
wire [0:0] direct_interc_265_out ;
wire [0:0] direct_interc_266_out ;
wire [0:0] direct_interc_267_out ;
wire [0:0] direct_interc_268_out ;
wire [0:0] direct_interc_269_out ;
wire [0:0] direct_interc_26_out ;
wire [0:0] direct_interc_270_out ;
wire [0:0] direct_interc_271_out ;
wire [0:0] direct_interc_272_out ;
wire [0:0] direct_interc_273_out ;
wire [0:0] direct_interc_274_out ;
wire [0:0] direct_interc_275_out ;
wire [0:0] direct_interc_276_out ;
wire [0:0] direct_interc_277_out ;
wire [0:0] direct_interc_278_out ;
wire [0:0] direct_interc_279_out ;
wire [0:0] direct_interc_27_out ;
wire [0:0] direct_interc_280_out ;
wire [0:0] direct_interc_281_out ;
wire [0:0] direct_interc_282_out ;
wire [0:0] direct_interc_283_out ;
wire [0:0] direct_interc_284_out ;
wire [0:0] direct_interc_285_out ;
wire [0:0] direct_interc_28_out ;
wire [0:0] direct_interc_29_out ;
wire [0:0] direct_interc_2_out ;
wire [0:0] direct_interc_30_out ;
wire [0:0] direct_interc_31_out ;
wire [0:0] direct_interc_32_out ;
wire [0:0] direct_interc_33_out ;
wire [0:0] direct_interc_34_out ;
wire [0:0] direct_interc_35_out ;
wire [0:0] direct_interc_36_out ;
wire [0:0] direct_interc_37_out ;
wire [0:0] direct_interc_38_out ;
wire [0:0] direct_interc_39_out ;
wire [0:0] direct_interc_3_out ;
wire [0:0] direct_interc_40_out ;
wire [0:0] direct_interc_41_out ;
wire [0:0] direct_interc_42_out ;
wire [0:0] direct_interc_43_out ;
wire [0:0] direct_interc_44_out ;
wire [0:0] direct_interc_45_out ;
wire [0:0] direct_interc_46_out ;
wire [0:0] direct_interc_47_out ;
wire [0:0] direct_interc_48_out ;
wire [0:0] direct_interc_49_out ;
wire [0:0] direct_interc_4_out ;
wire [0:0] direct_interc_50_out ;
wire [0:0] direct_interc_51_out ;
wire [0:0] direct_interc_52_out ;
wire [0:0] direct_interc_53_out ;
wire [0:0] direct_interc_54_out ;
wire [0:0] direct_interc_55_out ;
wire [0:0] direct_interc_56_out ;
wire [0:0] direct_interc_57_out ;
wire [0:0] direct_interc_58_out ;
wire [0:0] direct_interc_59_out ;
wire [0:0] direct_interc_5_out ;
wire [0:0] direct_interc_60_out ;
wire [0:0] direct_interc_61_out ;
wire [0:0] direct_interc_62_out ;
wire [0:0] direct_interc_63_out ;
wire [0:0] direct_interc_64_out ;
wire [0:0] direct_interc_65_out ;
wire [0:0] direct_interc_66_out ;
wire [0:0] direct_interc_67_out ;
wire [0:0] direct_interc_68_out ;
wire [0:0] direct_interc_69_out ;
wire [0:0] direct_interc_6_out ;
wire [0:0] direct_interc_70_out ;
wire [0:0] direct_interc_71_out ;
wire [0:0] direct_interc_72_out ;
wire [0:0] direct_interc_73_out ;
wire [0:0] direct_interc_74_out ;
wire [0:0] direct_interc_75_out ;
wire [0:0] direct_interc_76_out ;
wire [0:0] direct_interc_77_out ;
wire [0:0] direct_interc_78_out ;
wire [0:0] direct_interc_79_out ;
wire [0:0] direct_interc_7_out ;
wire [0:0] direct_interc_80_out ;
wire [0:0] direct_interc_81_out ;
wire [0:0] direct_interc_82_out ;
wire [0:0] direct_interc_83_out ;
wire [0:0] direct_interc_84_out ;
wire [0:0] direct_interc_85_out ;
wire [0:0] direct_interc_86_out ;
wire [0:0] direct_interc_87_out ;
wire [0:0] direct_interc_88_out ;
wire [0:0] direct_interc_89_out ;
wire [0:0] direct_interc_8_out ;
wire [0:0] direct_interc_90_out ;
wire [0:0] direct_interc_91_out ;
wire [0:0] direct_interc_92_out ;
wire [0:0] direct_interc_93_out ;
wire [0:0] direct_interc_94_out ;
wire [0:0] direct_interc_95_out ;
wire [0:0] direct_interc_96_out ;
wire [0:0] direct_interc_97_out ;
wire [0:0] direct_interc_98_out ;
wire [0:0] direct_interc_99_out ;
wire [0:0] direct_interc_9_out ;
wire [0:0] grid_clb_0_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_0_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_0_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_0_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_0_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_0_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_0_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_0_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_0_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_0_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_0_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_0_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_0_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_0_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_0_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_0_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_0_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_0_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_0_ccff_tail ;
wire [0:0] grid_clb_0_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_0_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_0_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_0_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_0_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_0_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_0_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_0_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_0_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_0_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_0_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_0_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_0_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_0_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_0_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_0_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_100_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_100_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_100_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_100_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_100_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_100_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_100_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_100_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_100_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_100_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_100_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_100_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_100_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_100_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_100_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_100_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_100_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_100_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_100_ccff_tail ;
wire [0:0] grid_clb_100_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_100_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_100_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_100_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_100_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_100_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_100_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_100_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_100_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_100_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_100_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_100_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_100_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_100_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_100_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_100_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_101_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_101_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_101_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_101_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_101_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_101_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_101_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_101_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_101_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_101_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_101_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_101_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_101_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_101_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_101_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_101_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_101_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_101_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_101_ccff_tail ;
wire [0:0] grid_clb_101_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_101_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_101_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_101_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_101_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_101_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_101_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_101_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_101_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_101_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_101_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_101_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_101_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_101_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_101_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_101_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_102_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_102_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_102_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_102_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_102_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_102_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_102_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_102_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_102_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_102_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_102_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_102_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_102_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_102_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_102_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_102_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_102_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_102_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_102_ccff_tail ;
wire [0:0] grid_clb_102_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_102_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_102_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_102_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_102_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_102_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_102_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_102_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_102_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_102_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_102_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_102_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_102_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_102_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_102_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_102_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_103_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_103_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_103_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_103_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_103_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_103_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_103_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_103_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_103_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_103_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_103_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_103_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_103_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_103_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_103_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_103_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_103_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_103_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_103_ccff_tail ;
wire [0:0] grid_clb_103_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_103_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_103_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_103_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_103_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_103_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_103_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_103_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_103_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_103_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_103_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_103_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_103_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_103_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_103_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_103_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_104_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_104_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_104_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_104_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_104_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_104_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_104_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_104_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_104_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_104_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_104_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_104_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_104_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_104_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_104_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_104_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_104_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_104_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_104_ccff_tail ;
wire [0:0] grid_clb_104_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_104_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_104_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_104_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_104_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_104_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_104_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_104_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_104_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_104_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_104_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_104_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_104_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_104_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_104_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_104_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_105_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_105_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_105_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_105_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_105_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_105_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_105_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_105_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_105_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_105_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_105_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_105_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_105_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_105_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_105_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_105_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_105_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_105_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_105_ccff_tail ;
wire [0:0] grid_clb_105_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_105_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_105_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_105_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_105_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_105_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_105_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_105_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_105_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_105_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_105_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_105_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_105_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_105_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_105_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_105_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_106_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_106_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_106_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_106_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_106_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_106_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_106_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_106_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_106_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_106_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_106_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_106_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_106_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_106_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_106_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_106_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_106_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_106_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_106_ccff_tail ;
wire [0:0] grid_clb_106_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_106_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_106_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_106_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_106_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_106_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_106_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_106_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_106_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_106_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_106_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_106_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_106_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_106_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_106_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_106_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_107_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_107_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_107_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_107_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_107_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_107_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_107_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_107_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_107_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_107_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_107_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_107_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_107_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_107_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_107_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_107_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_107_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_107_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_107_ccff_tail ;
wire [0:0] grid_clb_107_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_107_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_107_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_107_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_107_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_107_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_107_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_107_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_107_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_107_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_107_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_107_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_107_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_107_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_107_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_107_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_108_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_108_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_108_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_108_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_108_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_108_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_108_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_108_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_108_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_108_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_108_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_108_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_108_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_108_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_108_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_108_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_108_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_108_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_108_ccff_tail ;
wire [0:0] grid_clb_108_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_108_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_108_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_108_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_108_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_108_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_108_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_108_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_108_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_108_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_108_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_108_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_108_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_108_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_108_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_108_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_109_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_109_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_109_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_109_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_109_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_109_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_109_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_109_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_109_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_109_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_109_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_109_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_109_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_109_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_109_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_109_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_109_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_109_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_109_ccff_tail ;
wire [0:0] grid_clb_109_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_109_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_109_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_109_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_109_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_109_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_109_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_109_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_109_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_109_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_109_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_109_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_109_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_109_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_109_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_109_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_10_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_10_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_10_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_10_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_10_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_10_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_10_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_10_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_10_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_10_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_10_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_10_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_10_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_10_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_10_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_10_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_10_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_10_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_10_ccff_tail ;
wire [0:0] grid_clb_10_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_10_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_10_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_10_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_10_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_10_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_10_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_10_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_10_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_10_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_10_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_10_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_10_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_10_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_10_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_10_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_110_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_110_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_110_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_110_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_110_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_110_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_110_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_110_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_110_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_110_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_110_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_110_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_110_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_110_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_110_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_110_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_110_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_110_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_110_ccff_tail ;
wire [0:0] grid_clb_110_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_110_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_110_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_110_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_110_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_110_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_110_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_110_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_110_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_110_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_110_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_110_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_110_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_110_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_110_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_110_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_111_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_111_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_111_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_111_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_111_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_111_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_111_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_111_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_111_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_111_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_111_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_111_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_111_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_111_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_111_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_111_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_111_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_111_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_111_ccff_tail ;
wire [0:0] grid_clb_111_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_111_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_111_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_111_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_111_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_111_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_111_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_111_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_111_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_111_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_111_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_111_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_111_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_111_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_111_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_111_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_112_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_112_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_112_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_112_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_112_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_112_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_112_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_112_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_112_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_112_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_112_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_112_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_112_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_112_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_112_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_112_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_112_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_112_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_112_ccff_tail ;
wire [0:0] grid_clb_112_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_112_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_112_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_112_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_112_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_112_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_112_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_112_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_112_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_112_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_112_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_112_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_112_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_112_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_112_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_112_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_113_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_113_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_113_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_113_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_113_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_113_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_113_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_113_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_113_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_113_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_113_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_113_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_113_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_113_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_113_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_113_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_113_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_113_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_113_ccff_tail ;
wire [0:0] grid_clb_113_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_113_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_113_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_113_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_113_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_113_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_113_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_113_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_113_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_113_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_113_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_113_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_113_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_113_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_113_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_113_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_114_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_114_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_114_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_114_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_114_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_114_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_114_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_114_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_114_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_114_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_114_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_114_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_114_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_114_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_114_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_114_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_114_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_114_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_114_ccff_tail ;
wire [0:0] grid_clb_114_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_114_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_114_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_114_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_114_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_114_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_114_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_114_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_114_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_114_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_114_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_114_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_114_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_114_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_114_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_114_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_115_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_115_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_115_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_115_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_115_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_115_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_115_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_115_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_115_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_115_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_115_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_115_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_115_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_115_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_115_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_115_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_115_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_115_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_115_ccff_tail ;
wire [0:0] grid_clb_115_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_115_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_115_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_115_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_115_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_115_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_115_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_115_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_115_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_115_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_115_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_115_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_115_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_115_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_115_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_115_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_116_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_116_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_116_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_116_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_116_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_116_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_116_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_116_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_116_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_116_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_116_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_116_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_116_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_116_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_116_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_116_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_116_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_116_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_116_ccff_tail ;
wire [0:0] grid_clb_116_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_116_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_116_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_116_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_116_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_116_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_116_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_116_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_116_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_116_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_116_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_116_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_116_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_116_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_116_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_116_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_117_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_117_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_117_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_117_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_117_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_117_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_117_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_117_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_117_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_117_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_117_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_117_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_117_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_117_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_117_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_117_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_117_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_117_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_117_ccff_tail ;
wire [0:0] grid_clb_117_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_117_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_117_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_117_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_117_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_117_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_117_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_117_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_117_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_117_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_117_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_117_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_117_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_117_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_117_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_117_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_118_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_118_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_118_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_118_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_118_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_118_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_118_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_118_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_118_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_118_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_118_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_118_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_118_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_118_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_118_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_118_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_118_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_118_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_118_ccff_tail ;
wire [0:0] grid_clb_118_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_118_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_118_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_118_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_118_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_118_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_118_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_118_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_118_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_118_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_118_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_118_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_118_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_118_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_118_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_118_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_119_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_119_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_119_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_119_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_119_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_119_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_119_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_119_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_119_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_119_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_119_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_119_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_119_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_119_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_119_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_119_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_119_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_119_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_119_ccff_tail ;
wire [0:0] grid_clb_119_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_119_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_119_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_119_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_119_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_119_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_119_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_119_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_119_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_119_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_119_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_119_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_119_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_119_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_119_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_119_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_11_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_11_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_11_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_11_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_11_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_11_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_11_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_11_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_11_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_11_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_11_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_11_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_11_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_11_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_11_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_11_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_11_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_11_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_11_ccff_tail ;
wire [0:0] grid_clb_11_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_11_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_11_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_11_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_11_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_11_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_11_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_11_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_11_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_11_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_11_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_11_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_11_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_11_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_11_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_11_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_120_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_120_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_120_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_120_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_120_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_120_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_120_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_120_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_120_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_120_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_120_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_120_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_120_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_120_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_120_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_120_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_120_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_120_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_120_ccff_tail ;
wire [0:0] grid_clb_120_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_120_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_120_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_120_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_120_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_120_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_120_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_120_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_120_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_120_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_120_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_120_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_120_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_120_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_120_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_120_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_121_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_121_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_121_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_121_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_121_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_121_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_121_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_121_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_121_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_121_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_121_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_121_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_121_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_121_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_121_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_121_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_121_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_121_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_121_ccff_tail ;
wire [0:0] grid_clb_121_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_121_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_121_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_121_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_121_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_121_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_121_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_121_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_121_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_121_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_121_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_121_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_121_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_121_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_121_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_121_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_122_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_122_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_122_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_122_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_122_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_122_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_122_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_122_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_122_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_122_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_122_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_122_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_122_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_122_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_122_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_122_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_122_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_122_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_122_ccff_tail ;
wire [0:0] grid_clb_122_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_122_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_122_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_122_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_122_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_122_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_122_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_122_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_122_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_122_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_122_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_122_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_122_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_122_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_122_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_122_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_123_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_123_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_123_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_123_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_123_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_123_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_123_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_123_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_123_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_123_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_123_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_123_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_123_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_123_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_123_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_123_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_123_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_123_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_123_ccff_tail ;
wire [0:0] grid_clb_123_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_123_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_123_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_123_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_123_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_123_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_123_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_123_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_123_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_123_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_123_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_123_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_123_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_123_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_123_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_123_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_124_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_124_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_124_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_124_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_124_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_124_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_124_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_124_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_124_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_124_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_124_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_124_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_124_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_124_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_124_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_124_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_124_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_124_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_124_ccff_tail ;
wire [0:0] grid_clb_124_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_124_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_124_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_124_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_124_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_124_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_124_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_124_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_124_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_124_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_124_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_124_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_124_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_124_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_124_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_124_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_125_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_125_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_125_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_125_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_125_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_125_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_125_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_125_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_125_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_125_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_125_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_125_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_125_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_125_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_125_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_125_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_125_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_125_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_125_ccff_tail ;
wire [0:0] grid_clb_125_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_125_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_125_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_125_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_125_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_125_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_125_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_125_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_125_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_125_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_125_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_125_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_125_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_125_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_125_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_125_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_126_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_126_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_126_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_126_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_126_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_126_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_126_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_126_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_126_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_126_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_126_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_126_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_126_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_126_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_126_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_126_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_126_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_126_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_126_ccff_tail ;
wire [0:0] grid_clb_126_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_126_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_126_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_126_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_126_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_126_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_126_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_126_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_126_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_126_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_126_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_126_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_126_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_126_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_126_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_126_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_127_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_127_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_127_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_127_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_127_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_127_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_127_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_127_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_127_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_127_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_127_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_127_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_127_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_127_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_127_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_127_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_127_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_127_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_127_ccff_tail ;
wire [0:0] grid_clb_127_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_127_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_127_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_127_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_127_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_127_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_127_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_127_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_127_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_127_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_127_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_127_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_127_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_127_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_127_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_127_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_128_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_128_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_128_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_128_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_128_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_128_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_128_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_128_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_128_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_128_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_128_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_128_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_128_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_128_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_128_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_128_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_128_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_128_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_128_ccff_tail ;
wire [0:0] grid_clb_128_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_128_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_128_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_128_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_128_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_128_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_128_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_128_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_128_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_128_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_128_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_128_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_128_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_128_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_128_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_128_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_129_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_129_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_129_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_129_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_129_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_129_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_129_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_129_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_129_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_129_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_129_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_129_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_129_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_129_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_129_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_129_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_129_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_129_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_129_ccff_tail ;
wire [0:0] grid_clb_129_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_129_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_129_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_129_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_129_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_129_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_129_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_129_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_129_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_129_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_129_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_129_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_129_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_129_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_129_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_129_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_12__1__undriven_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_12__1__undriven_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_12_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_12_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_12_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_12_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_12_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_12_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_12_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_12_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_12_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_12_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_12_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_12_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_12_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_12_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_12_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_12_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_12_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_12_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_12_ccff_tail ;
wire [0:0] grid_clb_12_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_12_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_12_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_12_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_12_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_12_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_12_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_12_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_12_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_12_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_12_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_12_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_12_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_12_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_12_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_12_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_130_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_130_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_130_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_130_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_130_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_130_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_130_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_130_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_130_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_130_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_130_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_130_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_130_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_130_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_130_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_130_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_130_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_130_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_130_ccff_tail ;
wire [0:0] grid_clb_130_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_130_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_130_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_130_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_130_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_130_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_130_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_130_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_130_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_130_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_130_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_130_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_130_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_130_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_130_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_130_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_131_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_131_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_131_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_131_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_131_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_131_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_131_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_131_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_131_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_131_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_131_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_131_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_131_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_131_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_131_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_131_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_131_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_131_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_131_ccff_tail ;
wire [0:0] grid_clb_131_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_131_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_131_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_131_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_131_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_131_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_131_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_131_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_131_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_131_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_131_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_131_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_131_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_131_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_131_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_131_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_132_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_132_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_132_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_132_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_132_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_132_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_132_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_132_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_132_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_132_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_132_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_132_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_132_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_132_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_132_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_132_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_132_ccff_tail ;
wire [0:0] grid_clb_132_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_132_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_132_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_132_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_132_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_132_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_132_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_132_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_132_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_132_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_132_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_132_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_132_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_132_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_132_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_132_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_133_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_133_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_133_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_133_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_133_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_133_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_133_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_133_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_133_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_133_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_133_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_133_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_133_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_133_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_133_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_133_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_133_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_133_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_133_ccff_tail ;
wire [0:0] grid_clb_133_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_133_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_133_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_133_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_133_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_133_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_133_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_133_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_133_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_133_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_133_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_133_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_133_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_133_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_133_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_133_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_134_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_134_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_134_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_134_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_134_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_134_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_134_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_134_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_134_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_134_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_134_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_134_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_134_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_134_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_134_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_134_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_134_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_134_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_134_ccff_tail ;
wire [0:0] grid_clb_134_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_134_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_134_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_134_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_134_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_134_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_134_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_134_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_134_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_134_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_134_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_134_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_134_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_134_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_134_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_134_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_135_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_135_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_135_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_135_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_135_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_135_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_135_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_135_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_135_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_135_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_135_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_135_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_135_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_135_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_135_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_135_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_135_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_135_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_135_ccff_tail ;
wire [0:0] grid_clb_135_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_135_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_135_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_135_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_135_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_135_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_135_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_135_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_135_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_135_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_135_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_135_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_135_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_135_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_135_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_135_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_136_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_136_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_136_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_136_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_136_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_136_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_136_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_136_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_136_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_136_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_136_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_136_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_136_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_136_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_136_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_136_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_136_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_136_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_136_ccff_tail ;
wire [0:0] grid_clb_136_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_136_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_136_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_136_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_136_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_136_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_136_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_136_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_136_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_136_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_136_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_136_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_136_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_136_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_136_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_136_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_137_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_137_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_137_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_137_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_137_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_137_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_137_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_137_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_137_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_137_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_137_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_137_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_137_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_137_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_137_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_137_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_137_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_137_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_137_ccff_tail ;
wire [0:0] grid_clb_137_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_137_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_137_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_137_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_137_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_137_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_137_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_137_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_137_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_137_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_137_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_137_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_137_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_137_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_137_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_137_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_138_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_138_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_138_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_138_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_138_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_138_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_138_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_138_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_138_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_138_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_138_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_138_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_138_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_138_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_138_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_138_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_138_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_138_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_138_ccff_tail ;
wire [0:0] grid_clb_138_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_138_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_138_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_138_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_138_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_138_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_138_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_138_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_138_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_138_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_138_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_138_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_138_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_138_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_138_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_138_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_139_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_139_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_139_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_139_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_139_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_139_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_139_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_139_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_139_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_139_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_139_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_139_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_139_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_139_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_139_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_139_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_139_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_139_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_139_ccff_tail ;
wire [0:0] grid_clb_139_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_139_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_139_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_139_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_139_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_139_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_139_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_139_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_139_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_139_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_139_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_139_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_139_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_139_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_139_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_139_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_13_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_13_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_13_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_13_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_13_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_13_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_13_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_13_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_13_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_13_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_13_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_13_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_13_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_13_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_13_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_13_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_13_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_13_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_13_ccff_tail ;
wire [0:0] grid_clb_13_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_13_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_13_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_13_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_13_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_13_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_13_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_13_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_13_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_13_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_13_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_13_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_13_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_13_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_13_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_13_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_140_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_140_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_140_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_140_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_140_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_140_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_140_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_140_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_140_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_140_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_140_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_140_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_140_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_140_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_140_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_140_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_140_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_140_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_140_ccff_tail ;
wire [0:0] grid_clb_140_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_140_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_140_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_140_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_140_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_140_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_140_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_140_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_140_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_140_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_140_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_140_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_140_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_140_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_140_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_140_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_141_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_141_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_141_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_141_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_141_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_141_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_141_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_141_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_141_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_141_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_141_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_141_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_141_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_141_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_141_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_141_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_141_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_141_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_141_ccff_tail ;
wire [0:0] grid_clb_141_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_141_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_141_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_141_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_141_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_141_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_141_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_141_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_141_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_141_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_141_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_141_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_141_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_141_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_141_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_141_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_142_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_142_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_142_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_142_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_142_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_142_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_142_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_142_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_142_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_142_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_142_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_142_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_142_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_142_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_142_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_142_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_142_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_142_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_142_ccff_tail ;
wire [0:0] grid_clb_142_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_142_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_142_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_142_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_142_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_142_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_142_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_142_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_142_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_142_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_142_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_142_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_142_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_142_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_142_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_142_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_143_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_143_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_143_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_143_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_143_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_143_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_143_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_143_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_143_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_143_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_143_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_143_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_143_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_143_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_143_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_143_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_143_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_143_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_143_ccff_tail ;
wire [0:0] grid_clb_143_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_143_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_143_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_143_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_143_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_143_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_143_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_143_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_143_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_143_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_143_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_143_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_143_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_143_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_143_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_143_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_14_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_14_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_14_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_14_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_14_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_14_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_14_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_14_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_14_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_14_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_14_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_14_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_14_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_14_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_14_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_14_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_14_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_14_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_14_ccff_tail ;
wire [0:0] grid_clb_14_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_14_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_14_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_14_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_14_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_14_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_14_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_14_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_14_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_14_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_14_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_14_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_14_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_14_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_14_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_14_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_15_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_15_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_15_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_15_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_15_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_15_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_15_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_15_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_15_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_15_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_15_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_15_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_15_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_15_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_15_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_15_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_15_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_15_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_15_ccff_tail ;
wire [0:0] grid_clb_15_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_15_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_15_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_15_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_15_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_15_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_15_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_15_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_15_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_15_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_15_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_15_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_15_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_15_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_15_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_15_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_16_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_16_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_16_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_16_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_16_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_16_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_16_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_16_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_16_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_16_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_16_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_16_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_16_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_16_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_16_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_16_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_16_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_16_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_16_ccff_tail ;
wire [0:0] grid_clb_16_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_16_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_16_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_16_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_16_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_16_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_16_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_16_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_16_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_16_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_16_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_16_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_16_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_16_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_16_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_16_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_17_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_17_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_17_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_17_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_17_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_17_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_17_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_17_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_17_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_17_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_17_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_17_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_17_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_17_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_17_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_17_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_17_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_17_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_17_ccff_tail ;
wire [0:0] grid_clb_17_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_17_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_17_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_17_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_17_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_17_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_17_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_17_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_17_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_17_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_17_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_17_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_17_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_17_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_17_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_17_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_18_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_18_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_18_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_18_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_18_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_18_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_18_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_18_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_18_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_18_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_18_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_18_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_18_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_18_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_18_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_18_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_18_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_18_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_18_ccff_tail ;
wire [0:0] grid_clb_18_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_18_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_18_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_18_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_18_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_18_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_18_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_18_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_18_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_18_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_18_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_18_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_18_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_18_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_18_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_18_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_19_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_19_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_19_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_19_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_19_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_19_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_19_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_19_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_19_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_19_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_19_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_19_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_19_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_19_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_19_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_19_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_19_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_19_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_19_ccff_tail ;
wire [0:0] grid_clb_19_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_19_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_19_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_19_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_19_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_19_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_19_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_19_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_19_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_19_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_19_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_19_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_19_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_19_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_19_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_19_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_1__12__undriven_top_width_0_height_0__pin_32_ ;
wire [0:0] grid_clb_1__12__undriven_top_width_0_height_0__pin_33_ ;
wire [0:0] grid_clb_1_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_1_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_1_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_1_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_1_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_1_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_1_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_1_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_1_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_1_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_1_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_1_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_1_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_1_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_1_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_1_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_1_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_1_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_1_ccff_tail ;
wire [0:0] grid_clb_1_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_1_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_1_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_1_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_1_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_1_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_1_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_1_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_1_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_1_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_1_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_1_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_1_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_1_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_1_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_1_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_20_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_20_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_20_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_20_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_20_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_20_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_20_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_20_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_20_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_20_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_20_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_20_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_20_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_20_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_20_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_20_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_20_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_20_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_20_ccff_tail ;
wire [0:0] grid_clb_20_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_20_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_20_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_20_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_20_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_20_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_20_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_20_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_20_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_20_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_20_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_20_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_20_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_20_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_20_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_20_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_21_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_21_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_21_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_21_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_21_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_21_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_21_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_21_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_21_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_21_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_21_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_21_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_21_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_21_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_21_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_21_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_21_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_21_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_21_ccff_tail ;
wire [0:0] grid_clb_21_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_21_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_21_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_21_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_21_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_21_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_21_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_21_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_21_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_21_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_21_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_21_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_21_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_21_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_21_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_21_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_22_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_22_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_22_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_22_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_22_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_22_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_22_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_22_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_22_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_22_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_22_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_22_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_22_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_22_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_22_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_22_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_22_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_22_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_22_ccff_tail ;
wire [0:0] grid_clb_22_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_22_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_22_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_22_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_22_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_22_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_22_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_22_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_22_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_22_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_22_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_22_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_22_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_22_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_22_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_22_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_23_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_23_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_23_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_23_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_23_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_23_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_23_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_23_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_23_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_23_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_23_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_23_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_23_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_23_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_23_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_23_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_23_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_23_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_23_ccff_tail ;
wire [0:0] grid_clb_23_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_23_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_23_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_23_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_23_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_23_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_23_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_23_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_23_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_23_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_23_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_23_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_23_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_23_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_23_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_23_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_24_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_24_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_24_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_24_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_24_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_24_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_24_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_24_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_24_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_24_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_24_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_24_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_24_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_24_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_24_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_24_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_24_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_24_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_24_ccff_tail ;
wire [0:0] grid_clb_24_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_24_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_24_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_24_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_24_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_24_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_24_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_24_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_24_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_24_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_24_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_24_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_24_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_24_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_24_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_24_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_25_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_25_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_25_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_25_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_25_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_25_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_25_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_25_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_25_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_25_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_25_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_25_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_25_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_25_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_25_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_25_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_25_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_25_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_25_ccff_tail ;
wire [0:0] grid_clb_25_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_25_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_25_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_25_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_25_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_25_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_25_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_25_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_25_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_25_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_25_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_25_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_25_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_25_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_25_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_25_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_26_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_26_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_26_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_26_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_26_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_26_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_26_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_26_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_26_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_26_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_26_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_26_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_26_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_26_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_26_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_26_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_26_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_26_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_26_ccff_tail ;
wire [0:0] grid_clb_26_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_26_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_26_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_26_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_26_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_26_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_26_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_26_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_26_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_26_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_26_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_26_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_26_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_26_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_26_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_26_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_27_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_27_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_27_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_27_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_27_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_27_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_27_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_27_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_27_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_27_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_27_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_27_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_27_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_27_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_27_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_27_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_27_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_27_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_27_ccff_tail ;
wire [0:0] grid_clb_27_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_27_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_27_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_27_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_27_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_27_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_27_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_27_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_27_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_27_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_27_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_27_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_27_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_27_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_27_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_27_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_28_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_28_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_28_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_28_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_28_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_28_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_28_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_28_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_28_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_28_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_28_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_28_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_28_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_28_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_28_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_28_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_28_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_28_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_28_ccff_tail ;
wire [0:0] grid_clb_28_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_28_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_28_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_28_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_28_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_28_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_28_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_28_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_28_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_28_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_28_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_28_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_28_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_28_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_28_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_28_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_29_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_29_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_29_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_29_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_29_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_29_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_29_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_29_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_29_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_29_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_29_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_29_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_29_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_29_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_29_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_29_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_29_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_29_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_29_ccff_tail ;
wire [0:0] grid_clb_29_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_29_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_29_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_29_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_29_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_29_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_29_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_29_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_29_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_29_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_29_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_29_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_29_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_29_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_29_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_29_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_2_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_2_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_2_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_2_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_2_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_2_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_2_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_2_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_2_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_2_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_2_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_2_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_2_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_2_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_2_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_2_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_2_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_2_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_2_ccff_tail ;
wire [0:0] grid_clb_2_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_2_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_2_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_2_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_2_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_2_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_2_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_2_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_2_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_2_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_2_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_2_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_2_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_2_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_2_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_2_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_30_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_30_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_30_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_30_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_30_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_30_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_30_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_30_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_30_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_30_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_30_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_30_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_30_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_30_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_30_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_30_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_30_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_30_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_30_ccff_tail ;
wire [0:0] grid_clb_30_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_30_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_30_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_30_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_30_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_30_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_30_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_30_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_30_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_30_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_30_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_30_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_30_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_30_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_30_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_30_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_31_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_31_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_31_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_31_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_31_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_31_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_31_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_31_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_31_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_31_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_31_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_31_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_31_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_31_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_31_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_31_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_31_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_31_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_31_ccff_tail ;
wire [0:0] grid_clb_31_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_31_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_31_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_31_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_31_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_31_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_31_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_31_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_31_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_31_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_31_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_31_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_31_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_31_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_31_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_31_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_32_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_32_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_32_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_32_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_32_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_32_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_32_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_32_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_32_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_32_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_32_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_32_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_32_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_32_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_32_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_32_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_32_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_32_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_32_ccff_tail ;
wire [0:0] grid_clb_32_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_32_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_32_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_32_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_32_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_32_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_32_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_32_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_32_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_32_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_32_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_32_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_32_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_32_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_32_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_32_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_33_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_33_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_33_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_33_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_33_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_33_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_33_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_33_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_33_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_33_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_33_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_33_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_33_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_33_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_33_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_33_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_33_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_33_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_33_ccff_tail ;
wire [0:0] grid_clb_33_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_33_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_33_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_33_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_33_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_33_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_33_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_33_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_33_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_33_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_33_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_33_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_33_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_33_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_33_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_33_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_34_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_34_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_34_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_34_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_34_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_34_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_34_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_34_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_34_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_34_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_34_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_34_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_34_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_34_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_34_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_34_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_34_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_34_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_34_ccff_tail ;
wire [0:0] grid_clb_34_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_34_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_34_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_34_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_34_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_34_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_34_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_34_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_34_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_34_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_34_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_34_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_34_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_34_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_34_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_34_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_35_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_35_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_35_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_35_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_35_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_35_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_35_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_35_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_35_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_35_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_35_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_35_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_35_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_35_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_35_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_35_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_35_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_35_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_35_ccff_tail ;
wire [0:0] grid_clb_35_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_35_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_35_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_35_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_35_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_35_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_35_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_35_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_35_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_35_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_35_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_35_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_35_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_35_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_35_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_35_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_36_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_36_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_36_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_36_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_36_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_36_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_36_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_36_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_36_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_36_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_36_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_36_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_36_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_36_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_36_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_36_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_36_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_36_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_36_ccff_tail ;
wire [0:0] grid_clb_36_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_36_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_36_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_36_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_36_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_36_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_36_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_36_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_36_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_36_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_36_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_36_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_36_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_36_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_36_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_36_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_37_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_37_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_37_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_37_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_37_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_37_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_37_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_37_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_37_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_37_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_37_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_37_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_37_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_37_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_37_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_37_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_37_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_37_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_37_ccff_tail ;
wire [0:0] grid_clb_37_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_37_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_37_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_37_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_37_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_37_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_37_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_37_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_37_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_37_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_37_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_37_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_37_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_37_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_37_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_37_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_38_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_38_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_38_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_38_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_38_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_38_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_38_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_38_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_38_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_38_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_38_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_38_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_38_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_38_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_38_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_38_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_38_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_38_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_38_ccff_tail ;
wire [0:0] grid_clb_38_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_38_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_38_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_38_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_38_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_38_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_38_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_38_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_38_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_38_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_38_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_38_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_38_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_38_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_38_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_38_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_39_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_39_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_39_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_39_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_39_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_39_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_39_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_39_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_39_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_39_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_39_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_39_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_39_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_39_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_39_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_39_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_39_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_39_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_39_ccff_tail ;
wire [0:0] grid_clb_39_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_39_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_39_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_39_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_39_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_39_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_39_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_39_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_39_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_39_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_39_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_39_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_39_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_39_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_39_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_39_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_3_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_3_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_3_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_3_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_3_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_3_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_3_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_3_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_3_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_3_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_3_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_3_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_3_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_3_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_3_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_3_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_3_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_3_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_3_ccff_tail ;
wire [0:0] grid_clb_3_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_3_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_3_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_3_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_3_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_3_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_3_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_3_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_3_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_3_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_3_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_3_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_3_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_3_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_3_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_3_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_40_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_40_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_40_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_40_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_40_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_40_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_40_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_40_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_40_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_40_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_40_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_40_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_40_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_40_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_40_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_40_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_40_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_40_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_40_ccff_tail ;
wire [0:0] grid_clb_40_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_40_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_40_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_40_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_40_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_40_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_40_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_40_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_40_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_40_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_40_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_40_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_40_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_40_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_40_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_40_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_41_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_41_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_41_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_41_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_41_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_41_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_41_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_41_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_41_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_41_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_41_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_41_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_41_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_41_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_41_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_41_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_41_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_41_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_41_ccff_tail ;
wire [0:0] grid_clb_41_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_41_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_41_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_41_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_41_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_41_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_41_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_41_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_41_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_41_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_41_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_41_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_41_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_41_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_41_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_41_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_42_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_42_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_42_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_42_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_42_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_42_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_42_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_42_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_42_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_42_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_42_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_42_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_42_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_42_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_42_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_42_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_42_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_42_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_42_ccff_tail ;
wire [0:0] grid_clb_42_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_42_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_42_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_42_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_42_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_42_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_42_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_42_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_42_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_42_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_42_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_42_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_42_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_42_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_42_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_42_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_43_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_43_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_43_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_43_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_43_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_43_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_43_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_43_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_43_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_43_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_43_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_43_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_43_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_43_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_43_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_43_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_43_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_43_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_43_ccff_tail ;
wire [0:0] grid_clb_43_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_43_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_43_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_43_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_43_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_43_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_43_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_43_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_43_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_43_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_43_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_43_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_43_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_43_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_43_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_43_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_44_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_44_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_44_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_44_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_44_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_44_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_44_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_44_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_44_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_44_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_44_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_44_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_44_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_44_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_44_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_44_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_44_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_44_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_44_ccff_tail ;
wire [0:0] grid_clb_44_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_44_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_44_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_44_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_44_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_44_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_44_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_44_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_44_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_44_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_44_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_44_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_44_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_44_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_44_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_44_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_45_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_45_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_45_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_45_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_45_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_45_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_45_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_45_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_45_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_45_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_45_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_45_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_45_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_45_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_45_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_45_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_45_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_45_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_45_ccff_tail ;
wire [0:0] grid_clb_45_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_45_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_45_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_45_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_45_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_45_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_45_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_45_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_45_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_45_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_45_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_45_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_45_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_45_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_45_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_45_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_46_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_46_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_46_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_46_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_46_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_46_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_46_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_46_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_46_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_46_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_46_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_46_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_46_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_46_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_46_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_46_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_46_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_46_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_46_ccff_tail ;
wire [0:0] grid_clb_46_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_46_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_46_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_46_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_46_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_46_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_46_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_46_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_46_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_46_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_46_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_46_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_46_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_46_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_46_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_46_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_47_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_47_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_47_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_47_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_47_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_47_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_47_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_47_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_47_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_47_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_47_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_47_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_47_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_47_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_47_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_47_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_47_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_47_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_47_ccff_tail ;
wire [0:0] grid_clb_47_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_47_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_47_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_47_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_47_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_47_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_47_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_47_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_47_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_47_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_47_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_47_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_47_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_47_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_47_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_47_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_48_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_48_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_48_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_48_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_48_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_48_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_48_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_48_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_48_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_48_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_48_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_48_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_48_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_48_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_48_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_48_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_48_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_48_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_48_ccff_tail ;
wire [0:0] grid_clb_48_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_48_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_48_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_48_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_48_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_48_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_48_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_48_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_48_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_48_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_48_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_48_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_48_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_48_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_48_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_48_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_49_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_49_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_49_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_49_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_49_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_49_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_49_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_49_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_49_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_49_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_49_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_49_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_49_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_49_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_49_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_49_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_49_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_49_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_49_ccff_tail ;
wire [0:0] grid_clb_49_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_49_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_49_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_49_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_49_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_49_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_49_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_49_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_49_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_49_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_49_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_49_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_49_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_49_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_49_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_49_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_4_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_4_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_4_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_4_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_4_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_4_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_4_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_4_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_4_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_4_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_4_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_4_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_4_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_4_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_4_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_4_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_4_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_4_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_4_ccff_tail ;
wire [0:0] grid_clb_4_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_4_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_4_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_4_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_4_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_4_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_4_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_4_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_4_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_4_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_4_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_4_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_4_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_4_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_4_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_4_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_50_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_50_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_50_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_50_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_50_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_50_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_50_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_50_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_50_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_50_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_50_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_50_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_50_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_50_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_50_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_50_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_50_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_50_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_50_ccff_tail ;
wire [0:0] grid_clb_50_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_50_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_50_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_50_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_50_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_50_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_50_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_50_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_50_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_50_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_50_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_50_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_50_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_50_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_50_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_50_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_51_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_51_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_51_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_51_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_51_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_51_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_51_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_51_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_51_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_51_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_51_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_51_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_51_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_51_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_51_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_51_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_51_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_51_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_51_ccff_tail ;
wire [0:0] grid_clb_51_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_51_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_51_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_51_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_51_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_51_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_51_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_51_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_51_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_51_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_51_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_51_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_51_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_51_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_51_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_51_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_52_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_52_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_52_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_52_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_52_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_52_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_52_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_52_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_52_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_52_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_52_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_52_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_52_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_52_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_52_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_52_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_52_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_52_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_52_ccff_tail ;
wire [0:0] grid_clb_52_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_52_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_52_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_52_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_52_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_52_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_52_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_52_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_52_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_52_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_52_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_52_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_52_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_52_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_52_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_52_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_53_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_53_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_53_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_53_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_53_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_53_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_53_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_53_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_53_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_53_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_53_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_53_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_53_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_53_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_53_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_53_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_53_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_53_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_53_ccff_tail ;
wire [0:0] grid_clb_53_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_53_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_53_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_53_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_53_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_53_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_53_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_53_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_53_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_53_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_53_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_53_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_53_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_53_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_53_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_53_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_54_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_54_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_54_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_54_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_54_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_54_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_54_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_54_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_54_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_54_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_54_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_54_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_54_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_54_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_54_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_54_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_54_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_54_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_54_ccff_tail ;
wire [0:0] grid_clb_54_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_54_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_54_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_54_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_54_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_54_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_54_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_54_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_54_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_54_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_54_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_54_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_54_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_54_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_54_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_54_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_55_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_55_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_55_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_55_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_55_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_55_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_55_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_55_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_55_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_55_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_55_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_55_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_55_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_55_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_55_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_55_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_55_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_55_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_55_ccff_tail ;
wire [0:0] grid_clb_55_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_55_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_55_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_55_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_55_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_55_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_55_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_55_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_55_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_55_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_55_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_55_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_55_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_55_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_55_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_55_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_56_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_56_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_56_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_56_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_56_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_56_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_56_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_56_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_56_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_56_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_56_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_56_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_56_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_56_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_56_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_56_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_56_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_56_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_56_ccff_tail ;
wire [0:0] grid_clb_56_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_56_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_56_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_56_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_56_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_56_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_56_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_56_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_56_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_56_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_56_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_56_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_56_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_56_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_56_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_56_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_57_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_57_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_57_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_57_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_57_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_57_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_57_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_57_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_57_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_57_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_57_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_57_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_57_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_57_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_57_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_57_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_57_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_57_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_57_ccff_tail ;
wire [0:0] grid_clb_57_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_57_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_57_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_57_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_57_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_57_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_57_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_57_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_57_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_57_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_57_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_57_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_57_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_57_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_57_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_57_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_58_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_58_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_58_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_58_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_58_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_58_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_58_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_58_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_58_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_58_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_58_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_58_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_58_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_58_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_58_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_58_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_58_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_58_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_58_ccff_tail ;
wire [0:0] grid_clb_58_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_58_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_58_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_58_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_58_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_58_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_58_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_58_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_58_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_58_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_58_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_58_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_58_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_58_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_58_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_58_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_59_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_59_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_59_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_59_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_59_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_59_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_59_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_59_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_59_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_59_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_59_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_59_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_59_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_59_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_59_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_59_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_59_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_59_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_59_ccff_tail ;
wire [0:0] grid_clb_59_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_59_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_59_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_59_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_59_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_59_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_59_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_59_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_59_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_59_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_59_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_59_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_59_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_59_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_59_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_59_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_5_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_5_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_5_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_5_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_5_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_5_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_5_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_5_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_5_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_5_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_5_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_5_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_5_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_5_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_5_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_5_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_5_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_5_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_5_ccff_tail ;
wire [0:0] grid_clb_5_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_5_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_5_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_5_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_5_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_5_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_5_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_5_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_5_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_5_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_5_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_5_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_5_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_5_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_5_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_5_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_60_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_60_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_60_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_60_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_60_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_60_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_60_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_60_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_60_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_60_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_60_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_60_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_60_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_60_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_60_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_60_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_60_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_60_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_60_ccff_tail ;
wire [0:0] grid_clb_60_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_60_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_60_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_60_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_60_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_60_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_60_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_60_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_60_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_60_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_60_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_60_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_60_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_60_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_60_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_60_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_61_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_61_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_61_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_61_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_61_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_61_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_61_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_61_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_61_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_61_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_61_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_61_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_61_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_61_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_61_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_61_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_61_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_61_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_61_ccff_tail ;
wire [0:0] grid_clb_61_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_61_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_61_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_61_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_61_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_61_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_61_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_61_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_61_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_61_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_61_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_61_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_61_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_61_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_61_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_61_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_62_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_62_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_62_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_62_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_62_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_62_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_62_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_62_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_62_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_62_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_62_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_62_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_62_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_62_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_62_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_62_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_62_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_62_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_62_ccff_tail ;
wire [0:0] grid_clb_62_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_62_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_62_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_62_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_62_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_62_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_62_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_62_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_62_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_62_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_62_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_62_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_62_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_62_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_62_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_62_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_63_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_63_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_63_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_63_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_63_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_63_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_63_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_63_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_63_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_63_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_63_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_63_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_63_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_63_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_63_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_63_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_63_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_63_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_63_ccff_tail ;
wire [0:0] grid_clb_63_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_63_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_63_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_63_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_63_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_63_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_63_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_63_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_63_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_63_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_63_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_63_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_63_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_63_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_63_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_63_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_64_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_64_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_64_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_64_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_64_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_64_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_64_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_64_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_64_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_64_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_64_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_64_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_64_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_64_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_64_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_64_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_64_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_64_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_64_ccff_tail ;
wire [0:0] grid_clb_64_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_64_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_64_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_64_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_64_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_64_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_64_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_64_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_64_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_64_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_64_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_64_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_64_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_64_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_64_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_64_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_65_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_65_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_65_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_65_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_65_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_65_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_65_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_65_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_65_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_65_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_65_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_65_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_65_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_65_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_65_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_65_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_65_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_65_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_65_ccff_tail ;
wire [0:0] grid_clb_65_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_65_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_65_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_65_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_65_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_65_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_65_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_65_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_65_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_65_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_65_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_65_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_65_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_65_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_65_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_65_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_66_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_66_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_66_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_66_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_66_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_66_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_66_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_66_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_66_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_66_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_66_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_66_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_66_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_66_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_66_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_66_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_66_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_66_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_66_ccff_tail ;
wire [0:0] grid_clb_66_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_66_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_66_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_66_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_66_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_66_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_66_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_66_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_66_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_66_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_66_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_66_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_66_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_66_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_66_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_66_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_67_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_67_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_67_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_67_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_67_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_67_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_67_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_67_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_67_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_67_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_67_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_67_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_67_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_67_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_67_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_67_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_67_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_67_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_67_ccff_tail ;
wire [0:0] grid_clb_67_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_67_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_67_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_67_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_67_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_67_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_67_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_67_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_67_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_67_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_67_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_67_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_67_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_67_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_67_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_67_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_68_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_68_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_68_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_68_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_68_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_68_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_68_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_68_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_68_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_68_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_68_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_68_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_68_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_68_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_68_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_68_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_68_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_68_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_68_ccff_tail ;
wire [0:0] grid_clb_68_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_68_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_68_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_68_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_68_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_68_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_68_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_68_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_68_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_68_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_68_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_68_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_68_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_68_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_68_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_68_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_69_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_69_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_69_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_69_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_69_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_69_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_69_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_69_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_69_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_69_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_69_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_69_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_69_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_69_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_69_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_69_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_69_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_69_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_69_ccff_tail ;
wire [0:0] grid_clb_69_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_69_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_69_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_69_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_69_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_69_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_69_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_69_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_69_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_69_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_69_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_69_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_69_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_69_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_69_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_69_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_6_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_6_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_6_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_6_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_6_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_6_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_6_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_6_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_6_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_6_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_6_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_6_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_6_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_6_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_6_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_6_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_6_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_6_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_6_ccff_tail ;
wire [0:0] grid_clb_6_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_6_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_6_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_6_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_6_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_6_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_6_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_6_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_6_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_6_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_6_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_6_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_6_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_6_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_6_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_6_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_70_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_70_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_70_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_70_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_70_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_70_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_70_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_70_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_70_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_70_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_70_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_70_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_70_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_70_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_70_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_70_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_70_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_70_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_70_ccff_tail ;
wire [0:0] grid_clb_70_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_70_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_70_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_70_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_70_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_70_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_70_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_70_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_70_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_70_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_70_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_70_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_70_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_70_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_70_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_70_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_71_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_71_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_71_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_71_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_71_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_71_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_71_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_71_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_71_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_71_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_71_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_71_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_71_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_71_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_71_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_71_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_71_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_71_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_71_ccff_tail ;
wire [0:0] grid_clb_71_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_71_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_71_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_71_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_71_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_71_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_71_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_71_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_71_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_71_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_71_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_71_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_71_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_71_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_71_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_71_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_72_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_72_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_72_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_72_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_72_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_72_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_72_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_72_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_72_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_72_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_72_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_72_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_72_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_72_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_72_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_72_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_72_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_72_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_72_ccff_tail ;
wire [0:0] grid_clb_72_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_72_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_72_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_72_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_72_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_72_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_72_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_72_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_72_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_72_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_72_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_72_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_72_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_72_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_72_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_72_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_73_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_73_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_73_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_73_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_73_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_73_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_73_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_73_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_73_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_73_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_73_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_73_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_73_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_73_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_73_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_73_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_73_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_73_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_73_ccff_tail ;
wire [0:0] grid_clb_73_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_73_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_73_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_73_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_73_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_73_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_73_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_73_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_73_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_73_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_73_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_73_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_73_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_73_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_73_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_73_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_74_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_74_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_74_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_74_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_74_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_74_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_74_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_74_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_74_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_74_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_74_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_74_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_74_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_74_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_74_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_74_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_74_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_74_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_74_ccff_tail ;
wire [0:0] grid_clb_74_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_74_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_74_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_74_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_74_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_74_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_74_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_74_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_74_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_74_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_74_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_74_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_74_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_74_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_74_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_74_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_75_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_75_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_75_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_75_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_75_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_75_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_75_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_75_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_75_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_75_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_75_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_75_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_75_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_75_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_75_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_75_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_75_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_75_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_75_ccff_tail ;
wire [0:0] grid_clb_75_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_75_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_75_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_75_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_75_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_75_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_75_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_75_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_75_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_75_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_75_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_75_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_75_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_75_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_75_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_75_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_76_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_76_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_76_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_76_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_76_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_76_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_76_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_76_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_76_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_76_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_76_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_76_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_76_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_76_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_76_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_76_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_76_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_76_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_76_ccff_tail ;
wire [0:0] grid_clb_76_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_76_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_76_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_76_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_76_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_76_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_76_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_76_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_76_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_76_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_76_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_76_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_76_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_76_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_76_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_76_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_77_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_77_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_77_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_77_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_77_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_77_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_77_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_77_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_77_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_77_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_77_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_77_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_77_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_77_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_77_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_77_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_77_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_77_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_77_ccff_tail ;
wire [0:0] grid_clb_77_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_77_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_77_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_77_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_77_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_77_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_77_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_77_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_77_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_77_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_77_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_77_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_77_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_77_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_77_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_77_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_78_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_78_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_78_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_78_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_78_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_78_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_78_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_78_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_78_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_78_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_78_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_78_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_78_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_78_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_78_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_78_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_78_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_78_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_78_ccff_tail ;
wire [0:0] grid_clb_78_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_78_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_78_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_78_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_78_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_78_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_78_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_78_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_78_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_78_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_78_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_78_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_78_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_78_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_78_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_78_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_79_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_79_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_79_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_79_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_79_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_79_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_79_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_79_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_79_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_79_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_79_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_79_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_79_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_79_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_79_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_79_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_79_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_79_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_79_ccff_tail ;
wire [0:0] grid_clb_79_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_79_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_79_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_79_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_79_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_79_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_79_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_79_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_79_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_79_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_79_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_79_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_79_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_79_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_79_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_79_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_7_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_7_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_7_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_7_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_7_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_7_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_7_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_7_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_7_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_7_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_7_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_7_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_7_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_7_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_7_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_7_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_7_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_7_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_7_ccff_tail ;
wire [0:0] grid_clb_7_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_7_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_7_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_7_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_7_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_7_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_7_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_7_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_7_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_7_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_7_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_7_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_7_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_7_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_7_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_7_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_80_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_80_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_80_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_80_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_80_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_80_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_80_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_80_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_80_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_80_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_80_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_80_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_80_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_80_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_80_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_80_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_80_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_80_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_80_ccff_tail ;
wire [0:0] grid_clb_80_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_80_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_80_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_80_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_80_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_80_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_80_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_80_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_80_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_80_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_80_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_80_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_80_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_80_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_80_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_80_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_81_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_81_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_81_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_81_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_81_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_81_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_81_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_81_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_81_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_81_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_81_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_81_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_81_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_81_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_81_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_81_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_81_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_81_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_81_ccff_tail ;
wire [0:0] grid_clb_81_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_81_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_81_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_81_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_81_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_81_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_81_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_81_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_81_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_81_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_81_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_81_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_81_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_81_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_81_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_81_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_82_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_82_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_82_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_82_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_82_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_82_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_82_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_82_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_82_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_82_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_82_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_82_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_82_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_82_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_82_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_82_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_82_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_82_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_82_ccff_tail ;
wire [0:0] grid_clb_82_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_82_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_82_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_82_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_82_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_82_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_82_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_82_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_82_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_82_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_82_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_82_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_82_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_82_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_82_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_82_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_83_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_83_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_83_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_83_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_83_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_83_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_83_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_83_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_83_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_83_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_83_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_83_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_83_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_83_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_83_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_83_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_83_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_83_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_83_ccff_tail ;
wire [0:0] grid_clb_83_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_83_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_83_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_83_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_83_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_83_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_83_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_83_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_83_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_83_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_83_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_83_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_83_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_83_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_83_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_83_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_84_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_84_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_84_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_84_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_84_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_84_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_84_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_84_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_84_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_84_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_84_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_84_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_84_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_84_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_84_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_84_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_84_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_84_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_84_ccff_tail ;
wire [0:0] grid_clb_84_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_84_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_84_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_84_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_84_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_84_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_84_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_84_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_84_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_84_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_84_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_84_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_84_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_84_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_84_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_84_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_85_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_85_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_85_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_85_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_85_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_85_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_85_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_85_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_85_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_85_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_85_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_85_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_85_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_85_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_85_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_85_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_85_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_85_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_85_ccff_tail ;
wire [0:0] grid_clb_85_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_85_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_85_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_85_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_85_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_85_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_85_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_85_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_85_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_85_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_85_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_85_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_85_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_85_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_85_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_85_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_86_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_86_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_86_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_86_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_86_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_86_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_86_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_86_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_86_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_86_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_86_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_86_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_86_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_86_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_86_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_86_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_86_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_86_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_86_ccff_tail ;
wire [0:0] grid_clb_86_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_86_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_86_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_86_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_86_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_86_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_86_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_86_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_86_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_86_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_86_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_86_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_86_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_86_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_86_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_86_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_87_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_87_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_87_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_87_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_87_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_87_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_87_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_87_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_87_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_87_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_87_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_87_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_87_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_87_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_87_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_87_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_87_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_87_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_87_ccff_tail ;
wire [0:0] grid_clb_87_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_87_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_87_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_87_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_87_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_87_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_87_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_87_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_87_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_87_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_87_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_87_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_87_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_87_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_87_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_87_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_88_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_88_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_88_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_88_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_88_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_88_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_88_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_88_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_88_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_88_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_88_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_88_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_88_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_88_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_88_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_88_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_88_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_88_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_88_ccff_tail ;
wire [0:0] grid_clb_88_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_88_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_88_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_88_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_88_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_88_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_88_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_88_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_88_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_88_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_88_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_88_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_88_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_88_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_88_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_88_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_89_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_89_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_89_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_89_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_89_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_89_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_89_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_89_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_89_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_89_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_89_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_89_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_89_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_89_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_89_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_89_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_89_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_89_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_89_ccff_tail ;
wire [0:0] grid_clb_89_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_89_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_89_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_89_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_89_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_89_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_89_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_89_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_89_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_89_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_89_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_89_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_89_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_89_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_89_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_89_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_8_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_8_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_8_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_8_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_8_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_8_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_8_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_8_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_8_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_8_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_8_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_8_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_8_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_8_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_8_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_8_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_8_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_8_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_8_ccff_tail ;
wire [0:0] grid_clb_8_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_8_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_8_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_8_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_8_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_8_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_8_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_8_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_8_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_8_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_8_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_8_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_8_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_8_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_8_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_8_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_90_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_90_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_90_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_90_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_90_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_90_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_90_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_90_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_90_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_90_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_90_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_90_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_90_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_90_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_90_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_90_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_90_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_90_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_90_ccff_tail ;
wire [0:0] grid_clb_90_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_90_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_90_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_90_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_90_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_90_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_90_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_90_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_90_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_90_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_90_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_90_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_90_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_90_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_90_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_90_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_91_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_91_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_91_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_91_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_91_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_91_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_91_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_91_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_91_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_91_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_91_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_91_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_91_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_91_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_91_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_91_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_91_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_91_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_91_ccff_tail ;
wire [0:0] grid_clb_91_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_91_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_91_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_91_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_91_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_91_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_91_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_91_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_91_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_91_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_91_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_91_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_91_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_91_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_91_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_91_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_92_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_92_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_92_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_92_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_92_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_92_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_92_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_92_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_92_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_92_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_92_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_92_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_92_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_92_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_92_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_92_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_92_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_92_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_92_ccff_tail ;
wire [0:0] grid_clb_92_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_92_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_92_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_92_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_92_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_92_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_92_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_92_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_92_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_92_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_92_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_92_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_92_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_92_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_92_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_92_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_93_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_93_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_93_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_93_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_93_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_93_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_93_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_93_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_93_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_93_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_93_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_93_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_93_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_93_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_93_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_93_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_93_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_93_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_93_ccff_tail ;
wire [0:0] grid_clb_93_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_93_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_93_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_93_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_93_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_93_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_93_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_93_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_93_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_93_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_93_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_93_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_93_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_93_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_93_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_93_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_94_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_94_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_94_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_94_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_94_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_94_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_94_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_94_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_94_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_94_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_94_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_94_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_94_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_94_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_94_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_94_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_94_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_94_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_94_ccff_tail ;
wire [0:0] grid_clb_94_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_94_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_94_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_94_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_94_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_94_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_94_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_94_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_94_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_94_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_94_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_94_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_94_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_94_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_94_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_94_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_95_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_95_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_95_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_95_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_95_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_95_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_95_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_95_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_95_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_95_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_95_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_95_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_95_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_95_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_95_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_95_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_95_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_95_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_95_ccff_tail ;
wire [0:0] grid_clb_95_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_95_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_95_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_95_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_95_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_95_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_95_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_95_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_95_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_95_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_95_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_95_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_95_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_95_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_95_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_95_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_96_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_96_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_96_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_96_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_96_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_96_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_96_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_96_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_96_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_96_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_96_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_96_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_96_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_96_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_96_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_96_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_96_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_96_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_96_ccff_tail ;
wire [0:0] grid_clb_96_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_96_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_96_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_96_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_96_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_96_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_96_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_96_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_96_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_96_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_96_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_96_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_96_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_96_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_96_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_96_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_97_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_97_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_97_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_97_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_97_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_97_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_97_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_97_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_97_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_97_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_97_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_97_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_97_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_97_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_97_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_97_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_97_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_97_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_97_ccff_tail ;
wire [0:0] grid_clb_97_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_97_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_97_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_97_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_97_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_97_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_97_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_97_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_97_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_97_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_97_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_97_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_97_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_97_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_97_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_97_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_98_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_98_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_98_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_98_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_98_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_98_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_98_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_98_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_98_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_98_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_98_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_98_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_98_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_98_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_98_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_98_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_98_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_98_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_98_ccff_tail ;
wire [0:0] grid_clb_98_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_98_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_98_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_98_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_98_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_98_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_98_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_98_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_98_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_98_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_98_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_98_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_98_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_98_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_98_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_98_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_99_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_99_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_99_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_99_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_99_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_99_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_99_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_99_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_99_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_99_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_99_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_99_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_99_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_99_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_99_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_99_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_99_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_99_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_99_ccff_tail ;
wire [0:0] grid_clb_99_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_99_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_99_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_99_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_99_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_99_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_99_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_99_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_99_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_99_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_99_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_99_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_99_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_99_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_99_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_99_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_9_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_9_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_9_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_9_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_9_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_9_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_9_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_9_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_9_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_9_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_9_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_9_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_9_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_9_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_9_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_9_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_9_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_9_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_9_ccff_tail ;
wire [0:0] grid_clb_9_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_9_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_9_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_9_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_9_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_9_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_9_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_9_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_9_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_9_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_9_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_9_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_9_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_9_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_9_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_9_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_io_bottom_0_ccff_tail ;
wire [0:0] grid_io_bottom_0_top_width_0_height_0__pin_1_lower ;
wire [0:0] grid_io_bottom_0_top_width_0_height_0__pin_1_upper ;
wire [0:0] grid_io_bottom_10_ccff_tail ;
wire [0:0] grid_io_bottom_10_top_width_0_height_0__pin_1_lower ;
wire [0:0] grid_io_bottom_10_top_width_0_height_0__pin_1_upper ;
wire [0:0] grid_io_bottom_11_ccff_tail ;
wire [0:0] grid_io_bottom_11_top_width_0_height_0__pin_1_lower ;
wire [0:0] grid_io_bottom_11_top_width_0_height_0__pin_1_upper ;
wire [0:0] grid_io_bottom_1_ccff_tail ;
wire [0:0] grid_io_bottom_1_top_width_0_height_0__pin_1_lower ;
wire [0:0] grid_io_bottom_1_top_width_0_height_0__pin_1_upper ;
wire [0:0] grid_io_bottom_2_ccff_tail ;
wire [0:0] grid_io_bottom_2_top_width_0_height_0__pin_1_lower ;
wire [0:0] grid_io_bottom_2_top_width_0_height_0__pin_1_upper ;
wire [0:0] grid_io_bottom_3_ccff_tail ;
wire [0:0] grid_io_bottom_3_top_width_0_height_0__pin_1_lower ;
wire [0:0] grid_io_bottom_3_top_width_0_height_0__pin_1_upper ;
wire [0:0] grid_io_bottom_4_ccff_tail ;
wire [0:0] grid_io_bottom_4_top_width_0_height_0__pin_1_lower ;
wire [0:0] grid_io_bottom_4_top_width_0_height_0__pin_1_upper ;
wire [0:0] grid_io_bottom_5_ccff_tail ;
wire [0:0] grid_io_bottom_5_top_width_0_height_0__pin_1_lower ;
wire [0:0] grid_io_bottom_5_top_width_0_height_0__pin_1_upper ;
wire [0:0] grid_io_bottom_6_ccff_tail ;
wire [0:0] grid_io_bottom_6_top_width_0_height_0__pin_1_lower ;
wire [0:0] grid_io_bottom_6_top_width_0_height_0__pin_1_upper ;
wire [0:0] grid_io_bottom_7_ccff_tail ;
wire [0:0] grid_io_bottom_7_top_width_0_height_0__pin_1_lower ;
wire [0:0] grid_io_bottom_7_top_width_0_height_0__pin_1_upper ;
wire [0:0] grid_io_bottom_8_ccff_tail ;
wire [0:0] grid_io_bottom_8_top_width_0_height_0__pin_1_lower ;
wire [0:0] grid_io_bottom_8_top_width_0_height_0__pin_1_upper ;
wire [0:0] grid_io_bottom_9_ccff_tail ;
wire [0:0] grid_io_bottom_9_top_width_0_height_0__pin_1_lower ;
wire [0:0] grid_io_bottom_9_top_width_0_height_0__pin_1_upper ;
wire [0:0] grid_io_left_0_ccff_tail ;
wire [0:0] grid_io_left_0_right_width_0_height_0__pin_1_lower ;
wire [0:0] grid_io_left_0_right_width_0_height_0__pin_1_upper ;
wire [0:0] grid_io_left_10_ccff_tail ;
wire [0:0] grid_io_left_10_right_width_0_height_0__pin_1_lower ;
wire [0:0] grid_io_left_10_right_width_0_height_0__pin_1_upper ;
wire [0:0] grid_io_left_11_ccff_tail ;
wire [0:0] grid_io_left_11_right_width_0_height_0__pin_1_lower ;
wire [0:0] grid_io_left_11_right_width_0_height_0__pin_1_upper ;
wire [0:0] grid_io_left_1_ccff_tail ;
wire [0:0] grid_io_left_1_right_width_0_height_0__pin_1_lower ;
wire [0:0] grid_io_left_1_right_width_0_height_0__pin_1_upper ;
wire [0:0] grid_io_left_2_ccff_tail ;
wire [0:0] grid_io_left_2_right_width_0_height_0__pin_1_lower ;
wire [0:0] grid_io_left_2_right_width_0_height_0__pin_1_upper ;
wire [0:0] grid_io_left_3_ccff_tail ;
wire [0:0] grid_io_left_3_right_width_0_height_0__pin_1_lower ;
wire [0:0] grid_io_left_3_right_width_0_height_0__pin_1_upper ;
wire [0:0] grid_io_left_4_ccff_tail ;
wire [0:0] grid_io_left_4_right_width_0_height_0__pin_1_lower ;
wire [0:0] grid_io_left_4_right_width_0_height_0__pin_1_upper ;
wire [0:0] grid_io_left_5_ccff_tail ;
wire [0:0] grid_io_left_5_right_width_0_height_0__pin_1_lower ;
wire [0:0] grid_io_left_5_right_width_0_height_0__pin_1_upper ;
wire [0:0] grid_io_left_6_ccff_tail ;
wire [0:0] grid_io_left_6_right_width_0_height_0__pin_1_lower ;
wire [0:0] grid_io_left_6_right_width_0_height_0__pin_1_upper ;
wire [0:0] grid_io_left_7_ccff_tail ;
wire [0:0] grid_io_left_7_right_width_0_height_0__pin_1_lower ;
wire [0:0] grid_io_left_7_right_width_0_height_0__pin_1_upper ;
wire [0:0] grid_io_left_8_ccff_tail ;
wire [0:0] grid_io_left_8_right_width_0_height_0__pin_1_lower ;
wire [0:0] grid_io_left_8_right_width_0_height_0__pin_1_upper ;
wire [0:0] grid_io_left_9_ccff_tail ;
wire [0:0] grid_io_left_9_right_width_0_height_0__pin_1_lower ;
wire [0:0] grid_io_left_9_right_width_0_height_0__pin_1_upper ;
wire [0:0] grid_io_right_0_ccff_tail ;
wire [0:0] grid_io_right_0_left_width_0_height_0__pin_1_lower ;
wire [0:0] grid_io_right_0_left_width_0_height_0__pin_1_upper ;
wire [0:0] grid_io_right_10_ccff_tail ;
wire [0:0] grid_io_right_10_left_width_0_height_0__pin_1_lower ;
wire [0:0] grid_io_right_10_left_width_0_height_0__pin_1_upper ;
wire [0:0] grid_io_right_11_ccff_tail ;
wire [0:0] grid_io_right_11_left_width_0_height_0__pin_1_lower ;
wire [0:0] grid_io_right_11_left_width_0_height_0__pin_1_upper ;
wire [0:0] grid_io_right_1_ccff_tail ;
wire [0:0] grid_io_right_1_left_width_0_height_0__pin_1_lower ;
wire [0:0] grid_io_right_1_left_width_0_height_0__pin_1_upper ;
wire [0:0] grid_io_right_2_ccff_tail ;
wire [0:0] grid_io_right_2_left_width_0_height_0__pin_1_lower ;
wire [0:0] grid_io_right_2_left_width_0_height_0__pin_1_upper ;
wire [0:0] grid_io_right_3_ccff_tail ;
wire [0:0] grid_io_right_3_left_width_0_height_0__pin_1_lower ;
wire [0:0] grid_io_right_3_left_width_0_height_0__pin_1_upper ;
wire [0:0] grid_io_right_4_ccff_tail ;
wire [0:0] grid_io_right_4_left_width_0_height_0__pin_1_lower ;
wire [0:0] grid_io_right_4_left_width_0_height_0__pin_1_upper ;
wire [0:0] grid_io_right_5_ccff_tail ;
wire [0:0] grid_io_right_5_left_width_0_height_0__pin_1_lower ;
wire [0:0] grid_io_right_5_left_width_0_height_0__pin_1_upper ;
wire [0:0] grid_io_right_6_ccff_tail ;
wire [0:0] grid_io_right_6_left_width_0_height_0__pin_1_lower ;
wire [0:0] grid_io_right_6_left_width_0_height_0__pin_1_upper ;
wire [0:0] grid_io_right_7_ccff_tail ;
wire [0:0] grid_io_right_7_left_width_0_height_0__pin_1_lower ;
wire [0:0] grid_io_right_7_left_width_0_height_0__pin_1_upper ;
wire [0:0] grid_io_right_8_ccff_tail ;
wire [0:0] grid_io_right_8_left_width_0_height_0__pin_1_lower ;
wire [0:0] grid_io_right_8_left_width_0_height_0__pin_1_upper ;
wire [0:0] grid_io_right_9_ccff_tail ;
wire [0:0] grid_io_right_9_left_width_0_height_0__pin_1_lower ;
wire [0:0] grid_io_right_9_left_width_0_height_0__pin_1_upper ;
wire [0:0] grid_io_top_0_bottom_width_0_height_0__pin_1_lower ;
wire [0:0] grid_io_top_0_bottom_width_0_height_0__pin_1_upper ;
wire [0:0] grid_io_top_0_ccff_tail ;
wire [0:0] grid_io_top_10_bottom_width_0_height_0__pin_1_lower ;
wire [0:0] grid_io_top_10_bottom_width_0_height_0__pin_1_upper ;
wire [0:0] grid_io_top_10_ccff_tail ;
wire [0:0] grid_io_top_11_bottom_width_0_height_0__pin_1_lower ;
wire [0:0] grid_io_top_11_bottom_width_0_height_0__pin_1_upper ;
wire [0:0] grid_io_top_11_ccff_tail ;
wire [0:0] grid_io_top_1_bottom_width_0_height_0__pin_1_lower ;
wire [0:0] grid_io_top_1_bottom_width_0_height_0__pin_1_upper ;
wire [0:0] grid_io_top_1_ccff_tail ;
wire [0:0] grid_io_top_2_bottom_width_0_height_0__pin_1_lower ;
wire [0:0] grid_io_top_2_bottom_width_0_height_0__pin_1_upper ;
wire [0:0] grid_io_top_2_ccff_tail ;
wire [0:0] grid_io_top_3_bottom_width_0_height_0__pin_1_lower ;
wire [0:0] grid_io_top_3_bottom_width_0_height_0__pin_1_upper ;
wire [0:0] grid_io_top_3_ccff_tail ;
wire [0:0] grid_io_top_4_bottom_width_0_height_0__pin_1_lower ;
wire [0:0] grid_io_top_4_bottom_width_0_height_0__pin_1_upper ;
wire [0:0] grid_io_top_4_ccff_tail ;
wire [0:0] grid_io_top_5_bottom_width_0_height_0__pin_1_lower ;
wire [0:0] grid_io_top_5_bottom_width_0_height_0__pin_1_upper ;
wire [0:0] grid_io_top_5_ccff_tail ;
wire [0:0] grid_io_top_6_bottom_width_0_height_0__pin_1_lower ;
wire [0:0] grid_io_top_6_bottom_width_0_height_0__pin_1_upper ;
wire [0:0] grid_io_top_6_ccff_tail ;
wire [0:0] grid_io_top_7_bottom_width_0_height_0__pin_1_lower ;
wire [0:0] grid_io_top_7_bottom_width_0_height_0__pin_1_upper ;
wire [0:0] grid_io_top_7_ccff_tail ;
wire [0:0] grid_io_top_8_bottom_width_0_height_0__pin_1_lower ;
wire [0:0] grid_io_top_8_bottom_width_0_height_0__pin_1_upper ;
wire [0:0] grid_io_top_8_ccff_tail ;
wire [0:0] grid_io_top_9_bottom_width_0_height_0__pin_1_lower ;
wire [0:0] grid_io_top_9_bottom_width_0_height_0__pin_1_upper ;
wire [0:0] grid_io_top_9_ccff_tail ;
wire [0:19] sb_0__0__0_chanx_right_out ;
wire [0:19] sb_0__0__0_chany_top_out ;
wire [0:0] sb_0__12__0_ccff_tail ;
wire [0:19] sb_0__12__0_chanx_right_out ;
wire [0:19] sb_0__12__0_chany_bottom_out ;
wire [0:0] sb_0__1__0_ccff_tail ;
wire [0:19] sb_0__1__0_chanx_right_out ;
wire [0:19] sb_0__1__0_chany_bottom_out ;
wire [0:19] sb_0__1__0_chany_top_out ;
wire [0:0] sb_0__1__10_ccff_tail ;
wire [0:19] sb_0__1__10_chanx_right_out ;
wire [0:19] sb_0__1__10_chany_bottom_out ;
wire [0:19] sb_0__1__10_chany_top_out ;
wire [0:0] sb_0__1__1_ccff_tail ;
wire [0:19] sb_0__1__1_chanx_right_out ;
wire [0:19] sb_0__1__1_chany_bottom_out ;
wire [0:19] sb_0__1__1_chany_top_out ;
wire [0:0] sb_0__1__2_ccff_tail ;
wire [0:19] sb_0__1__2_chanx_right_out ;
wire [0:19] sb_0__1__2_chany_bottom_out ;
wire [0:19] sb_0__1__2_chany_top_out ;
wire [0:0] sb_0__1__3_ccff_tail ;
wire [0:19] sb_0__1__3_chanx_right_out ;
wire [0:19] sb_0__1__3_chany_bottom_out ;
wire [0:19] sb_0__1__3_chany_top_out ;
wire [0:0] sb_0__1__4_ccff_tail ;
wire [0:19] sb_0__1__4_chanx_right_out ;
wire [0:19] sb_0__1__4_chany_bottom_out ;
wire [0:19] sb_0__1__4_chany_top_out ;
wire [0:0] sb_0__1__5_ccff_tail ;
wire [0:19] sb_0__1__5_chanx_right_out ;
wire [0:19] sb_0__1__5_chany_bottom_out ;
wire [0:19] sb_0__1__5_chany_top_out ;
wire [0:0] sb_0__1__6_ccff_tail ;
wire [0:19] sb_0__1__6_chanx_right_out ;
wire [0:19] sb_0__1__6_chany_bottom_out ;
wire [0:19] sb_0__1__6_chany_top_out ;
wire [0:0] sb_0__1__7_ccff_tail ;
wire [0:19] sb_0__1__7_chanx_right_out ;
wire [0:19] sb_0__1__7_chany_bottom_out ;
wire [0:19] sb_0__1__7_chany_top_out ;
wire [0:0] sb_0__1__8_ccff_tail ;
wire [0:19] sb_0__1__8_chanx_right_out ;
wire [0:19] sb_0__1__8_chany_bottom_out ;
wire [0:19] sb_0__1__8_chany_top_out ;
wire [0:0] sb_0__1__9_ccff_tail ;
wire [0:19] sb_0__1__9_chanx_right_out ;
wire [0:19] sb_0__1__9_chany_bottom_out ;
wire [0:19] sb_0__1__9_chany_top_out ;
wire [0:0] sb_12__0__0_ccff_tail ;
wire [0:19] sb_12__0__0_chanx_left_out ;
wire [0:19] sb_12__0__0_chany_top_out ;
wire [0:0] sb_12__12__0_ccff_tail ;
wire [0:19] sb_12__12__0_chanx_left_out ;
wire [0:19] sb_12__12__0_chany_bottom_out ;
wire [0:0] sb_12__1__0_ccff_tail ;
wire [0:19] sb_12__1__0_chanx_left_out ;
wire [0:19] sb_12__1__0_chany_bottom_out ;
wire [0:19] sb_12__1__0_chany_top_out ;
wire [0:0] sb_12__1__10_ccff_tail ;
wire [0:19] sb_12__1__10_chanx_left_out ;
wire [0:19] sb_12__1__10_chany_bottom_out ;
wire [0:19] sb_12__1__10_chany_top_out ;
wire [0:0] sb_12__1__1_ccff_tail ;
wire [0:19] sb_12__1__1_chanx_left_out ;
wire [0:19] sb_12__1__1_chany_bottom_out ;
wire [0:19] sb_12__1__1_chany_top_out ;
wire [0:0] sb_12__1__2_ccff_tail ;
wire [0:19] sb_12__1__2_chanx_left_out ;
wire [0:19] sb_12__1__2_chany_bottom_out ;
wire [0:19] sb_12__1__2_chany_top_out ;
wire [0:0] sb_12__1__3_ccff_tail ;
wire [0:19] sb_12__1__3_chanx_left_out ;
wire [0:19] sb_12__1__3_chany_bottom_out ;
wire [0:19] sb_12__1__3_chany_top_out ;
wire [0:0] sb_12__1__4_ccff_tail ;
wire [0:19] sb_12__1__4_chanx_left_out ;
wire [0:19] sb_12__1__4_chany_bottom_out ;
wire [0:19] sb_12__1__4_chany_top_out ;
wire [0:0] sb_12__1__5_ccff_tail ;
wire [0:19] sb_12__1__5_chanx_left_out ;
wire [0:19] sb_12__1__5_chany_bottom_out ;
wire [0:19] sb_12__1__5_chany_top_out ;
wire [0:0] sb_12__1__6_ccff_tail ;
wire [0:19] sb_12__1__6_chanx_left_out ;
wire [0:19] sb_12__1__6_chany_bottom_out ;
wire [0:19] sb_12__1__6_chany_top_out ;
wire [0:0] sb_12__1__7_ccff_tail ;
wire [0:19] sb_12__1__7_chanx_left_out ;
wire [0:19] sb_12__1__7_chany_bottom_out ;
wire [0:19] sb_12__1__7_chany_top_out ;
wire [0:0] sb_12__1__8_ccff_tail ;
wire [0:19] sb_12__1__8_chanx_left_out ;
wire [0:19] sb_12__1__8_chany_bottom_out ;
wire [0:19] sb_12__1__8_chany_top_out ;
wire [0:0] sb_12__1__9_ccff_tail ;
wire [0:19] sb_12__1__9_chanx_left_out ;
wire [0:19] sb_12__1__9_chany_bottom_out ;
wire [0:19] sb_12__1__9_chany_top_out ;
wire [0:0] sb_1__0__0_ccff_tail ;
wire [0:19] sb_1__0__0_chanx_left_out ;
wire [0:19] sb_1__0__0_chanx_right_out ;
wire [0:19] sb_1__0__0_chany_top_out ;
wire [0:0] sb_1__0__10_ccff_tail ;
wire [0:19] sb_1__0__10_chanx_left_out ;
wire [0:19] sb_1__0__10_chanx_right_out ;
wire [0:19] sb_1__0__10_chany_top_out ;
wire [0:0] sb_1__0__1_ccff_tail ;
wire [0:19] sb_1__0__1_chanx_left_out ;
wire [0:19] sb_1__0__1_chanx_right_out ;
wire [0:19] sb_1__0__1_chany_top_out ;
wire [0:0] sb_1__0__2_ccff_tail ;
wire [0:19] sb_1__0__2_chanx_left_out ;
wire [0:19] sb_1__0__2_chanx_right_out ;
wire [0:19] sb_1__0__2_chany_top_out ;
wire [0:0] sb_1__0__3_ccff_tail ;
wire [0:19] sb_1__0__3_chanx_left_out ;
wire [0:19] sb_1__0__3_chanx_right_out ;
wire [0:19] sb_1__0__3_chany_top_out ;
wire [0:0] sb_1__0__4_ccff_tail ;
wire [0:19] sb_1__0__4_chanx_left_out ;
wire [0:19] sb_1__0__4_chanx_right_out ;
wire [0:19] sb_1__0__4_chany_top_out ;
wire [0:0] sb_1__0__5_ccff_tail ;
wire [0:19] sb_1__0__5_chanx_left_out ;
wire [0:19] sb_1__0__5_chanx_right_out ;
wire [0:19] sb_1__0__5_chany_top_out ;
wire [0:0] sb_1__0__6_ccff_tail ;
wire [0:19] sb_1__0__6_chanx_left_out ;
wire [0:19] sb_1__0__6_chanx_right_out ;
wire [0:19] sb_1__0__6_chany_top_out ;
wire [0:0] sb_1__0__7_ccff_tail ;
wire [0:19] sb_1__0__7_chanx_left_out ;
wire [0:19] sb_1__0__7_chanx_right_out ;
wire [0:19] sb_1__0__7_chany_top_out ;
wire [0:0] sb_1__0__8_ccff_tail ;
wire [0:19] sb_1__0__8_chanx_left_out ;
wire [0:19] sb_1__0__8_chanx_right_out ;
wire [0:19] sb_1__0__8_chany_top_out ;
wire [0:0] sb_1__0__9_ccff_tail ;
wire [0:19] sb_1__0__9_chanx_left_out ;
wire [0:19] sb_1__0__9_chanx_right_out ;
wire [0:19] sb_1__0__9_chany_top_out ;
wire [0:0] sb_1__12__0_ccff_tail ;
wire [0:19] sb_1__12__0_chanx_left_out ;
wire [0:19] sb_1__12__0_chanx_right_out ;
wire [0:19] sb_1__12__0_chany_bottom_out ;
wire [0:0] sb_1__12__10_ccff_tail ;
wire [0:19] sb_1__12__10_chanx_left_out ;
wire [0:19] sb_1__12__10_chanx_right_out ;
wire [0:19] sb_1__12__10_chany_bottom_out ;
wire [0:0] sb_1__12__1_ccff_tail ;
wire [0:19] sb_1__12__1_chanx_left_out ;
wire [0:19] sb_1__12__1_chanx_right_out ;
wire [0:19] sb_1__12__1_chany_bottom_out ;
wire [0:0] sb_1__12__2_ccff_tail ;
wire [0:19] sb_1__12__2_chanx_left_out ;
wire [0:19] sb_1__12__2_chanx_right_out ;
wire [0:19] sb_1__12__2_chany_bottom_out ;
wire [0:0] sb_1__12__3_ccff_tail ;
wire [0:19] sb_1__12__3_chanx_left_out ;
wire [0:19] sb_1__12__3_chanx_right_out ;
wire [0:19] sb_1__12__3_chany_bottom_out ;
wire [0:0] sb_1__12__4_ccff_tail ;
wire [0:19] sb_1__12__4_chanx_left_out ;
wire [0:19] sb_1__12__4_chanx_right_out ;
wire [0:19] sb_1__12__4_chany_bottom_out ;
wire [0:0] sb_1__12__5_ccff_tail ;
wire [0:19] sb_1__12__5_chanx_left_out ;
wire [0:19] sb_1__12__5_chanx_right_out ;
wire [0:19] sb_1__12__5_chany_bottom_out ;
wire [0:0] sb_1__12__6_ccff_tail ;
wire [0:19] sb_1__12__6_chanx_left_out ;
wire [0:19] sb_1__12__6_chanx_right_out ;
wire [0:19] sb_1__12__6_chany_bottom_out ;
wire [0:0] sb_1__12__7_ccff_tail ;
wire [0:19] sb_1__12__7_chanx_left_out ;
wire [0:19] sb_1__12__7_chanx_right_out ;
wire [0:19] sb_1__12__7_chany_bottom_out ;
wire [0:0] sb_1__12__8_ccff_tail ;
wire [0:19] sb_1__12__8_chanx_left_out ;
wire [0:19] sb_1__12__8_chanx_right_out ;
wire [0:19] sb_1__12__8_chany_bottom_out ;
wire [0:0] sb_1__12__9_ccff_tail ;
wire [0:19] sb_1__12__9_chanx_left_out ;
wire [0:19] sb_1__12__9_chanx_right_out ;
wire [0:19] sb_1__12__9_chany_bottom_out ;
wire [0:0] sb_1__1__0_ccff_tail ;
wire [0:19] sb_1__1__0_chanx_left_out ;
wire [0:19] sb_1__1__0_chanx_right_out ;
wire [0:19] sb_1__1__0_chany_bottom_out ;
wire [0:19] sb_1__1__0_chany_top_out ;
wire [0:0] sb_1__1__100_ccff_tail ;
wire [0:19] sb_1__1__100_chanx_left_out ;
wire [0:19] sb_1__1__100_chanx_right_out ;
wire [0:19] sb_1__1__100_chany_bottom_out ;
wire [0:19] sb_1__1__100_chany_top_out ;
wire [0:0] sb_1__1__101_ccff_tail ;
wire [0:19] sb_1__1__101_chanx_left_out ;
wire [0:19] sb_1__1__101_chanx_right_out ;
wire [0:19] sb_1__1__101_chany_bottom_out ;
wire [0:19] sb_1__1__101_chany_top_out ;
wire [0:0] sb_1__1__102_ccff_tail ;
wire [0:19] sb_1__1__102_chanx_left_out ;
wire [0:19] sb_1__1__102_chanx_right_out ;
wire [0:19] sb_1__1__102_chany_bottom_out ;
wire [0:19] sb_1__1__102_chany_top_out ;
wire [0:0] sb_1__1__103_ccff_tail ;
wire [0:19] sb_1__1__103_chanx_left_out ;
wire [0:19] sb_1__1__103_chanx_right_out ;
wire [0:19] sb_1__1__103_chany_bottom_out ;
wire [0:19] sb_1__1__103_chany_top_out ;
wire [0:0] sb_1__1__104_ccff_tail ;
wire [0:19] sb_1__1__104_chanx_left_out ;
wire [0:19] sb_1__1__104_chanx_right_out ;
wire [0:19] sb_1__1__104_chany_bottom_out ;
wire [0:19] sb_1__1__104_chany_top_out ;
wire [0:0] sb_1__1__105_ccff_tail ;
wire [0:19] sb_1__1__105_chanx_left_out ;
wire [0:19] sb_1__1__105_chanx_right_out ;
wire [0:19] sb_1__1__105_chany_bottom_out ;
wire [0:19] sb_1__1__105_chany_top_out ;
wire [0:0] sb_1__1__106_ccff_tail ;
wire [0:19] sb_1__1__106_chanx_left_out ;
wire [0:19] sb_1__1__106_chanx_right_out ;
wire [0:19] sb_1__1__106_chany_bottom_out ;
wire [0:19] sb_1__1__106_chany_top_out ;
wire [0:0] sb_1__1__107_ccff_tail ;
wire [0:19] sb_1__1__107_chanx_left_out ;
wire [0:19] sb_1__1__107_chanx_right_out ;
wire [0:19] sb_1__1__107_chany_bottom_out ;
wire [0:19] sb_1__1__107_chany_top_out ;
wire [0:0] sb_1__1__108_ccff_tail ;
wire [0:19] sb_1__1__108_chanx_left_out ;
wire [0:19] sb_1__1__108_chanx_right_out ;
wire [0:19] sb_1__1__108_chany_bottom_out ;
wire [0:19] sb_1__1__108_chany_top_out ;
wire [0:0] sb_1__1__109_ccff_tail ;
wire [0:19] sb_1__1__109_chanx_left_out ;
wire [0:19] sb_1__1__109_chanx_right_out ;
wire [0:19] sb_1__1__109_chany_bottom_out ;
wire [0:19] sb_1__1__109_chany_top_out ;
wire [0:0] sb_1__1__10_ccff_tail ;
wire [0:19] sb_1__1__10_chanx_left_out ;
wire [0:19] sb_1__1__10_chanx_right_out ;
wire [0:19] sb_1__1__10_chany_bottom_out ;
wire [0:19] sb_1__1__10_chany_top_out ;
wire [0:0] sb_1__1__110_ccff_tail ;
wire [0:19] sb_1__1__110_chanx_left_out ;
wire [0:19] sb_1__1__110_chanx_right_out ;
wire [0:19] sb_1__1__110_chany_bottom_out ;
wire [0:19] sb_1__1__110_chany_top_out ;
wire [0:0] sb_1__1__111_ccff_tail ;
wire [0:19] sb_1__1__111_chanx_left_out ;
wire [0:19] sb_1__1__111_chanx_right_out ;
wire [0:19] sb_1__1__111_chany_bottom_out ;
wire [0:19] sb_1__1__111_chany_top_out ;
wire [0:0] sb_1__1__112_ccff_tail ;
wire [0:19] sb_1__1__112_chanx_left_out ;
wire [0:19] sb_1__1__112_chanx_right_out ;
wire [0:19] sb_1__1__112_chany_bottom_out ;
wire [0:19] sb_1__1__112_chany_top_out ;
wire [0:0] sb_1__1__113_ccff_tail ;
wire [0:19] sb_1__1__113_chanx_left_out ;
wire [0:19] sb_1__1__113_chanx_right_out ;
wire [0:19] sb_1__1__113_chany_bottom_out ;
wire [0:19] sb_1__1__113_chany_top_out ;
wire [0:0] sb_1__1__114_ccff_tail ;
wire [0:19] sb_1__1__114_chanx_left_out ;
wire [0:19] sb_1__1__114_chanx_right_out ;
wire [0:19] sb_1__1__114_chany_bottom_out ;
wire [0:19] sb_1__1__114_chany_top_out ;
wire [0:0] sb_1__1__115_ccff_tail ;
wire [0:19] sb_1__1__115_chanx_left_out ;
wire [0:19] sb_1__1__115_chanx_right_out ;
wire [0:19] sb_1__1__115_chany_bottom_out ;
wire [0:19] sb_1__1__115_chany_top_out ;
wire [0:0] sb_1__1__116_ccff_tail ;
wire [0:19] sb_1__1__116_chanx_left_out ;
wire [0:19] sb_1__1__116_chanx_right_out ;
wire [0:19] sb_1__1__116_chany_bottom_out ;
wire [0:19] sb_1__1__116_chany_top_out ;
wire [0:0] sb_1__1__117_ccff_tail ;
wire [0:19] sb_1__1__117_chanx_left_out ;
wire [0:19] sb_1__1__117_chanx_right_out ;
wire [0:19] sb_1__1__117_chany_bottom_out ;
wire [0:19] sb_1__1__117_chany_top_out ;
wire [0:0] sb_1__1__118_ccff_tail ;
wire [0:19] sb_1__1__118_chanx_left_out ;
wire [0:19] sb_1__1__118_chanx_right_out ;
wire [0:19] sb_1__1__118_chany_bottom_out ;
wire [0:19] sb_1__1__118_chany_top_out ;
wire [0:0] sb_1__1__119_ccff_tail ;
wire [0:19] sb_1__1__119_chanx_left_out ;
wire [0:19] sb_1__1__119_chanx_right_out ;
wire [0:19] sb_1__1__119_chany_bottom_out ;
wire [0:19] sb_1__1__119_chany_top_out ;
wire [0:0] sb_1__1__11_ccff_tail ;
wire [0:19] sb_1__1__11_chanx_left_out ;
wire [0:19] sb_1__1__11_chanx_right_out ;
wire [0:19] sb_1__1__11_chany_bottom_out ;
wire [0:19] sb_1__1__11_chany_top_out ;
wire [0:0] sb_1__1__120_ccff_tail ;
wire [0:19] sb_1__1__120_chanx_left_out ;
wire [0:19] sb_1__1__120_chanx_right_out ;
wire [0:19] sb_1__1__120_chany_bottom_out ;
wire [0:19] sb_1__1__120_chany_top_out ;
wire [0:0] sb_1__1__12_ccff_tail ;
wire [0:19] sb_1__1__12_chanx_left_out ;
wire [0:19] sb_1__1__12_chanx_right_out ;
wire [0:19] sb_1__1__12_chany_bottom_out ;
wire [0:19] sb_1__1__12_chany_top_out ;
wire [0:0] sb_1__1__13_ccff_tail ;
wire [0:19] sb_1__1__13_chanx_left_out ;
wire [0:19] sb_1__1__13_chanx_right_out ;
wire [0:19] sb_1__1__13_chany_bottom_out ;
wire [0:19] sb_1__1__13_chany_top_out ;
wire [0:0] sb_1__1__14_ccff_tail ;
wire [0:19] sb_1__1__14_chanx_left_out ;
wire [0:19] sb_1__1__14_chanx_right_out ;
wire [0:19] sb_1__1__14_chany_bottom_out ;
wire [0:19] sb_1__1__14_chany_top_out ;
wire [0:0] sb_1__1__15_ccff_tail ;
wire [0:19] sb_1__1__15_chanx_left_out ;
wire [0:19] sb_1__1__15_chanx_right_out ;
wire [0:19] sb_1__1__15_chany_bottom_out ;
wire [0:19] sb_1__1__15_chany_top_out ;
wire [0:0] sb_1__1__16_ccff_tail ;
wire [0:19] sb_1__1__16_chanx_left_out ;
wire [0:19] sb_1__1__16_chanx_right_out ;
wire [0:19] sb_1__1__16_chany_bottom_out ;
wire [0:19] sb_1__1__16_chany_top_out ;
wire [0:0] sb_1__1__17_ccff_tail ;
wire [0:19] sb_1__1__17_chanx_left_out ;
wire [0:19] sb_1__1__17_chanx_right_out ;
wire [0:19] sb_1__1__17_chany_bottom_out ;
wire [0:19] sb_1__1__17_chany_top_out ;
wire [0:0] sb_1__1__18_ccff_tail ;
wire [0:19] sb_1__1__18_chanx_left_out ;
wire [0:19] sb_1__1__18_chanx_right_out ;
wire [0:19] sb_1__1__18_chany_bottom_out ;
wire [0:19] sb_1__1__18_chany_top_out ;
wire [0:0] sb_1__1__19_ccff_tail ;
wire [0:19] sb_1__1__19_chanx_left_out ;
wire [0:19] sb_1__1__19_chanx_right_out ;
wire [0:19] sb_1__1__19_chany_bottom_out ;
wire [0:19] sb_1__1__19_chany_top_out ;
wire [0:0] sb_1__1__1_ccff_tail ;
wire [0:19] sb_1__1__1_chanx_left_out ;
wire [0:19] sb_1__1__1_chanx_right_out ;
wire [0:19] sb_1__1__1_chany_bottom_out ;
wire [0:19] sb_1__1__1_chany_top_out ;
wire [0:0] sb_1__1__20_ccff_tail ;
wire [0:19] sb_1__1__20_chanx_left_out ;
wire [0:19] sb_1__1__20_chanx_right_out ;
wire [0:19] sb_1__1__20_chany_bottom_out ;
wire [0:19] sb_1__1__20_chany_top_out ;
wire [0:0] sb_1__1__21_ccff_tail ;
wire [0:19] sb_1__1__21_chanx_left_out ;
wire [0:19] sb_1__1__21_chanx_right_out ;
wire [0:19] sb_1__1__21_chany_bottom_out ;
wire [0:19] sb_1__1__21_chany_top_out ;
wire [0:0] sb_1__1__22_ccff_tail ;
wire [0:19] sb_1__1__22_chanx_left_out ;
wire [0:19] sb_1__1__22_chanx_right_out ;
wire [0:19] sb_1__1__22_chany_bottom_out ;
wire [0:19] sb_1__1__22_chany_top_out ;
wire [0:0] sb_1__1__23_ccff_tail ;
wire [0:19] sb_1__1__23_chanx_left_out ;
wire [0:19] sb_1__1__23_chanx_right_out ;
wire [0:19] sb_1__1__23_chany_bottom_out ;
wire [0:19] sb_1__1__23_chany_top_out ;
wire [0:0] sb_1__1__24_ccff_tail ;
wire [0:19] sb_1__1__24_chanx_left_out ;
wire [0:19] sb_1__1__24_chanx_right_out ;
wire [0:19] sb_1__1__24_chany_bottom_out ;
wire [0:19] sb_1__1__24_chany_top_out ;
wire [0:0] sb_1__1__25_ccff_tail ;
wire [0:19] sb_1__1__25_chanx_left_out ;
wire [0:19] sb_1__1__25_chanx_right_out ;
wire [0:19] sb_1__1__25_chany_bottom_out ;
wire [0:19] sb_1__1__25_chany_top_out ;
wire [0:0] sb_1__1__26_ccff_tail ;
wire [0:19] sb_1__1__26_chanx_left_out ;
wire [0:19] sb_1__1__26_chanx_right_out ;
wire [0:19] sb_1__1__26_chany_bottom_out ;
wire [0:19] sb_1__1__26_chany_top_out ;
wire [0:0] sb_1__1__27_ccff_tail ;
wire [0:19] sb_1__1__27_chanx_left_out ;
wire [0:19] sb_1__1__27_chanx_right_out ;
wire [0:19] sb_1__1__27_chany_bottom_out ;
wire [0:19] sb_1__1__27_chany_top_out ;
wire [0:0] sb_1__1__28_ccff_tail ;
wire [0:19] sb_1__1__28_chanx_left_out ;
wire [0:19] sb_1__1__28_chanx_right_out ;
wire [0:19] sb_1__1__28_chany_bottom_out ;
wire [0:19] sb_1__1__28_chany_top_out ;
wire [0:0] sb_1__1__29_ccff_tail ;
wire [0:19] sb_1__1__29_chanx_left_out ;
wire [0:19] sb_1__1__29_chanx_right_out ;
wire [0:19] sb_1__1__29_chany_bottom_out ;
wire [0:19] sb_1__1__29_chany_top_out ;
wire [0:0] sb_1__1__2_ccff_tail ;
wire [0:19] sb_1__1__2_chanx_left_out ;
wire [0:19] sb_1__1__2_chanx_right_out ;
wire [0:19] sb_1__1__2_chany_bottom_out ;
wire [0:19] sb_1__1__2_chany_top_out ;
wire [0:0] sb_1__1__30_ccff_tail ;
wire [0:19] sb_1__1__30_chanx_left_out ;
wire [0:19] sb_1__1__30_chanx_right_out ;
wire [0:19] sb_1__1__30_chany_bottom_out ;
wire [0:19] sb_1__1__30_chany_top_out ;
wire [0:0] sb_1__1__31_ccff_tail ;
wire [0:19] sb_1__1__31_chanx_left_out ;
wire [0:19] sb_1__1__31_chanx_right_out ;
wire [0:19] sb_1__1__31_chany_bottom_out ;
wire [0:19] sb_1__1__31_chany_top_out ;
wire [0:0] sb_1__1__32_ccff_tail ;
wire [0:19] sb_1__1__32_chanx_left_out ;
wire [0:19] sb_1__1__32_chanx_right_out ;
wire [0:19] sb_1__1__32_chany_bottom_out ;
wire [0:19] sb_1__1__32_chany_top_out ;
wire [0:0] sb_1__1__33_ccff_tail ;
wire [0:19] sb_1__1__33_chanx_left_out ;
wire [0:19] sb_1__1__33_chanx_right_out ;
wire [0:19] sb_1__1__33_chany_bottom_out ;
wire [0:19] sb_1__1__33_chany_top_out ;
wire [0:0] sb_1__1__34_ccff_tail ;
wire [0:19] sb_1__1__34_chanx_left_out ;
wire [0:19] sb_1__1__34_chanx_right_out ;
wire [0:19] sb_1__1__34_chany_bottom_out ;
wire [0:19] sb_1__1__34_chany_top_out ;
wire [0:0] sb_1__1__35_ccff_tail ;
wire [0:19] sb_1__1__35_chanx_left_out ;
wire [0:19] sb_1__1__35_chanx_right_out ;
wire [0:19] sb_1__1__35_chany_bottom_out ;
wire [0:19] sb_1__1__35_chany_top_out ;
wire [0:0] sb_1__1__36_ccff_tail ;
wire [0:19] sb_1__1__36_chanx_left_out ;
wire [0:19] sb_1__1__36_chanx_right_out ;
wire [0:19] sb_1__1__36_chany_bottom_out ;
wire [0:19] sb_1__1__36_chany_top_out ;
wire [0:0] sb_1__1__37_ccff_tail ;
wire [0:19] sb_1__1__37_chanx_left_out ;
wire [0:19] sb_1__1__37_chanx_right_out ;
wire [0:19] sb_1__1__37_chany_bottom_out ;
wire [0:19] sb_1__1__37_chany_top_out ;
wire [0:0] sb_1__1__38_ccff_tail ;
wire [0:19] sb_1__1__38_chanx_left_out ;
wire [0:19] sb_1__1__38_chanx_right_out ;
wire [0:19] sb_1__1__38_chany_bottom_out ;
wire [0:19] sb_1__1__38_chany_top_out ;
wire [0:0] sb_1__1__39_ccff_tail ;
wire [0:19] sb_1__1__39_chanx_left_out ;
wire [0:19] sb_1__1__39_chanx_right_out ;
wire [0:19] sb_1__1__39_chany_bottom_out ;
wire [0:19] sb_1__1__39_chany_top_out ;
wire [0:0] sb_1__1__3_ccff_tail ;
wire [0:19] sb_1__1__3_chanx_left_out ;
wire [0:19] sb_1__1__3_chanx_right_out ;
wire [0:19] sb_1__1__3_chany_bottom_out ;
wire [0:19] sb_1__1__3_chany_top_out ;
wire [0:0] sb_1__1__40_ccff_tail ;
wire [0:19] sb_1__1__40_chanx_left_out ;
wire [0:19] sb_1__1__40_chanx_right_out ;
wire [0:19] sb_1__1__40_chany_bottom_out ;
wire [0:19] sb_1__1__40_chany_top_out ;
wire [0:0] sb_1__1__41_ccff_tail ;
wire [0:19] sb_1__1__41_chanx_left_out ;
wire [0:19] sb_1__1__41_chanx_right_out ;
wire [0:19] sb_1__1__41_chany_bottom_out ;
wire [0:19] sb_1__1__41_chany_top_out ;
wire [0:0] sb_1__1__42_ccff_tail ;
wire [0:19] sb_1__1__42_chanx_left_out ;
wire [0:19] sb_1__1__42_chanx_right_out ;
wire [0:19] sb_1__1__42_chany_bottom_out ;
wire [0:19] sb_1__1__42_chany_top_out ;
wire [0:0] sb_1__1__43_ccff_tail ;
wire [0:19] sb_1__1__43_chanx_left_out ;
wire [0:19] sb_1__1__43_chanx_right_out ;
wire [0:19] sb_1__1__43_chany_bottom_out ;
wire [0:19] sb_1__1__43_chany_top_out ;
wire [0:0] sb_1__1__44_ccff_tail ;
wire [0:19] sb_1__1__44_chanx_left_out ;
wire [0:19] sb_1__1__44_chanx_right_out ;
wire [0:19] sb_1__1__44_chany_bottom_out ;
wire [0:19] sb_1__1__44_chany_top_out ;
wire [0:0] sb_1__1__45_ccff_tail ;
wire [0:19] sb_1__1__45_chanx_left_out ;
wire [0:19] sb_1__1__45_chanx_right_out ;
wire [0:19] sb_1__1__45_chany_bottom_out ;
wire [0:19] sb_1__1__45_chany_top_out ;
wire [0:0] sb_1__1__46_ccff_tail ;
wire [0:19] sb_1__1__46_chanx_left_out ;
wire [0:19] sb_1__1__46_chanx_right_out ;
wire [0:19] sb_1__1__46_chany_bottom_out ;
wire [0:19] sb_1__1__46_chany_top_out ;
wire [0:0] sb_1__1__47_ccff_tail ;
wire [0:19] sb_1__1__47_chanx_left_out ;
wire [0:19] sb_1__1__47_chanx_right_out ;
wire [0:19] sb_1__1__47_chany_bottom_out ;
wire [0:19] sb_1__1__47_chany_top_out ;
wire [0:0] sb_1__1__48_ccff_tail ;
wire [0:19] sb_1__1__48_chanx_left_out ;
wire [0:19] sb_1__1__48_chanx_right_out ;
wire [0:19] sb_1__1__48_chany_bottom_out ;
wire [0:19] sb_1__1__48_chany_top_out ;
wire [0:0] sb_1__1__49_ccff_tail ;
wire [0:19] sb_1__1__49_chanx_left_out ;
wire [0:19] sb_1__1__49_chanx_right_out ;
wire [0:19] sb_1__1__49_chany_bottom_out ;
wire [0:19] sb_1__1__49_chany_top_out ;
wire [0:0] sb_1__1__4_ccff_tail ;
wire [0:19] sb_1__1__4_chanx_left_out ;
wire [0:19] sb_1__1__4_chanx_right_out ;
wire [0:19] sb_1__1__4_chany_bottom_out ;
wire [0:19] sb_1__1__4_chany_top_out ;
wire [0:0] sb_1__1__50_ccff_tail ;
wire [0:19] sb_1__1__50_chanx_left_out ;
wire [0:19] sb_1__1__50_chanx_right_out ;
wire [0:19] sb_1__1__50_chany_bottom_out ;
wire [0:19] sb_1__1__50_chany_top_out ;
wire [0:0] sb_1__1__51_ccff_tail ;
wire [0:19] sb_1__1__51_chanx_left_out ;
wire [0:19] sb_1__1__51_chanx_right_out ;
wire [0:19] sb_1__1__51_chany_bottom_out ;
wire [0:19] sb_1__1__51_chany_top_out ;
wire [0:0] sb_1__1__52_ccff_tail ;
wire [0:19] sb_1__1__52_chanx_left_out ;
wire [0:19] sb_1__1__52_chanx_right_out ;
wire [0:19] sb_1__1__52_chany_bottom_out ;
wire [0:19] sb_1__1__52_chany_top_out ;
wire [0:0] sb_1__1__53_ccff_tail ;
wire [0:19] sb_1__1__53_chanx_left_out ;
wire [0:19] sb_1__1__53_chanx_right_out ;
wire [0:19] sb_1__1__53_chany_bottom_out ;
wire [0:19] sb_1__1__53_chany_top_out ;
wire [0:0] sb_1__1__54_ccff_tail ;
wire [0:19] sb_1__1__54_chanx_left_out ;
wire [0:19] sb_1__1__54_chanx_right_out ;
wire [0:19] sb_1__1__54_chany_bottom_out ;
wire [0:19] sb_1__1__54_chany_top_out ;
wire [0:0] sb_1__1__55_ccff_tail ;
wire [0:19] sb_1__1__55_chanx_left_out ;
wire [0:19] sb_1__1__55_chanx_right_out ;
wire [0:19] sb_1__1__55_chany_bottom_out ;
wire [0:19] sb_1__1__55_chany_top_out ;
wire [0:0] sb_1__1__56_ccff_tail ;
wire [0:19] sb_1__1__56_chanx_left_out ;
wire [0:19] sb_1__1__56_chanx_right_out ;
wire [0:19] sb_1__1__56_chany_bottom_out ;
wire [0:19] sb_1__1__56_chany_top_out ;
wire [0:0] sb_1__1__57_ccff_tail ;
wire [0:19] sb_1__1__57_chanx_left_out ;
wire [0:19] sb_1__1__57_chanx_right_out ;
wire [0:19] sb_1__1__57_chany_bottom_out ;
wire [0:19] sb_1__1__57_chany_top_out ;
wire [0:0] sb_1__1__58_ccff_tail ;
wire [0:19] sb_1__1__58_chanx_left_out ;
wire [0:19] sb_1__1__58_chanx_right_out ;
wire [0:19] sb_1__1__58_chany_bottom_out ;
wire [0:19] sb_1__1__58_chany_top_out ;
wire [0:0] sb_1__1__59_ccff_tail ;
wire [0:19] sb_1__1__59_chanx_left_out ;
wire [0:19] sb_1__1__59_chanx_right_out ;
wire [0:19] sb_1__1__59_chany_bottom_out ;
wire [0:19] sb_1__1__59_chany_top_out ;
wire [0:0] sb_1__1__5_ccff_tail ;
wire [0:19] sb_1__1__5_chanx_left_out ;
wire [0:19] sb_1__1__5_chanx_right_out ;
wire [0:19] sb_1__1__5_chany_bottom_out ;
wire [0:19] sb_1__1__5_chany_top_out ;
wire [0:0] sb_1__1__60_ccff_tail ;
wire [0:19] sb_1__1__60_chanx_left_out ;
wire [0:19] sb_1__1__60_chanx_right_out ;
wire [0:19] sb_1__1__60_chany_bottom_out ;
wire [0:19] sb_1__1__60_chany_top_out ;
wire [0:0] sb_1__1__61_ccff_tail ;
wire [0:19] sb_1__1__61_chanx_left_out ;
wire [0:19] sb_1__1__61_chanx_right_out ;
wire [0:19] sb_1__1__61_chany_bottom_out ;
wire [0:19] sb_1__1__61_chany_top_out ;
wire [0:0] sb_1__1__62_ccff_tail ;
wire [0:19] sb_1__1__62_chanx_left_out ;
wire [0:19] sb_1__1__62_chanx_right_out ;
wire [0:19] sb_1__1__62_chany_bottom_out ;
wire [0:19] sb_1__1__62_chany_top_out ;
wire [0:0] sb_1__1__63_ccff_tail ;
wire [0:19] sb_1__1__63_chanx_left_out ;
wire [0:19] sb_1__1__63_chanx_right_out ;
wire [0:19] sb_1__1__63_chany_bottom_out ;
wire [0:19] sb_1__1__63_chany_top_out ;
wire [0:0] sb_1__1__64_ccff_tail ;
wire [0:19] sb_1__1__64_chanx_left_out ;
wire [0:19] sb_1__1__64_chanx_right_out ;
wire [0:19] sb_1__1__64_chany_bottom_out ;
wire [0:19] sb_1__1__64_chany_top_out ;
wire [0:0] sb_1__1__65_ccff_tail ;
wire [0:19] sb_1__1__65_chanx_left_out ;
wire [0:19] sb_1__1__65_chanx_right_out ;
wire [0:19] sb_1__1__65_chany_bottom_out ;
wire [0:19] sb_1__1__65_chany_top_out ;
wire [0:0] sb_1__1__66_ccff_tail ;
wire [0:19] sb_1__1__66_chanx_left_out ;
wire [0:19] sb_1__1__66_chanx_right_out ;
wire [0:19] sb_1__1__66_chany_bottom_out ;
wire [0:19] sb_1__1__66_chany_top_out ;
wire [0:0] sb_1__1__67_ccff_tail ;
wire [0:19] sb_1__1__67_chanx_left_out ;
wire [0:19] sb_1__1__67_chanx_right_out ;
wire [0:19] sb_1__1__67_chany_bottom_out ;
wire [0:19] sb_1__1__67_chany_top_out ;
wire [0:0] sb_1__1__68_ccff_tail ;
wire [0:19] sb_1__1__68_chanx_left_out ;
wire [0:19] sb_1__1__68_chanx_right_out ;
wire [0:19] sb_1__1__68_chany_bottom_out ;
wire [0:19] sb_1__1__68_chany_top_out ;
wire [0:0] sb_1__1__69_ccff_tail ;
wire [0:19] sb_1__1__69_chanx_left_out ;
wire [0:19] sb_1__1__69_chanx_right_out ;
wire [0:19] sb_1__1__69_chany_bottom_out ;
wire [0:19] sb_1__1__69_chany_top_out ;
wire [0:0] sb_1__1__6_ccff_tail ;
wire [0:19] sb_1__1__6_chanx_left_out ;
wire [0:19] sb_1__1__6_chanx_right_out ;
wire [0:19] sb_1__1__6_chany_bottom_out ;
wire [0:19] sb_1__1__6_chany_top_out ;
wire [0:0] sb_1__1__70_ccff_tail ;
wire [0:19] sb_1__1__70_chanx_left_out ;
wire [0:19] sb_1__1__70_chanx_right_out ;
wire [0:19] sb_1__1__70_chany_bottom_out ;
wire [0:19] sb_1__1__70_chany_top_out ;
wire [0:0] sb_1__1__71_ccff_tail ;
wire [0:19] sb_1__1__71_chanx_left_out ;
wire [0:19] sb_1__1__71_chanx_right_out ;
wire [0:19] sb_1__1__71_chany_bottom_out ;
wire [0:19] sb_1__1__71_chany_top_out ;
wire [0:0] sb_1__1__72_ccff_tail ;
wire [0:19] sb_1__1__72_chanx_left_out ;
wire [0:19] sb_1__1__72_chanx_right_out ;
wire [0:19] sb_1__1__72_chany_bottom_out ;
wire [0:19] sb_1__1__72_chany_top_out ;
wire [0:0] sb_1__1__73_ccff_tail ;
wire [0:19] sb_1__1__73_chanx_left_out ;
wire [0:19] sb_1__1__73_chanx_right_out ;
wire [0:19] sb_1__1__73_chany_bottom_out ;
wire [0:19] sb_1__1__73_chany_top_out ;
wire [0:0] sb_1__1__74_ccff_tail ;
wire [0:19] sb_1__1__74_chanx_left_out ;
wire [0:19] sb_1__1__74_chanx_right_out ;
wire [0:19] sb_1__1__74_chany_bottom_out ;
wire [0:19] sb_1__1__74_chany_top_out ;
wire [0:0] sb_1__1__75_ccff_tail ;
wire [0:19] sb_1__1__75_chanx_left_out ;
wire [0:19] sb_1__1__75_chanx_right_out ;
wire [0:19] sb_1__1__75_chany_bottom_out ;
wire [0:19] sb_1__1__75_chany_top_out ;
wire [0:0] sb_1__1__76_ccff_tail ;
wire [0:19] sb_1__1__76_chanx_left_out ;
wire [0:19] sb_1__1__76_chanx_right_out ;
wire [0:19] sb_1__1__76_chany_bottom_out ;
wire [0:19] sb_1__1__76_chany_top_out ;
wire [0:0] sb_1__1__77_ccff_tail ;
wire [0:19] sb_1__1__77_chanx_left_out ;
wire [0:19] sb_1__1__77_chanx_right_out ;
wire [0:19] sb_1__1__77_chany_bottom_out ;
wire [0:19] sb_1__1__77_chany_top_out ;
wire [0:0] sb_1__1__78_ccff_tail ;
wire [0:19] sb_1__1__78_chanx_left_out ;
wire [0:19] sb_1__1__78_chanx_right_out ;
wire [0:19] sb_1__1__78_chany_bottom_out ;
wire [0:19] sb_1__1__78_chany_top_out ;
wire [0:0] sb_1__1__79_ccff_tail ;
wire [0:19] sb_1__1__79_chanx_left_out ;
wire [0:19] sb_1__1__79_chanx_right_out ;
wire [0:19] sb_1__1__79_chany_bottom_out ;
wire [0:19] sb_1__1__79_chany_top_out ;
wire [0:0] sb_1__1__7_ccff_tail ;
wire [0:19] sb_1__1__7_chanx_left_out ;
wire [0:19] sb_1__1__7_chanx_right_out ;
wire [0:19] sb_1__1__7_chany_bottom_out ;
wire [0:19] sb_1__1__7_chany_top_out ;
wire [0:0] sb_1__1__80_ccff_tail ;
wire [0:19] sb_1__1__80_chanx_left_out ;
wire [0:19] sb_1__1__80_chanx_right_out ;
wire [0:19] sb_1__1__80_chany_bottom_out ;
wire [0:19] sb_1__1__80_chany_top_out ;
wire [0:0] sb_1__1__81_ccff_tail ;
wire [0:19] sb_1__1__81_chanx_left_out ;
wire [0:19] sb_1__1__81_chanx_right_out ;
wire [0:19] sb_1__1__81_chany_bottom_out ;
wire [0:19] sb_1__1__81_chany_top_out ;
wire [0:0] sb_1__1__82_ccff_tail ;
wire [0:19] sb_1__1__82_chanx_left_out ;
wire [0:19] sb_1__1__82_chanx_right_out ;
wire [0:19] sb_1__1__82_chany_bottom_out ;
wire [0:19] sb_1__1__82_chany_top_out ;
wire [0:0] sb_1__1__83_ccff_tail ;
wire [0:19] sb_1__1__83_chanx_left_out ;
wire [0:19] sb_1__1__83_chanx_right_out ;
wire [0:19] sb_1__1__83_chany_bottom_out ;
wire [0:19] sb_1__1__83_chany_top_out ;
wire [0:0] sb_1__1__84_ccff_tail ;
wire [0:19] sb_1__1__84_chanx_left_out ;
wire [0:19] sb_1__1__84_chanx_right_out ;
wire [0:19] sb_1__1__84_chany_bottom_out ;
wire [0:19] sb_1__1__84_chany_top_out ;
wire [0:0] sb_1__1__85_ccff_tail ;
wire [0:19] sb_1__1__85_chanx_left_out ;
wire [0:19] sb_1__1__85_chanx_right_out ;
wire [0:19] sb_1__1__85_chany_bottom_out ;
wire [0:19] sb_1__1__85_chany_top_out ;
wire [0:0] sb_1__1__86_ccff_tail ;
wire [0:19] sb_1__1__86_chanx_left_out ;
wire [0:19] sb_1__1__86_chanx_right_out ;
wire [0:19] sb_1__1__86_chany_bottom_out ;
wire [0:19] sb_1__1__86_chany_top_out ;
wire [0:0] sb_1__1__87_ccff_tail ;
wire [0:19] sb_1__1__87_chanx_left_out ;
wire [0:19] sb_1__1__87_chanx_right_out ;
wire [0:19] sb_1__1__87_chany_bottom_out ;
wire [0:19] sb_1__1__87_chany_top_out ;
wire [0:0] sb_1__1__88_ccff_tail ;
wire [0:19] sb_1__1__88_chanx_left_out ;
wire [0:19] sb_1__1__88_chanx_right_out ;
wire [0:19] sb_1__1__88_chany_bottom_out ;
wire [0:19] sb_1__1__88_chany_top_out ;
wire [0:0] sb_1__1__89_ccff_tail ;
wire [0:19] sb_1__1__89_chanx_left_out ;
wire [0:19] sb_1__1__89_chanx_right_out ;
wire [0:19] sb_1__1__89_chany_bottom_out ;
wire [0:19] sb_1__1__89_chany_top_out ;
wire [0:0] sb_1__1__8_ccff_tail ;
wire [0:19] sb_1__1__8_chanx_left_out ;
wire [0:19] sb_1__1__8_chanx_right_out ;
wire [0:19] sb_1__1__8_chany_bottom_out ;
wire [0:19] sb_1__1__8_chany_top_out ;
wire [0:0] sb_1__1__90_ccff_tail ;
wire [0:19] sb_1__1__90_chanx_left_out ;
wire [0:19] sb_1__1__90_chanx_right_out ;
wire [0:19] sb_1__1__90_chany_bottom_out ;
wire [0:19] sb_1__1__90_chany_top_out ;
wire [0:0] sb_1__1__91_ccff_tail ;
wire [0:19] sb_1__1__91_chanx_left_out ;
wire [0:19] sb_1__1__91_chanx_right_out ;
wire [0:19] sb_1__1__91_chany_bottom_out ;
wire [0:19] sb_1__1__91_chany_top_out ;
wire [0:0] sb_1__1__92_ccff_tail ;
wire [0:19] sb_1__1__92_chanx_left_out ;
wire [0:19] sb_1__1__92_chanx_right_out ;
wire [0:19] sb_1__1__92_chany_bottom_out ;
wire [0:19] sb_1__1__92_chany_top_out ;
wire [0:0] sb_1__1__93_ccff_tail ;
wire [0:19] sb_1__1__93_chanx_left_out ;
wire [0:19] sb_1__1__93_chanx_right_out ;
wire [0:19] sb_1__1__93_chany_bottom_out ;
wire [0:19] sb_1__1__93_chany_top_out ;
wire [0:0] sb_1__1__94_ccff_tail ;
wire [0:19] sb_1__1__94_chanx_left_out ;
wire [0:19] sb_1__1__94_chanx_right_out ;
wire [0:19] sb_1__1__94_chany_bottom_out ;
wire [0:19] sb_1__1__94_chany_top_out ;
wire [0:0] sb_1__1__95_ccff_tail ;
wire [0:19] sb_1__1__95_chanx_left_out ;
wire [0:19] sb_1__1__95_chanx_right_out ;
wire [0:19] sb_1__1__95_chany_bottom_out ;
wire [0:19] sb_1__1__95_chany_top_out ;
wire [0:0] sb_1__1__96_ccff_tail ;
wire [0:19] sb_1__1__96_chanx_left_out ;
wire [0:19] sb_1__1__96_chanx_right_out ;
wire [0:19] sb_1__1__96_chany_bottom_out ;
wire [0:19] sb_1__1__96_chany_top_out ;
wire [0:0] sb_1__1__97_ccff_tail ;
wire [0:19] sb_1__1__97_chanx_left_out ;
wire [0:19] sb_1__1__97_chanx_right_out ;
wire [0:19] sb_1__1__97_chany_bottom_out ;
wire [0:19] sb_1__1__97_chany_top_out ;
wire [0:0] sb_1__1__98_ccff_tail ;
wire [0:19] sb_1__1__98_chanx_left_out ;
wire [0:19] sb_1__1__98_chanx_right_out ;
wire [0:19] sb_1__1__98_chany_bottom_out ;
wire [0:19] sb_1__1__98_chany_top_out ;
wire [0:0] sb_1__1__99_ccff_tail ;
wire [0:19] sb_1__1__99_chanx_left_out ;
wire [0:19] sb_1__1__99_chanx_right_out ;
wire [0:19] sb_1__1__99_chany_bottom_out ;
wire [0:19] sb_1__1__99_chany_top_out ;
wire [0:0] sb_1__1__9_ccff_tail ;
wire [0:19] sb_1__1__9_chanx_left_out ;
wire [0:19] sb_1__1__9_chanx_right_out ;
wire [0:19] sb_1__1__9_chany_bottom_out ;
wire [0:19] sb_1__1__9_chany_top_out ;
//

grid_clb grid_clb_1__1_ (
    .prog_clk ( { ctsbuf_net_4422424 } ) ,
    .Test_en ( { BUF_net_583 } ) ,
    .clk ( { ctsbuf_net_21984 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_0_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_143_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__0_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__0_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__0_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__0_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__0_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__0_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__0_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__0_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__0_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__0_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__0_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__0_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__0_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__0_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__0_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__0_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__0__0_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__0__0_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__0__0_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__0__0_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__0__0_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__0__0_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__0__0_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__0__0_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__0__0_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__0__0_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__0__0_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__0__0_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__0__0_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__0__0_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__0__0_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__0__0_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_0__1__0_right_grid_pin_52_ ) , 
    .ccff_head ( grid_io_left_0_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_0_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_0_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_0_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_0_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_0_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_0_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_0_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_0_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_0_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_0_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_0_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_0_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_0_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_0_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_0_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_0_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_0_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_0_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_0_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_0_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_0_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_0_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_0_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_0_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_0_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_0_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_0_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_0_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_0_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_0_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_0_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_0_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_0_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_0_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_0_ccff_tail ) ) ;
grid_clb grid_clb_1__2_ (
    .prog_clk ( { ctsbuf_net_4842466 } ) ,
    .Test_en ( { BUF_net_582 } ) ,
    .clk ( { ctsbuf_net_21984 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_1_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_144_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__1_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__1_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__1_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__1_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__1_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__1_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__1_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__1_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__1_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__1_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__1_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__1_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__1_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__1_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__1_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__1_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__0_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__0_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__0_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__0_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__0_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__0_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__0_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__0_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__0_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__0_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__0_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__0_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__0_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__0_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__0_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__0_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_0__1__1_right_grid_pin_52_ ) , 
    .ccff_head ( grid_io_left_1_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_1_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_1_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_1_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_1_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_1_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_1_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_1_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_1_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_1_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_1_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_1_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_1_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_1_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_1_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_1_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_1_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_1_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_1_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_1_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_1_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_1_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_1_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_1_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_1_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_1_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_1_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_1_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_1_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_1_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_1_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_1_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_1_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_1_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_1_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_1_ccff_tail ) ) ;
grid_clb grid_clb_1__3_ (
    .prog_clk ( { ctsbuf_net_5172499 } ) ,
    .Test_en ( { BUF_net_581 } ) ,
    .clk ( { ctsbuf_net_51987 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_2_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_145_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__2_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__2_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__2_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__2_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__2_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__2_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__2_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__2_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__2_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__2_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__2_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__2_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__2_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__2_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__2_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__2_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__1_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__1_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__1_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__1_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__1_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__1_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__1_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__1_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__1_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__1_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__1_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__1_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__1_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__1_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__1_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__1_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_0__1__2_right_grid_pin_52_ ) , 
    .ccff_head ( grid_io_left_2_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_2_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_2_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_2_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_2_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_2_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_2_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_2_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_2_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_2_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_2_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_2_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_2_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_2_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_2_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_2_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_2_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_2_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_2_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_2_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_2_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_2_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_2_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_2_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_2_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_2_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_2_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_2_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_2_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_2_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_2_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_2_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_2_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_2_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_2_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_2_ccff_tail ) ) ;
grid_clb grid_clb_1__4_ (
    .prog_clk ( { ctsbuf_net_5452527 } ) ,
    .Test_en ( { BUF_net_580 } ) ,
    .clk ( { ctsbuf_net_51987 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_3_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_146_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__3_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__3_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__3_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__3_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__3_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__3_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__3_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__3_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__3_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__3_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__3_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__3_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__3_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__3_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__3_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__3_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__2_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__2_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__2_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__2_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__2_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__2_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__2_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__2_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__2_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__2_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__2_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__2_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__2_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__2_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__2_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__2_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_0__1__3_right_grid_pin_52_ ) , 
    .ccff_head ( grid_io_left_3_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_3_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_3_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_3_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_3_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_3_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_3_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_3_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_3_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_3_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_3_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_3_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_3_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_3_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_3_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_3_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_3_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_3_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_3_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_3_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_3_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_3_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_3_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_3_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_3_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_3_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_3_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_3_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_3_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_3_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_3_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_3_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_3_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_3_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_3_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_3_ccff_tail ) ) ;
grid_clb grid_clb_1__5_ (
    .prog_clk ( { ctsbuf_net_5652547 } ) ,
    .Test_en ( { BUF_net_579 } ) ,
    .clk ( { ctsbuf_net_101992 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_4_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_147_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__4_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__4_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__4_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__4_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__4_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__4_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__4_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__4_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__4_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__4_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__4_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__4_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__4_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__4_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__4_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__4_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__3_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__3_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__3_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__3_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__3_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__3_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__3_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__3_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__3_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__3_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__3_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__3_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__3_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__3_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__3_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__3_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_0__1__4_right_grid_pin_52_ ) , 
    .ccff_head ( grid_io_left_4_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_4_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_4_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_4_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_4_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_4_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_4_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_4_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_4_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_4_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_4_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_4_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_4_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_4_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_4_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_4_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_4_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_4_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_4_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_4_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_4_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_4_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_4_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_4_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_4_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_4_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_4_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_4_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_4_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_4_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_4_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_4_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_4_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_4_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_4_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_4_ccff_tail ) ) ;
grid_clb grid_clb_1__6_ (
    .prog_clk ( { ctsbuf_net_5782560 } ) ,
    .Test_en ( { BUF_net_578 } ) ,
    .clk ( { ctsbuf_net_101992 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_5_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_148_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__5_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__5_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__5_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__5_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__5_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__5_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__5_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__5_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__5_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__5_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__5_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__5_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__5_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__5_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__5_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__5_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__4_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__4_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__4_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__4_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__4_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__4_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__4_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__4_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__4_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__4_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__4_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__4_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__4_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__4_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__4_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__4_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_0__1__5_right_grid_pin_52_ ) , 
    .ccff_head ( grid_io_left_5_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_5_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_5_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_5_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_5_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_5_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_5_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_5_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_5_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_5_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_5_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_5_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_5_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_5_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_5_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_5_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_5_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_5_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_5_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_5_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_5_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_5_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_5_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_5_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_5_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_5_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_5_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_5_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_5_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_5_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_5_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_5_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_5_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_5_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_5_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_5_ccff_tail ) ) ;
grid_clb grid_clb_1__7_ (
    .prog_clk ( { ctsbuf_net_5812563 } ) ,
    .Test_en ( { BUF_net_577 } ) ,
    .clk ( { ctsbuf_net_151997 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_6_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_149_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__6_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__6_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__6_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__6_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__6_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__6_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__6_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__6_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__6_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__6_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__6_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__6_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__6_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__6_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__6_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__6_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__5_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__5_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__5_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__5_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__5_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__5_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__5_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__5_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__5_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__5_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__5_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__5_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__5_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__5_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__5_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__5_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_0__1__6_right_grid_pin_52_ ) , 
    .ccff_head ( grid_io_left_6_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_6_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_6_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_6_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_6_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_6_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_6_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_6_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_6_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_6_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_6_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_6_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_6_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_6_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_6_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_6_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_6_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_6_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_6_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_6_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_6_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_6_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_6_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_6_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_6_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_6_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_6_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_6_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_6_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_6_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_6_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_6_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_6_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_6_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_6_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_6_ccff_tail ) ) ;
grid_clb grid_clb_1__8_ (
    .prog_clk ( { ctsbuf_net_5722554 } ) ,
    .Test_en ( { BUF_net_576 } ) ,
    .clk ( { ctsbuf_net_151997 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_7_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_150_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__7_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__7_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__7_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__7_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__7_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__7_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__7_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__7_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__7_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__7_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__7_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__7_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__7_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__7_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__7_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__7_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__6_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__6_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__6_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__6_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__6_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__6_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__6_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__6_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__6_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__6_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__6_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__6_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__6_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__6_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__6_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__6_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_0__1__7_right_grid_pin_52_ ) , 
    .ccff_head ( grid_io_left_7_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_7_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_7_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_7_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_7_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_7_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_7_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_7_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_7_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_7_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_7_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_7_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_7_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_7_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_7_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_7_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_7_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_7_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_7_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_7_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_7_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_7_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_7_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_7_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_7_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_7_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_7_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_7_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_7_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_7_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_7_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_7_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_7_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_7_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_7_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_7_ccff_tail ) ) ;
grid_clb grid_clb_1__9_ (
    .prog_clk ( { ctsbuf_net_5562538 } ) ,
    .Test_en ( { BUF_net_575 } ) ,
    .clk ( { ctsbuf_net_202002 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_8_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_151_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__8_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__8_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__8_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__8_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__8_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__8_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__8_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__8_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__8_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__8_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__8_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__8_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__8_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__8_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__8_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__8_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__7_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__7_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__7_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__7_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__7_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__7_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__7_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__7_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__7_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__7_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__7_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__7_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__7_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__7_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__7_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__7_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_0__1__8_right_grid_pin_52_ ) , 
    .ccff_head ( grid_io_left_8_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_8_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_8_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_8_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_8_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_8_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_8_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_8_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_8_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_8_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_8_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_8_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_8_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_8_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_8_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_8_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_8_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_8_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_8_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_8_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_8_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_8_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_8_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_8_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_8_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_8_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_8_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_8_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_8_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_8_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_8_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_8_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_8_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_8_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_8_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_8_ccff_tail ) ) ;
grid_clb grid_clb_1__10_ (
    .prog_clk ( { ctsbuf_net_5322514 } ) ,
    .Test_en ( { BUF_net_574 } ) ,
    .clk ( { ctsbuf_net_202002 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_9_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_152_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__9_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__9_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__9_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__9_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__9_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__9_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__9_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__9_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__9_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__9_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__9_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__9_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__9_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__9_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__9_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__9_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__8_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__8_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__8_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__8_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__8_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__8_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__8_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__8_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__8_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__8_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__8_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__8_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__8_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__8_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__8_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__8_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_0__1__9_right_grid_pin_52_ ) , 
    .ccff_head ( grid_io_left_9_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_9_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_9_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_9_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_9_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_9_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_9_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_9_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_9_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_9_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_9_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_9_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_9_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_9_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_9_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_9_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_9_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_9_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_9_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_9_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_9_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_9_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_9_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_9_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_9_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_9_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_9_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_9_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_9_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_9_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_9_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_9_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_9_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_9_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_9_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_9_ccff_tail ) ) ;
grid_clb grid_clb_1__11_ (
    .prog_clk ( { ctsbuf_net_5032485 } ) ,
    .Test_en ( { BUF_net_573 } ) ,
    .clk ( { ctsbuf_net_252007 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_10_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_153_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__10_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__10_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__10_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__10_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__10_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__10_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__10_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__10_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__10_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__10_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__10_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__10_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__10_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__10_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__10_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__10_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__9_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__9_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__9_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__9_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__9_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__9_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__9_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__9_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__9_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__9_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__9_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__9_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__9_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__9_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__9_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__9_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_0__1__10_right_grid_pin_52_ ) , 
    .ccff_head ( grid_io_left_10_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_10_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_10_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_10_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_10_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_10_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_10_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_10_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_10_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_10_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_10_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_10_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_10_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_10_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_10_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_10_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_10_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_10_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_10_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_10_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_10_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_10_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_10_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_10_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_10_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_10_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_10_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_10_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_10_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_10_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_10_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_10_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_10_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_10_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_10_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_10_ccff_tail ) ) ;
grid_clb grid_clb_1__12_ (
    .prog_clk ( { ctsbuf_net_4652447 } ) ,
    .Test_en ( { BUF_net_572 } ) ,
    .clk ( { ctsbuf_net_252007 } ) ,
    
    .top_width_0_height_0__pin_32_ ( grid_clb_1__12__undriven_top_width_0_height_0__pin_32_ ) , 
    .top_width_0_height_0__pin_33_ ( grid_clb_1__12__undriven_top_width_0_height_0__pin_33_ ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__11_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__11_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__11_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__11_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__11_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__11_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__11_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__11_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__11_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__11_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__11_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__11_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__11_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__11_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__11_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__11_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__10_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__10_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__10_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__10_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__10_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__10_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__10_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__10_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__10_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__10_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__10_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__10_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__10_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__10_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__10_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__10_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_0__1__11_right_grid_pin_52_ ) , 
    .ccff_head ( grid_io_left_11_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_11_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_11_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_11_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_11_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_11_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_11_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_11_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_11_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_11_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_11_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_11_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_11_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_11_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_11_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_11_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_11_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_11_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_11_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_11_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_11_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_11_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_11_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_11_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_11_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_11_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_11_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_11_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_11_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_11_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_11_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_11_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_11_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_11_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_11_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_11_ccff_tail ) ) ;
grid_clb grid_clb_2__1_ (
    .prog_clk ( { ctsbuf_net_3982380 } ) ,
    .Test_en ( { BUF_net_571 } ) ,
    .clk ( { ctsbuf_net_21984 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_11_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_154_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__12_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__12_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__12_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__12_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__12_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__12_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__12_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__12_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__12_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__12_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__12_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__12_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__12_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__12_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__12_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__12_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__0__1_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__0__1_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__0__1_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__0__1_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__0__1_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__0__1_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__0__1_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__0__1_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__0__1_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__0__1_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__0__1_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__0__1_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__0__1_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__0__1_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__0__1_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__0__1_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__0_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__0_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_12_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_12_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_12_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_12_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_12_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_12_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_12_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_12_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_12_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_12_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_12_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_12_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_12_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_12_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_12_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_12_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_12_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_12_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_12_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_12_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_12_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_12_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_12_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_12_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_12_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_12_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_12_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_12_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_12_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_12_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_12_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_12_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_12_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_12_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_12_ccff_tail ) ) ;
grid_clb grid_clb_2__2_ (
    .prog_clk ( { ctsbuf_net_4432425 } ) ,
    .Test_en ( { BUF_net_846 } ) ,
    .clk ( { ctsbuf_net_21984 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_12_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_155_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__13_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__13_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__13_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__13_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__13_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__13_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__13_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__13_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__13_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__13_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__13_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__13_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__13_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__13_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__13_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__13_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__11_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__11_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__11_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__11_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__11_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__11_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__11_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__11_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__11_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__11_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__11_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__11_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__11_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__11_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__11_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__11_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__1_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__1_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_13_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_13_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_13_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_13_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_13_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_13_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_13_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_13_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_13_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_13_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_13_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_13_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_13_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_13_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_13_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_13_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_13_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_13_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_13_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_13_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_13_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_13_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_13_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_13_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_13_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_13_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_13_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_13_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_13_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_13_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_13_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_13_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_13_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_13_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_13_ccff_tail ) ) ;
grid_clb grid_clb_2__3_ (
    .prog_clk ( { ctsbuf_net_4852467 } ) ,
    .Test_en ( { BUF_net_718 } ) ,
    .clk ( { ctsbuf_net_51987 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_13_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_156_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__14_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__14_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__14_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__14_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__14_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__14_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__14_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__14_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__14_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__14_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__14_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__14_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__14_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__14_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__14_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__14_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__12_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__12_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__12_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__12_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__12_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__12_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__12_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__12_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__12_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__12_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__12_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__12_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__12_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__12_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__12_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__12_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__2_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__2_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_14_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_14_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_14_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_14_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_14_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_14_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_14_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_14_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_14_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_14_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_14_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_14_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_14_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_14_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_14_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_14_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_14_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_14_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_14_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_14_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_14_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_14_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_14_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_14_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_14_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_14_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_14_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_14_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_14_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_14_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_14_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_14_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_14_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_14_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_14_ccff_tail ) ) ;
grid_clb grid_clb_2__4_ (
    .prog_clk ( { ctsbuf_net_5182500 } ) ,
    .Test_en ( { BUF_net_720 } ) ,
    .clk ( { ctsbuf_net_51987 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_14_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_157_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__15_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__15_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__15_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__15_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__15_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__15_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__15_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__15_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__15_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__15_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__15_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__15_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__15_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__15_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__15_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__15_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__13_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__13_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__13_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__13_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__13_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__13_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__13_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__13_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__13_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__13_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__13_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__13_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__13_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__13_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__13_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__13_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__3_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__3_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_15_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_15_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_15_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_15_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_15_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_15_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_15_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_15_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_15_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_15_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_15_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_15_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_15_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_15_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_15_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_15_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_15_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_15_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_15_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_15_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_15_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_15_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_15_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_15_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_15_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_15_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_15_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_15_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_15_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_15_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_15_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_15_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_15_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_15_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_15_ccff_tail ) ) ;
grid_clb grid_clb_2__5_ (
    .prog_clk ( { ctsbuf_net_5462528 } ) ,
    .Test_en ( { BUF_net_849 } ) ,
    .clk ( { ctsbuf_net_101992 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_15_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_158_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__16_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__16_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__16_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__16_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__16_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__16_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__16_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__16_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__16_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__16_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__16_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__16_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__16_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__16_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__16_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__16_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__14_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__14_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__14_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__14_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__14_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__14_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__14_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__14_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__14_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__14_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__14_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__14_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__14_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__14_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__14_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__14_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__4_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__4_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_16_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_16_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_16_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_16_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_16_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_16_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_16_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_16_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_16_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_16_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_16_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_16_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_16_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_16_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_16_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_16_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_16_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_16_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_16_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_16_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_16_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_16_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_16_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_16_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_16_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_16_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_16_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_16_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_16_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_16_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_16_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_16_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_16_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_16_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_16_ccff_tail ) ) ;
grid_clb grid_clb_2__6_ (
    .prog_clk ( { ctsbuf_net_5662548 } ) ,
    .Test_en ( { BUF_net_566 } ) ,
    .clk ( { ctsbuf_net_101992 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_16_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_159_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__17_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__17_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__17_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__17_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__17_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__17_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__17_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__17_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__17_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__17_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__17_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__17_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__17_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__17_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__17_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__17_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__15_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__15_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__15_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__15_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__15_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__15_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__15_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__15_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__15_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__15_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__15_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__15_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__15_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__15_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__15_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__15_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__5_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__5_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_17_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_17_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_17_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_17_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_17_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_17_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_17_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_17_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_17_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_17_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_17_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_17_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_17_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_17_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_17_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_17_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_17_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_17_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_17_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_17_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_17_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_17_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_17_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_17_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_17_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_17_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_17_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_17_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_17_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_17_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_17_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_17_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_17_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_17_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_17_ccff_tail ) ) ;
grid_clb grid_clb_2__7_ (
    .prog_clk ( { ctsbuf_net_5732555 } ) ,
    .Test_en ( { BUF_net_851 } ) ,
    .clk ( { ctsbuf_net_151997 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_17_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_160_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__18_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__18_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__18_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__18_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__18_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__18_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__18_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__18_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__18_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__18_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__18_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__18_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__18_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__18_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__18_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__18_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__16_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__16_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__16_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__16_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__16_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__16_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__16_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__16_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__16_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__16_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__16_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__16_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__16_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__16_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__16_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__16_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__6_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__6_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_18_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_18_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_18_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_18_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_18_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_18_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_18_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_18_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_18_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_18_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_18_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_18_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_18_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_18_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_18_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_18_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_18_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_18_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_18_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_18_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_18_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_18_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_18_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_18_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_18_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_18_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_18_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_18_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_18_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_18_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_18_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_18_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_18_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_18_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_18_ccff_tail ) ) ;
grid_clb grid_clb_2__8_ (
    .prog_clk ( { ctsbuf_net_5572539 } ) ,
    .Test_en ( { BUF_net_726 } ) ,
    .clk ( { ctsbuf_net_151997 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_18_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_161_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__19_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__19_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__19_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__19_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__19_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__19_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__19_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__19_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__19_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__19_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__19_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__19_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__19_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__19_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__19_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__19_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__17_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__17_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__17_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__17_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__17_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__17_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__17_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__17_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__17_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__17_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__17_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__17_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__17_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__17_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__17_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__17_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__7_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__7_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_19_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_19_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_19_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_19_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_19_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_19_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_19_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_19_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_19_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_19_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_19_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_19_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_19_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_19_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_19_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_19_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_19_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_19_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_19_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_19_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_19_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_19_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_19_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_19_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_19_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_19_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_19_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_19_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_19_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_19_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_19_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_19_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_19_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_19_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_19_ccff_tail ) ) ;
grid_clb grid_clb_2__9_ (
    .prog_clk ( { ctsbuf_net_5332515 } ) ,
    .Test_en ( { BUF_net_853 } ) ,
    .clk ( { ctsbuf_net_202002 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_19_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_162_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__20_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__20_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__20_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__20_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__20_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__20_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__20_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__20_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__20_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__20_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__20_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__20_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__20_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__20_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__20_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__20_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__18_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__18_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__18_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__18_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__18_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__18_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__18_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__18_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__18_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__18_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__18_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__18_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__18_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__18_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__18_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__18_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__8_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__8_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_20_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_20_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_20_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_20_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_20_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_20_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_20_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_20_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_20_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_20_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_20_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_20_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_20_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_20_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_20_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_20_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_20_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_20_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_20_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_20_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_20_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_20_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_20_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_20_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_20_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_20_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_20_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_20_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_20_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_20_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_20_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_20_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_20_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_20_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_20_ccff_tail ) ) ;
grid_clb grid_clb_2__10_ (
    .prog_clk ( { ctsbuf_net_5042486 } ) ,
    .Test_en ( { BUF_net_730 } ) ,
    .clk ( { ctsbuf_net_202002 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_20_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_163_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__21_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__21_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__21_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__21_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__21_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__21_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__21_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__21_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__21_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__21_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__21_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__21_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__21_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__21_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__21_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__21_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__19_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__19_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__19_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__19_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__19_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__19_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__19_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__19_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__19_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__19_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__19_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__19_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__19_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__19_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__19_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__19_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__9_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__9_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_21_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_21_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_21_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_21_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_21_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_21_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_21_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_21_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_21_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_21_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_21_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_21_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_21_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_21_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_21_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_21_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_21_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_21_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_21_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_21_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_21_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_21_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_21_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_21_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_21_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_21_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_21_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_21_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_21_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_21_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_21_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_21_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_21_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_21_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_21_ccff_tail ) ) ;
grid_clb grid_clb_2__11_ (
    .prog_clk ( { ctsbuf_net_4662448 } ) ,
    .Test_en ( { BUF_net_857 } ) ,
    .clk ( { ctsbuf_net_252007 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_21_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_164_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__22_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__22_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__22_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__22_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__22_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__22_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__22_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__22_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__22_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__22_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__22_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__22_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__22_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__22_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__22_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__22_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__20_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__20_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__20_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__20_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__20_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__20_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__20_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__20_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__20_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__20_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__20_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__20_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__20_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__20_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__20_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__20_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__10_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__10_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_22_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_22_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_22_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_22_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_22_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_22_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_22_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_22_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_22_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_22_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_22_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_22_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_22_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_22_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_22_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_22_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_22_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_22_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_22_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_22_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_22_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_22_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_22_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_22_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_22_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_22_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_22_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_22_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_22_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_22_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_22_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_22_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_22_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_22_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_22_ccff_tail ) ) ;
grid_clb grid_clb_2__12_ (
    .prog_clk ( { ctsbuf_net_4232405 } ) ,
    .Test_en ( { BUF_net_560 } ) ,
    .clk ( { ctsbuf_net_252007 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_132_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_275_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__23_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__23_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__23_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__23_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__23_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__23_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__23_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__23_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__23_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__23_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__23_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__23_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__23_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__23_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__23_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__23_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__21_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__21_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__21_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__21_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__21_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__21_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__21_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__21_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__21_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__21_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__21_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__21_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__21_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__21_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__21_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__21_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__11_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__11_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_23_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_23_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_23_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_23_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_23_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_23_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_23_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_23_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_23_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_23_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_23_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_23_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_23_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_23_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_23_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_23_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_23_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_23_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_23_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_23_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_23_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_23_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_23_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_23_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_23_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_23_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_23_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_23_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_23_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_23_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_23_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_23_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_23_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_23_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_23_ccff_tail ) ) ;
grid_clb grid_clb_3__1_ (
    .prog_clk ( { ctsbuf_net_3552337 } ) ,
    .Test_en ( { BUF_net_559 } ) ,
    .clk ( { ctsbuf_net_21984 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_22_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_165_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__24_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__24_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__24_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__24_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__24_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__24_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__24_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__24_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__24_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__24_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__24_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__24_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__24_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__24_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__24_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__24_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__0__2_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__0__2_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__0__2_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__0__2_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__0__2_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__0__2_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__0__2_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__0__2_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__0__2_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__0__2_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__0__2_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__0__2_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__0__2_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__0__2_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__0__2_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__0__2_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__12_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__12_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_24_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_24_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_24_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_24_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_24_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_24_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_24_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_24_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_24_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_24_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_24_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_24_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_24_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_24_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_24_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_24_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_24_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_24_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_24_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_24_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_24_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_24_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_24_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_24_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_24_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_24_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_24_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_24_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_24_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_24_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_24_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_24_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_24_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_24_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_24_ccff_tail ) ) ;
grid_clb grid_clb_3__2_ (
    .prog_clk ( { ctsbuf_net_3992381 } ) ,
    .Test_en ( { BUF_net_1185 } ) ,
    .clk ( { ctsbuf_net_81990 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_23_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_166_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__25_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__25_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__25_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__25_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__25_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__25_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__25_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__25_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__25_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__25_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__25_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__25_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__25_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__25_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__25_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__25_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__22_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__22_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__22_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__22_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__22_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__22_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__22_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__22_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__22_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__22_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__22_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__22_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__22_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__22_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__22_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__22_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__13_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__13_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_25_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_25_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_25_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_25_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_25_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_25_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_25_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_25_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_25_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_25_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_25_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_25_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_25_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_25_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_25_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_25_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_25_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_25_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_25_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_25_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_25_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_25_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_25_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_25_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_25_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_25_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_25_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_25_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_25_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_25_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_25_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_25_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_25_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_25_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_25_ccff_tail ) ) ;
grid_clb grid_clb_3__3_ (
    .prog_clk ( { ctsbuf_net_4442426 } ) ,
    .Test_en ( { BUF_net_966 } ) ,
    .clk ( { ctsbuf_net_81990 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_24_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_167_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__26_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__26_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__26_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__26_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__26_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__26_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__26_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__26_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__26_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__26_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__26_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__26_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__26_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__26_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__26_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__26_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__23_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__23_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__23_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__23_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__23_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__23_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__23_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__23_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__23_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__23_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__23_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__23_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__23_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__23_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__23_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__23_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__14_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__14_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_26_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_26_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_26_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_26_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_26_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_26_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_26_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_26_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_26_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_26_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_26_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_26_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_26_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_26_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_26_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_26_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_26_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_26_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_26_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_26_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_26_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_26_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_26_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_26_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_26_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_26_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_26_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_26_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_26_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_26_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_26_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_26_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_26_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_26_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_26_ccff_tail ) ) ;
grid_clb grid_clb_3__4_ (
    .prog_clk ( { ctsbuf_net_4862468 } ) ,
    .Test_en ( { BUF_net_968 } ) ,
    .clk ( { ctsbuf_net_121994 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_25_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_168_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__27_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__27_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__27_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__27_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__27_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__27_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__27_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__27_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__27_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__27_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__27_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__27_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__27_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__27_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__27_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__27_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__24_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__24_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__24_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__24_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__24_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__24_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__24_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__24_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__24_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__24_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__24_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__24_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__24_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__24_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__24_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__24_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__15_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__15_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_27_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_27_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_27_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_27_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_27_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_27_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_27_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_27_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_27_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_27_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_27_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_27_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_27_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_27_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_27_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_27_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_27_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_27_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_27_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_27_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_27_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_27_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_27_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_27_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_27_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_27_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_27_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_27_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_27_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_27_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_27_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_27_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_27_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_27_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_27_ccff_tail ) ) ;
grid_clb grid_clb_3__5_ (
    .prog_clk ( { ctsbuf_net_5192501 } ) ,
    .Test_en ( { BUF_net_1200 } ) ,
    .clk ( { ctsbuf_net_101992 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_26_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_169_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__28_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__28_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__28_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__28_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__28_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__28_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__28_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__28_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__28_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__28_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__28_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__28_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__28_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__28_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__28_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__28_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__25_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__25_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__25_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__25_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__25_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__25_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__25_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__25_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__25_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__25_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__25_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__25_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__25_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__25_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__25_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__25_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__16_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__16_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_28_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_28_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_28_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_28_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_28_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_28_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_28_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_28_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_28_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_28_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_28_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_28_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_28_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_28_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_28_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_28_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_28_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_28_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_28_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_28_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_28_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_28_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_28_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_28_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_28_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_28_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_28_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_28_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_28_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_28_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_28_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_28_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_28_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_28_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_28_ccff_tail ) ) ;
grid_clb grid_clb_3__6_ (
    .prog_clk ( { ctsbuf_net_5472529 } ) ,
    .Test_en ( { BUF_net_554 } ) ,
    .clk ( { ctsbuf_net_101992 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_27_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_170_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__29_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__29_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__29_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__29_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__29_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__29_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__29_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__29_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__29_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__29_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__29_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__29_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__29_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__29_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__29_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__29_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__26_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__26_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__26_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__26_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__26_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__26_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__26_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__26_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__26_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__26_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__26_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__26_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__26_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__26_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__26_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__26_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__17_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__17_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_29_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_29_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_29_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_29_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_29_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_29_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_29_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_29_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_29_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_29_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_29_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_29_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_29_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_29_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_29_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_29_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_29_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_29_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_29_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_29_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_29_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_29_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_29_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_29_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_29_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_29_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_29_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_29_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_29_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_29_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_29_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_29_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_29_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_29_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_29_ccff_tail ) ) ;
grid_clb grid_clb_3__7_ (
    .prog_clk ( { ctsbuf_net_5592541 } ) ,
    .Test_en ( { BUF_net_1094 } ) ,
    .clk ( { ctsbuf_net_151997 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_28_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_171_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__30_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__30_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__30_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__30_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__30_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__30_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__30_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__30_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__30_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__30_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__30_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__30_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__30_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__30_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__30_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__30_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__27_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__27_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__27_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__27_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__27_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__27_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__27_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__27_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__27_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__27_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__27_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__27_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__27_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__27_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__27_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__27_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__18_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__18_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_30_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_30_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_30_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_30_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_30_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_30_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_30_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_30_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_30_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_30_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_30_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_30_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_30_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_30_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_30_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_30_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_30_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_30_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_30_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_30_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_30_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_30_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_30_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_30_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_30_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_30_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_30_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_30_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_30_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_30_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_30_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_30_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_30_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_30_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_30_ccff_tail ) ) ;
grid_clb grid_clb_3__8_ (
    .prog_clk ( { ctsbuf_net_5352517 } ) ,
    .Test_en ( { BUF_net_975 } ) ,
    .clk ( { ctsbuf_net_192001 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_29_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_172_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__31_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__31_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__31_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__31_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__31_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__31_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__31_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__31_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__31_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__31_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__31_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__31_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__31_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__31_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__31_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__31_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__28_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__28_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__28_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__28_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__28_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__28_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__28_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__28_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__28_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__28_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__28_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__28_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__28_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__28_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__28_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__28_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__19_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__19_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_31_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_31_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_31_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_31_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_31_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_31_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_31_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_31_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_31_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_31_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_31_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_31_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_31_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_31_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_31_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_31_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_31_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_31_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_31_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_31_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_31_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_31_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_31_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_31_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_31_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_31_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_31_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_31_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_31_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_31_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_31_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_31_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_31_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_31_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_31_ccff_tail ) ) ;
grid_clb grid_clb_3__9_ (
    .prog_clk ( { ctsbuf_net_5052487 } ) ,
    .Test_en ( { BUF_net_1206 } ) ,
    .clk ( { ctsbuf_net_202002 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_30_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_173_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__32_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__32_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__32_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__32_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__32_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__32_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__32_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__32_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__32_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__32_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__32_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__32_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__32_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__32_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__32_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__32_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__29_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__29_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__29_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__29_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__29_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__29_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__29_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__29_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__29_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__29_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__29_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__29_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__29_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__29_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__29_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__29_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__20_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__20_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_32_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_32_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_32_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_32_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_32_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_32_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_32_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_32_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_32_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_32_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_32_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_32_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_32_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_32_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_32_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_32_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_32_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_32_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_32_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_32_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_32_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_32_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_32_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_32_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_32_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_32_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_32_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_32_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_32_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_32_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_32_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_32_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_32_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_32_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_32_ccff_tail ) ) ;
grid_clb grid_clb_3__10_ (
    .prog_clk ( { ctsbuf_net_4682450 } ) ,
    .Test_en ( { BUF_net_979 } ) ,
    .clk ( { ctsbuf_net_232005 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_31_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_174_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__33_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__33_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__33_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__33_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__33_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__33_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__33_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__33_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__33_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__33_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__33_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__33_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__33_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__33_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__33_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__33_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__30_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__30_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__30_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__30_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__30_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__30_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__30_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__30_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__30_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__30_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__30_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__30_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__30_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__30_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__30_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__30_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__21_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__21_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_33_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_33_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_33_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_33_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_33_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_33_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_33_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_33_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_33_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_33_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_33_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_33_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_33_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_33_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_33_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_33_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_33_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_33_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_33_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_33_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_33_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_33_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_33_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_33_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_33_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_33_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_33_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_33_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_33_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_33_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_33_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_33_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_33_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_33_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_33_ccff_tail ) ) ;
grid_clb grid_clb_3__11_ (
    .prog_clk ( { ctsbuf_net_4242406 } ) ,
    .Test_en ( { BUF_net_1209 } ) ,
    .clk ( { ctsbuf_net_252007 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_32_out ) ,
    .top_width_0_height_0__pin_33_ ( { ropt_net_2645 } ) ,
    .right_width_0_height_0__pin_0_ ( cby_1__1__34_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__34_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__34_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__34_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__34_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__34_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__34_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__34_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__34_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__34_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__34_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__34_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__34_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__34_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__34_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__34_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__31_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__31_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__31_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__31_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__31_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__31_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__31_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__31_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__31_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__31_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__31_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__31_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__31_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__31_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__31_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__31_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__22_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__22_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_34_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_34_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_34_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_34_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_34_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_34_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_34_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_34_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_34_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_34_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_34_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_34_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_34_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_34_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_34_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_34_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_34_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_34_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_34_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_34_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_34_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_34_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_34_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_34_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_34_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_34_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_34_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_34_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_34_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_34_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_34_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_34_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_34_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_34_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_34_ccff_tail ) ) ;
grid_clb grid_clb_3__12_ (
    .prog_clk ( { ctsbuf_net_3792361 } ) ,
    .Test_en ( { BUF_net_548 } ) ,
    .clk ( { ctsbuf_net_302012 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_133_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_276_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__35_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__35_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__35_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__35_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__35_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__35_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__35_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__35_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__35_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__35_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__35_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__35_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__35_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__35_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__35_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__35_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__32_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__32_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__32_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__32_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__32_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__32_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__32_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__32_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__32_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__32_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__32_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__32_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__32_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__32_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__32_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__32_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__23_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__23_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_35_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_35_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_35_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_35_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_35_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_35_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_35_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_35_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_35_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_35_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_35_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_35_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_35_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_35_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_35_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_35_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_35_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_35_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_35_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_35_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_35_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_35_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_35_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_35_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_35_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_35_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_35_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_35_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_35_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_35_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_35_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_35_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_35_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_35_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_35_ccff_tail ) ) ;
grid_clb grid_clb_4__1_ (
    .prog_clk ( { ctsbuf_net_3112293 } ) ,
    .Test_en ( { BUF_net_547 } ) ,
    .clk ( { ctsbuf_net_71989 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_33_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_176_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__36_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__36_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__36_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__36_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__36_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__36_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__36_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__36_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__36_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__36_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__36_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__36_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__36_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__36_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__36_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__36_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__0__3_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__0__3_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__0__3_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__0__3_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__0__3_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__0__3_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__0__3_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__0__3_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__0__3_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__0__3_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__0__3_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__0__3_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__0__3_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__0__3_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__0__3_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__0__3_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__24_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__24_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_36_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_36_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_36_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_36_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_36_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_36_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_36_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_36_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_36_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_36_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_36_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_36_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_36_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_36_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_36_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_36_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_36_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_36_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_36_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_36_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_36_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_36_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_36_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_36_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_36_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_36_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_36_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_36_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_36_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_36_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_36_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_36_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_36_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_36_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_36_ccff_tail ) ) ;
grid_clb grid_clb_4__2_ (
    .prog_clk ( { ctsbuf_net_3562338 } ) ,
    .Test_en ( { BUF_net_1444 } ) ,
    .clk ( { ctsbuf_net_71989 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_34_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_177_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__37_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__37_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__37_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__37_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__37_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__37_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__37_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__37_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__37_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__37_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__37_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__37_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__37_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__37_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__37_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__37_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__33_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__33_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__33_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__33_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__33_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__33_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__33_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__33_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__33_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__33_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__33_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__33_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__33_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__33_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__33_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__33_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__25_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__25_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_37_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_37_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_37_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_37_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_37_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_37_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_37_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_37_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_37_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_37_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_37_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_37_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_37_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_37_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_37_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_37_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_37_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_37_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_37_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_37_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_37_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_37_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_37_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_37_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_37_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_37_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_37_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_37_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_37_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_37_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_37_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_37_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_37_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_37_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_37_ccff_tail ) ) ;
grid_clb grid_clb_4__3_ (
    .prog_clk ( { ctsbuf_net_4002382 } ) ,
    .Test_en ( { BUF_net_1288 } ) ,
    .clk ( { ctsbuf_net_81990 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_35_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_178_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__38_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__38_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__38_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__38_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__38_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__38_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__38_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__38_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__38_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__38_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__38_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__38_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__38_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__38_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__38_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__38_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__34_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__34_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__34_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__34_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__34_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__34_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__34_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__34_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__34_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__34_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__34_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__34_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__34_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__34_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__34_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__34_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__26_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__26_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_38_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_38_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_38_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_38_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_38_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_38_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_38_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_38_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_38_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_38_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_38_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_38_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_38_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_38_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_38_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_38_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_38_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_38_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_38_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_38_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_38_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_38_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_38_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_38_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_38_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_38_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_38_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_38_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_38_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_38_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_38_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_38_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_38_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_38_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_38_ccff_tail ) ) ;
grid_clb grid_clb_4__4_ (
    .prog_clk ( { ctsbuf_net_4452427 } ) ,
    .Test_en ( { BUF_net_1188 } ) ,
    .clk ( { ctsbuf_net_121994 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_36_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_179_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__39_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__39_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__39_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__39_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__39_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__39_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__39_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__39_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__39_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__39_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__39_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__39_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__39_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__39_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__39_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__39_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__35_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__35_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__35_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__35_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__35_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__35_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__35_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__35_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__35_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__35_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__35_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__35_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__35_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__35_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__35_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__35_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__27_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__27_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_39_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_39_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_39_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_39_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_39_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_39_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_39_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_39_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_39_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_39_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_39_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_39_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_39_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_39_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_39_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_39_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_39_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_39_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_39_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_39_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_39_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_39_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_39_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_39_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_39_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_39_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_39_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_39_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_39_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_39_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_39_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_39_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_39_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_39_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_39_ccff_tail ) ) ;
grid_clb grid_clb_4__5_ (
    .prog_clk ( { ctsbuf_net_4872469 } ) ,
    .Test_en ( { BUF_net_1448 } ) ,
    .clk ( { ctsbuf_net_121994 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_37_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_180_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__40_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__40_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__40_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__40_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__40_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__40_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__40_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__40_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__40_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__40_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__40_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__40_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__40_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__40_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__40_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__40_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__36_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__36_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__36_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__36_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__36_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__36_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__36_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__36_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__36_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__36_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__36_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__36_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__36_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__36_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__36_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__36_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__28_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__28_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_40_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_40_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_40_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_40_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_40_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_40_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_40_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_40_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_40_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_40_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_40_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_40_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_40_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_40_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_40_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_40_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_40_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_40_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_40_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_40_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_40_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_40_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_40_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_40_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_40_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_40_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_40_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_40_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_40_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_40_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_40_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_40_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_40_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_40_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_40_ccff_tail ) ) ;
grid_clb grid_clb_4__6_ (
    .prog_clk ( { ctsbuf_net_5202502 } ) ,
    .Test_en ( { BUF_net_542 } ) ,
    .clk ( { ctsbuf_net_182000 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_38_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_181_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__41_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__41_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__41_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__41_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__41_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__41_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__41_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__41_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__41_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__41_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__41_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__41_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__41_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__41_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__41_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__41_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__37_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__37_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__37_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__37_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__37_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__37_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__37_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__37_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__37_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__37_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__37_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__37_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__37_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__37_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__37_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__37_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__29_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__29_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_41_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_41_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_41_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_41_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_41_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_41_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_41_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_41_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_41_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_41_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_41_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_41_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_41_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_41_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_41_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_41_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_41_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_41_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_41_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_41_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_41_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_41_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_41_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_41_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_41_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_41_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_41_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_41_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_41_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_41_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_41_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_41_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_41_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_41_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_41_ccff_tail ) ) ;
grid_clb grid_clb_4__7_ (
    .prog_clk ( { ctsbuf_net_5372519 } ) ,
    .Test_en ( { BUF_net_541 } ) ,
    .clk ( { ctsbuf_net_192001 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_39_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_182_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__42_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__42_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__42_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__42_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__42_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__42_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__42_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__42_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__42_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__42_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__42_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__42_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__42_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__42_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__42_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__42_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__38_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__38_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__38_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__38_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__38_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__38_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__38_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__38_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__38_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__38_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__38_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__38_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__38_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__38_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__38_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__38_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__30_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__30_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_42_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_42_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_42_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_42_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_42_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_42_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_42_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_42_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_42_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_42_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_42_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_42_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_42_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_42_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_42_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_42_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_42_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_42_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_42_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_42_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_42_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_42_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_42_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_42_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_42_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_42_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_42_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_42_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_42_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_42_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_42_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_42_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_42_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_42_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_42_ccff_tail ) ) ;
grid_clb grid_clb_4__8_ (
    .prog_clk ( { ctsbuf_net_5072489 } ) ,
    .Test_en ( { BUF_net_1450 } ) ,
    .clk ( { ctsbuf_net_192001 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_40_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_183_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__43_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__43_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__43_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__43_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__43_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__43_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__43_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__43_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__43_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__43_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__43_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__43_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__43_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__43_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__43_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__43_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__39_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__39_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__39_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__39_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__39_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__39_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__39_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__39_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__39_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__39_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__39_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__39_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__39_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__39_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__39_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__39_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__31_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__31_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_43_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_43_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_43_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_43_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_43_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_43_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_43_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_43_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_43_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_43_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_43_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_43_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_43_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_43_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_43_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_43_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_43_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_43_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_43_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_43_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_43_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_43_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_43_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_43_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_43_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_43_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_43_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_43_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_43_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_43_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_43_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_43_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_43_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_43_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_43_ccff_tail ) ) ;
grid_clb grid_clb_4__9_ (
    .prog_clk ( { ctsbuf_net_4692451 } ) ,
    .Test_en ( { BUF_net_1451 } ) ,
    .clk ( { ctsbuf_net_232005 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_41_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_184_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__44_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__44_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__44_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__44_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__44_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__44_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__44_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__44_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__44_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__44_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__44_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__44_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__44_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__44_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__44_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__44_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__40_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__40_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__40_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__40_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__40_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__40_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__40_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__40_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__40_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__40_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__40_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__40_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__40_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__40_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__40_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__40_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__32_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__32_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_44_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_44_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_44_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_44_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_44_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_44_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_44_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_44_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_44_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_44_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_44_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_44_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_44_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_44_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_44_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_44_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_44_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_44_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_44_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_44_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_44_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_44_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_44_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_44_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_44_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_44_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_44_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_44_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_44_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_44_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_44_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_44_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_44_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_44_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_44_ccff_tail ) ) ;
grid_clb grid_clb_4__10_ (
    .prog_clk ( { ctsbuf_net_4262408 } ) ,
    .Test_en ( { BUF_net_1194 } ) ,
    .clk ( { ctsbuf_net_232005 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_42_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_185_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__45_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__45_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__45_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__45_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__45_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__45_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__45_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__45_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__45_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__45_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__45_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__45_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__45_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__45_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__45_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__45_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__41_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__41_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__41_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__41_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__41_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__41_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__41_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__41_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__41_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__41_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__41_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__41_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__41_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__41_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__41_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__41_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__33_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__33_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_45_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_45_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_45_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_45_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_45_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_45_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_45_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_45_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_45_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_45_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_45_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_45_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_45_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_45_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_45_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_45_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_45_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_45_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_45_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_45_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_45_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_45_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_45_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_45_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_45_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_45_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_45_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_45_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_45_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_45_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_45_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_45_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_45_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_45_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_45_ccff_tail ) ) ;
grid_clb grid_clb_4__11_ (
    .prog_clk ( { ctsbuf_net_3802362 } ) ,
    .Test_en ( { BUF_net_1549 } ) ,
    .clk ( { ctsbuf_net_282010 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_43_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_186_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__46_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__46_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__46_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__46_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__46_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__46_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__46_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__46_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__46_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__46_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__46_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__46_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__46_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__46_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__46_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__46_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__42_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__42_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__42_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__42_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__42_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__42_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__42_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__42_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__42_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__42_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__42_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__42_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__42_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__42_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__42_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__42_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__34_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__34_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_46_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_46_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_46_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_46_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_46_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_46_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_46_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_46_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_46_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_46_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_46_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_46_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_46_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_46_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_46_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_46_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_46_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_46_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_46_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_46_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_46_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_46_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_46_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_46_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_46_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_46_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_46_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_46_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_46_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_46_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_46_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_46_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_46_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_46_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_46_ccff_tail ) ) ;
grid_clb grid_clb_4__12_ (
    .prog_clk ( { ctsbuf_net_3362318 } ) ,
    .Test_en ( { BUF_net_536 } ) ,
    .clk ( { ctsbuf_net_302012 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_134_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_277_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__47_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__47_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__47_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__47_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__47_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__47_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__47_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__47_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__47_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__47_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__47_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__47_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__47_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__47_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__47_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__47_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__43_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__43_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__43_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__43_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__43_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__43_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__43_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__43_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__43_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__43_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__43_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__43_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__43_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__43_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__43_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__43_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__35_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__35_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_47_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_47_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_47_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_47_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_47_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_47_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_47_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_47_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_47_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_47_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_47_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_47_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_47_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_47_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_47_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_47_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_47_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_47_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_47_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_47_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_47_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_47_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_47_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_47_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_47_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_47_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_47_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_47_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_47_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_47_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_47_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_47_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_47_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_47_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_47_ccff_tail ) ) ;
grid_clb grid_clb_5__1_ (
    .prog_clk ( { ctsbuf_net_2662248 } ) ,
    .Test_en ( { BUF_net_535 } ) ,
    .clk ( { ctsbuf_net_71989 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_44_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_187_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__48_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__48_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__48_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__48_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__48_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__48_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__48_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__48_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__48_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__48_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__48_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__48_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__48_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__48_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__48_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__48_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__0__4_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__0__4_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__0__4_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__0__4_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__0__4_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__0__4_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__0__4_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__0__4_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__0__4_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__0__4_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__0__4_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__0__4_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__0__4_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__0__4_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__0__4_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__0__4_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__36_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__36_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_48_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_48_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_48_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_48_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_48_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_48_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_48_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_48_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_48_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_48_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_48_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_48_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_48_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_48_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_48_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_48_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_48_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_48_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_48_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_48_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_48_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_48_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_48_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_48_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_48_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_48_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_48_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_48_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_48_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_48_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_48_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_48_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_48_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_48_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_48_ccff_tail ) ) ;
grid_clb grid_clb_5__2_ (
    .prog_clk ( { ctsbuf_net_3122294 } ) ,
    .Test_en ( { BUF_net_1615 } ) ,
    .clk ( { ctsbuf_net_81990 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_45_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_188_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__49_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__49_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__49_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__49_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__49_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__49_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__49_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__49_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__49_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__49_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__49_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__49_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__49_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__49_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__49_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__49_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__44_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__44_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__44_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__44_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__44_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__44_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__44_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__44_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__44_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__44_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__44_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__44_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__44_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__44_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__44_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__44_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__37_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__37_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_49_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_49_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_49_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_49_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_49_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_49_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_49_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_49_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_49_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_49_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_49_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_49_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_49_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_49_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_49_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_49_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_49_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_49_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_49_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_49_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_49_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_49_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_49_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_49_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_49_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_49_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_49_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_49_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_49_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_49_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_49_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_49_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_49_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_49_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_49_ccff_tail ) ) ;
grid_clb grid_clb_5__3_ (
    .prog_clk ( { ctsbuf_net_3572339 } ) ,
    .Test_en ( { BUF_net_1446 } ) ,
    .clk ( { ctsbuf_net_81990 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_46_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_189_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__50_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__50_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__50_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__50_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__50_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__50_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__50_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__50_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__50_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__50_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__50_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__50_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__50_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__50_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__50_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__50_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__45_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__45_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__45_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__45_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__45_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__45_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__45_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__45_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__45_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__45_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__45_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__45_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__45_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__45_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__45_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__45_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__38_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__38_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_50_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_50_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_50_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_50_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_50_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_50_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_50_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_50_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_50_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_50_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_50_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_50_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_50_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_50_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_50_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_50_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_50_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_50_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_50_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_50_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_50_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_50_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_50_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_50_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_50_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_50_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_50_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_50_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_50_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_50_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_50_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_50_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_50_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_50_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_50_ccff_tail ) ) ;
grid_clb grid_clb_5__4_ (
    .prog_clk ( { ctsbuf_net_4012383 } ) ,
    .Test_en ( { BUF_net_1375 } ) ,
    .clk ( { ctsbuf_net_121994 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_47_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_190_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__51_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__51_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__51_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__51_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__51_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__51_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__51_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__51_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__51_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__51_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__51_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__51_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__51_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__51_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__51_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__51_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__46_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__46_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__46_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__46_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__46_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__46_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__46_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__46_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__46_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__46_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__46_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__46_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__46_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__46_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__46_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__46_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__39_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__39_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_51_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_51_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_51_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_51_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_51_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_51_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_51_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_51_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_51_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_51_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_51_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_51_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_51_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_51_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_51_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_51_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_51_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_51_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_51_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_51_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_51_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_51_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_51_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_51_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_51_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_51_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_51_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_51_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_51_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_51_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_51_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_51_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_51_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_51_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_51_ccff_tail ) ) ;
grid_clb grid_clb_5__5_ (
    .prog_clk ( { ctsbuf_net_4462428 } ) ,
    .Test_en ( { BUF_net_1627 } ) ,
    .clk ( { ctsbuf_net_182000 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_48_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_191_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__52_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__52_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__52_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__52_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__52_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__52_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__52_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__52_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__52_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__52_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__52_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__52_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__52_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__52_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__52_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__52_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__47_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__47_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__47_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__47_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__47_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__47_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__47_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__47_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__47_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__47_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__47_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__47_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__47_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__47_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__47_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__47_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__40_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__40_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_52_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_52_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_52_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_52_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_52_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_52_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_52_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_52_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_52_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_52_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_52_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_52_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_52_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_52_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_52_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_52_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_52_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_52_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_52_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_52_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_52_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_52_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_52_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_52_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_52_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_52_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_52_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_52_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_52_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_52_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_52_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_52_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_52_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_52_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_52_ccff_tail ) ) ;
grid_clb grid_clb_5__6_ (
    .prog_clk ( { ctsbuf_net_4882470 } ) ,
    .Test_en ( { BUF_net_530 } ) ,
    .clk ( { ctsbuf_net_182000 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_49_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_192_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__53_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__53_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__53_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__53_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__53_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__53_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__53_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__53_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__53_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__53_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__53_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__53_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__53_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__53_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__53_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__53_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__48_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__48_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__48_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__48_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__48_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__48_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__48_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__48_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__48_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__48_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__48_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__48_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__48_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__48_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__48_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__48_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__41_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__41_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_53_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_53_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_53_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_53_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_53_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_53_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_53_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_53_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_53_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_53_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_53_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_53_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_53_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_53_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_53_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_53_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_53_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_53_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_53_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_53_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_53_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_53_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_53_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_53_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_53_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_53_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_53_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_53_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_53_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_53_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_53_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_53_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_53_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_53_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_53_ccff_tail ) ) ;
grid_clb grid_clb_5__7_ (
    .prog_clk ( { ctsbuf_net_5082490 } ) ,
    .Test_en ( { BUF_net_1109 } ) ,
    .clk ( { ctsbuf_net_192001 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_50_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_193_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__54_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__54_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__54_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__54_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__54_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__54_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__54_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__54_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__54_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__54_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__54_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__54_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__54_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__54_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__54_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__54_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__49_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__49_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__49_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__49_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__49_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__49_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__49_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__49_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__49_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__49_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__49_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__49_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__49_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__49_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__49_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__49_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__42_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__42_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_54_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_54_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_54_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_54_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_54_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_54_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_54_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_54_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_54_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_54_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_54_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_54_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_54_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_54_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_54_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_54_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_54_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_54_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_54_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_54_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_54_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_54_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_54_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_54_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_54_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_54_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_54_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_54_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_54_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_54_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_54_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_54_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_54_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_54_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_54_ccff_tail ) ) ;
grid_clb grid_clb_5__8_ (
    .prog_clk ( { ctsbuf_net_4712453 } ) ,
    .Test_en ( { BUF_net_1576 } ) ,
    .clk ( { ctsbuf_net_192001 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_51_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_194_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__55_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__55_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__55_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__55_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__55_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__55_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__55_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__55_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__55_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__55_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__55_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__55_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__55_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__55_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__55_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__55_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__50_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__50_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__50_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__50_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__50_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__50_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__50_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__50_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__50_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__50_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__50_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__50_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__50_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__50_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__50_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__50_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__43_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__43_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_55_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_55_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_55_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_55_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_55_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_55_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_55_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_55_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_55_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_55_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_55_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_55_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_55_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_55_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_55_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_55_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_55_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_55_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_55_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_55_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_55_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_55_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_55_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_55_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_55_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_55_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_55_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_55_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_55_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_55_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_55_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_55_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_55_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_55_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_55_ccff_tail ) ) ;
grid_clb grid_clb_5__9_ (
    .prog_clk ( { ctsbuf_net_4272409 } ) ,
    .Test_en ( { BUF_net_1626 } ) ,
    .clk ( { ctsbuf_net_232005 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_52_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_195_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__56_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__56_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__56_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__56_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__56_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__56_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__56_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__56_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__56_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__56_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__56_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__56_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__56_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__56_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__56_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__56_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__51_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__51_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__51_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__51_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__51_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__51_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__51_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__51_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__51_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__51_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__51_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__51_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__51_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__51_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__51_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__51_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__44_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__44_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_56_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_56_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_56_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_56_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_56_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_56_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_56_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_56_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_56_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_56_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_56_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_56_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_56_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_56_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_56_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_56_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_56_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_56_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_56_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_56_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_56_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_56_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_56_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_56_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_56_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_56_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_56_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_56_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_56_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_56_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_56_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_56_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_56_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_56_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_56_ccff_tail ) ) ;
grid_clb grid_clb_5__10_ (
    .prog_clk ( { ctsbuf_net_3822364 } ) ,
    .Test_en ( { BUF_net_1376 } ) ,
    .clk ( { ctsbuf_net_232005 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_53_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_196_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__57_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__57_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__57_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__57_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__57_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__57_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__57_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__57_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__57_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__57_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__57_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__57_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__57_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__57_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__57_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__57_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__52_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__52_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__52_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__52_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__52_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__52_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__52_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__52_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__52_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__52_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__52_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__52_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__52_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__52_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__52_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__52_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__45_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__45_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_57_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_57_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_57_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_57_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_57_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_57_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_57_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_57_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_57_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_57_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_57_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_57_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_57_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_57_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_57_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_57_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_57_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_57_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_57_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_57_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_57_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_57_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_57_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_57_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_57_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_57_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_57_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_57_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_57_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_57_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_57_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_57_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_57_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_57_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_57_ccff_tail ) ) ;
grid_clb grid_clb_5__11_ (
    .prog_clk ( { ctsbuf_net_3372319 } ) ,
    .Test_en ( { BUF_net_1679 } ) ,
    .clk ( { ctsbuf_net_282010 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_54_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_197_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__58_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__58_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__58_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__58_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__58_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__58_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__58_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__58_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__58_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__58_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__58_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__58_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__58_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__58_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__58_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__58_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__53_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__53_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__53_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__53_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__53_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__53_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__53_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__53_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__53_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__53_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__53_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__53_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__53_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__53_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__53_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__53_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__46_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__46_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_58_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_58_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_58_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_58_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_58_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_58_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_58_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_58_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_58_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_58_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_58_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_58_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_58_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_58_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_58_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_58_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_58_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_58_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_58_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_58_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_58_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_58_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_58_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_58_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_58_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_58_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_58_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_58_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_58_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_58_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_58_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_58_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_58_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_58_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_58_ccff_tail ) ) ;
grid_clb grid_clb_5__12_ (
    .prog_clk ( { ctsbuf_net_2902272 } ) ,
    .Test_en ( Test_en ) ,
    .clk ( { ctsbuf_net_302012 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_135_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_278_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__59_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__59_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__59_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__59_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__59_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__59_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__59_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__59_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__59_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__59_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__59_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__59_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__59_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__59_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__59_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__59_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__54_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__54_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__54_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__54_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__54_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__54_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__54_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__54_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__54_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__54_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__54_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__54_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__54_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__54_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__54_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__54_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__47_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__47_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_59_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_59_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_59_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_59_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_59_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_59_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_59_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_59_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_59_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_59_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_59_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_59_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_59_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_59_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_59_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_59_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_59_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_59_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_59_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_59_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_59_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_59_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_59_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_59_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_59_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_59_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_59_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_59_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_59_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_59_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_59_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_59_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_59_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_59_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_59_ccff_tail ) ) ;
grid_clb grid_clb_6__1_ (
    .prog_clk ( { ctsbuf_net_2212203 } ) ,
    .Test_en ( { BUF_net_523 } ) ,
    .clk ( { ctsbuf_net_71989 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_55_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_198_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__60_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__60_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__60_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__60_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__60_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__60_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__60_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__60_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__60_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__60_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__60_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__60_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__60_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__60_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__60_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__60_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__0__5_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__0__5_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__0__5_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__0__5_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__0__5_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__0__5_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__0__5_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__0__5_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__0__5_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__0__5_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__0__5_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__0__5_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__0__5_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__0__5_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__0__5_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__0__5_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__48_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__48_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_60_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_60_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_60_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_60_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_60_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_60_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_60_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_60_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_60_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_60_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_60_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_60_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_60_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_60_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_60_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_60_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_60_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_60_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_60_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_60_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_60_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_60_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_60_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_60_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_60_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_60_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_60_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_60_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_60_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_60_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_60_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_60_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_60_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_60_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_60_ccff_tail ) ) ;
grid_clb grid_clb_6__2_ (
    .prog_clk ( { ctsbuf_net_2672249 } ) ,
    .Test_en ( { BUF_net_1715 } ) ,
    .clk ( { ctsbuf_net_131995 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_56_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_199_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__61_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__61_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__61_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__61_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__61_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__61_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__61_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__61_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__61_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__61_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__61_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__61_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__61_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__61_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__61_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__61_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__55_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__55_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__55_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__55_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__55_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__55_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__55_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__55_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__55_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__55_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__55_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__55_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__55_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__55_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__55_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__55_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__49_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__49_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_61_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_61_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_61_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_61_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_61_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_61_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_61_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_61_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_61_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_61_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_61_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_61_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_61_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_61_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_61_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_61_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_61_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_61_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_61_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_61_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_61_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_61_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_61_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_61_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_61_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_61_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_61_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_61_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_61_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_61_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_61_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_61_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_61_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_61_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_61_ccff_tail ) ) ;
grid_clb grid_clb_6__3_ (
    .prog_clk ( { ctsbuf_net_3132295 } ) ,
    .Test_en ( { BUF_net_1569 } ) ,
    .clk ( { ctsbuf_net_131995 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_57_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_200_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__62_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__62_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__62_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__62_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__62_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__62_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__62_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__62_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__62_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__62_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__62_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__62_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__62_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__62_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__62_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__62_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__56_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__56_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__56_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__56_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__56_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__56_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__56_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__56_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__56_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__56_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__56_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__56_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__56_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__56_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__56_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__56_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__50_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__50_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_62_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_62_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_62_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_62_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_62_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_62_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_62_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_62_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_62_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_62_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_62_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_62_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_62_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_62_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_62_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_62_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_62_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_62_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_62_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_62_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_62_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_62_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_62_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_62_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_62_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_62_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_62_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_62_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_62_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_62_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_62_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_62_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_62_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_62_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_62_ccff_tail ) ) ;
grid_clb grid_clb_6__4_ (
    .prog_clk ( { ctsbuf_net_3582340 } ) ,
    .Test_en ( { BUF_net_1571 } ) ,
    .clk ( { ctsbuf_net_131995 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_58_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_201_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__63_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__63_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__63_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__63_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__63_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__63_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__63_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__63_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__63_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__63_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__63_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__63_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__63_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__63_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__63_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__63_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__57_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__57_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__57_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__57_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__57_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__57_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__57_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__57_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__57_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__57_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__57_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__57_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__57_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__57_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__57_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__57_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__51_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__51_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_63_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_63_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_63_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_63_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_63_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_63_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_63_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_63_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_63_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_63_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_63_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_63_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_63_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_63_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_63_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_63_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_63_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_63_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_63_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_63_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_63_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_63_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_63_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_63_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_63_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_63_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_63_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_63_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_63_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_63_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_63_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_63_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_63_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_63_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_63_ccff_tail ) ) ;
grid_clb grid_clb_6__5_ (
    .prog_clk ( { ctsbuf_net_4022384 } ) ,
    .Test_en ( { BUF_net_519 } ) ,
    .clk ( { ctsbuf_net_182000 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_59_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_202_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__64_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__64_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__64_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__64_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__64_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__64_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__64_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__64_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__64_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__64_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__64_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__64_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__64_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__64_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__64_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__64_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__58_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__58_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__58_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__58_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__58_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__58_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__58_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__58_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__58_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__58_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__58_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__58_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__58_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__58_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__58_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__58_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__52_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__52_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_64_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_64_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_64_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_64_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_64_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_64_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_64_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_64_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_64_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_64_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_64_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_64_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_64_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_64_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_64_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_64_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_64_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_64_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_64_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_64_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_64_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_64_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_64_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_64_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_64_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_64_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_64_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_64_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_64_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_64_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_64_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_64_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_64_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_64_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_64_ccff_tail ) ) ;
grid_clb grid_clb_6__6_ (
    .prog_clk ( { ctsbuf_net_4472429 } ) ,
    .Test_en ( { BUF_net_518 } ) ,
    .clk ( { ctsbuf_net_182000 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_60_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_203_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__65_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__65_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__65_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__65_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__65_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__65_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__65_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__65_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__65_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__65_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__65_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__65_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__65_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__65_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__65_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__65_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__59_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__59_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__59_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__59_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__59_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__59_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__59_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__59_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__59_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__59_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__59_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__59_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__59_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__59_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__59_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__59_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__53_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__53_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_65_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_65_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_65_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_65_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_65_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_65_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_65_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_65_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_65_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_65_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_65_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_65_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_65_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_65_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_65_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_65_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_65_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_65_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_65_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_65_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_65_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_65_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_65_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_65_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_65_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_65_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_65_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_65_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_65_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_65_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_65_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_65_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_65_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_65_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_65_ccff_tail ) ) ;
grid_clb grid_clb_6__7_ (
    .prog_clk ( { ctsbuf_net_4732455 } ) ,
    .Test_en ( { BUF_net_517 } ) ,
    .clk ( { ctsbuf_net_192001 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_61_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_204_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__66_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__66_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__66_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__66_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__66_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__66_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__66_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__66_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__66_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__66_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__66_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__66_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__66_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__66_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__66_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__66_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__60_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__60_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__60_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__60_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__60_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__60_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__60_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__60_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__60_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__60_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__60_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__60_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__60_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__60_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__60_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__60_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__54_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__54_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_66_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_66_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_66_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_66_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_66_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_66_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_66_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_66_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_66_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_66_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_66_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_66_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_66_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_66_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_66_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_66_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_66_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_66_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_66_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_66_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_66_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_66_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_66_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_66_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_66_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_66_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_66_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_66_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_66_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_66_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_66_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_66_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_66_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_66_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_66_ccff_tail ) ) ;
grid_clb grid_clb_6__8_ (
    .prog_clk ( { ctsbuf_net_4292411 } ) ,
    .Test_en ( { BUF_net_1764 } ) ,
    .clk ( { ctsbuf_net_262008 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_62_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_205_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__67_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__67_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__67_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__67_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__67_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__67_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__67_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__67_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__67_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__67_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__67_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__67_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__67_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__67_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__67_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__67_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__61_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__61_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__61_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__61_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__61_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__61_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__61_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__61_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__61_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__61_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__61_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__61_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__61_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__61_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__61_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__61_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__55_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__55_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_67_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_67_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_67_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_67_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_67_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_67_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_67_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_67_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_67_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_67_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_67_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_67_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_67_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_67_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_67_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_67_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_67_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_67_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_67_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_67_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_67_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_67_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_67_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_67_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_67_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_67_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_67_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_67_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_67_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_67_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_67_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_67_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_67_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_67_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_67_ccff_tail ) ) ;
grid_clb grid_clb_6__9_ (
    .prog_clk ( { ctsbuf_net_3832365 } ) ,
    .Test_en ( { BUF_net_1724 } ) ,
    .clk ( { ctsbuf_net_262008 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_63_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_206_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__68_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__68_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__68_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__68_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__68_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__68_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__68_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__68_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__68_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__68_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__68_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__68_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__68_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__68_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__68_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__68_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__62_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__62_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__62_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__62_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__62_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__62_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__62_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__62_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__62_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__62_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__62_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__62_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__62_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__62_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__62_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__62_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__56_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__56_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_68_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_68_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_68_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_68_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_68_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_68_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_68_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_68_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_68_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_68_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_68_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_68_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_68_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_68_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_68_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_68_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_68_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_68_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_68_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_68_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_68_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_68_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_68_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_68_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_68_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_68_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_68_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_68_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_68_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_68_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_68_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_68_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_68_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_68_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_68_ccff_tail ) ) ;
grid_clb grid_clb_6__10_ (
    .prog_clk ( { ctsbuf_net_3392321 } ) ,
    .Test_en ( { BUF_net_1522 } ) ,
    .clk ( { ctsbuf_net_282010 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_64_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_207_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__69_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__69_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__69_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__69_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__69_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__69_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__69_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__69_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__69_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__69_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__69_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__69_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__69_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__69_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__69_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__69_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__63_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__63_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__63_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__63_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__63_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__63_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__63_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__63_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__63_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__63_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__63_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__63_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__63_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__63_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__63_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__63_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__57_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__57_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_69_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_69_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_69_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_69_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_69_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_69_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_69_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_69_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_69_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_69_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_69_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_69_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_69_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_69_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_69_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_69_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_69_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_69_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_69_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_69_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_69_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_69_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_69_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_69_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_69_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_69_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_69_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_69_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_69_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_69_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_69_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_69_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_69_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_69_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_69_ccff_tail ) ) ;
grid_clb grid_clb_6__11_ (
    .prog_clk ( { ctsbuf_net_2912273 } ) ,
    .Test_en ( { BUF_net_1725 } ) ,
    .clk ( { ctsbuf_net_282010 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_65_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_208_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__70_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__70_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__70_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__70_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__70_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__70_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__70_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__70_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__70_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__70_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__70_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__70_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__70_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__70_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__70_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__70_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__64_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__64_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__64_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__64_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__64_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__64_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__64_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__64_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__64_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__64_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__64_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__64_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__64_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__64_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__64_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__64_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__58_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__58_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_70_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_70_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_70_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_70_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_70_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_70_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_70_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_70_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_70_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_70_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_70_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_70_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_70_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_70_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_70_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_70_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_70_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_70_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_70_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_70_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_70_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_70_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_70_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_70_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_70_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_70_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_70_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_70_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_70_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_70_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_70_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_70_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_70_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_70_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_70_ccff_tail ) ) ;
grid_clb grid_clb_6__12_ (
    .prog_clk ( { ctsbuf_net_2462228 } ) ,
    .Test_en ( Test_en ) ,
    .clk ( { ctsbuf_net_302012 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_136_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_279_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__71_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__71_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__71_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__71_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__71_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__71_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__71_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__71_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__71_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__71_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__71_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__71_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__71_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__71_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__71_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__71_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__65_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__65_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__65_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__65_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__65_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__65_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__65_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__65_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__65_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__65_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__65_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__65_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__65_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__65_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__65_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__65_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__59_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__59_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_71_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_71_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_71_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_71_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_71_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_71_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_71_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_71_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_71_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_71_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_71_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_71_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_71_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_71_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_71_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_71_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_71_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_71_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_71_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_71_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_71_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_71_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_71_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_71_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_71_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_71_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_71_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_71_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_71_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_71_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_71_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_71_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_71_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_71_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_71_ccff_tail ) ) ;
grid_clb grid_clb_7__1_ (
    .prog_clk ( { ctsbuf_net_1772159 } ) ,
    .Test_en ( { BUF_net_511 } ) ,
    .clk ( { ctsbuf_net_61988 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_66_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_209_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__72_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__72_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__72_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__72_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__72_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__72_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__72_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__72_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__72_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__72_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__72_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__72_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__72_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__72_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__72_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__72_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__0__6_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__0__6_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__0__6_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__0__6_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__0__6_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__0__6_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__0__6_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__0__6_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__0__6_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__0__6_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__0__6_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__0__6_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__0__6_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__0__6_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__0__6_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__0__6_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__60_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__60_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_72_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_72_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_72_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_72_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_72_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_72_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_72_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_72_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_72_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_72_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_72_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_72_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_72_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_72_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_72_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_72_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_72_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_72_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_72_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_72_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_72_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_72_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_72_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_72_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_72_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_72_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_72_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_72_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_72_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_72_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_72_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_72_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_72_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_72_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_72_ccff_tail ) ) ;
grid_clb grid_clb_7__2_ (
    .prog_clk ( { ctsbuf_net_2222204 } ) ,
    .Test_en ( { BUF_net_1727 } ) ,
    .clk ( { ctsbuf_net_131995 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_67_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_210_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__73_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__73_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__73_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__73_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__73_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__73_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__73_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__73_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__73_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__73_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__73_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__73_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__73_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__73_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__73_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__73_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__66_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__66_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__66_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__66_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__66_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__66_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__66_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__66_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__66_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__66_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__66_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__66_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__66_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__66_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__66_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__66_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__61_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__61_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_73_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_73_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_73_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_73_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_73_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_73_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_73_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_73_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_73_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_73_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_73_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_73_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_73_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_73_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_73_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_73_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_73_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_73_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_73_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_73_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_73_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_73_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_73_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_73_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_73_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_73_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_73_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_73_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_73_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_73_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_73_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_73_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_73_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_73_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_73_ccff_tail ) ) ;
grid_clb grid_clb_7__3_ (
    .prog_clk ( { ctsbuf_net_2682250 } ) ,
    .Test_en ( { BUF_net_1514 } ) ,
    .clk ( { ctsbuf_net_111993 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_68_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_211_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__74_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__74_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__74_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__74_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__74_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__74_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__74_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__74_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__74_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__74_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__74_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__74_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__74_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__74_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__74_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__74_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__67_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__67_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__67_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__67_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__67_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__67_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__67_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__67_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__67_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__67_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__67_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__67_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__67_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__67_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__67_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__67_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__62_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__62_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_74_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_74_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_74_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_74_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_74_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_74_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_74_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_74_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_74_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_74_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_74_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_74_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_74_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_74_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_74_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_74_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_74_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_74_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_74_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_74_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_74_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_74_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_74_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_74_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_74_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_74_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_74_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_74_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_74_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_74_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_74_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_74_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_74_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_74_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_74_ccff_tail ) ) ;
grid_clb grid_clb_7__4_ (
    .prog_clk ( { ctsbuf_net_3142296 } ) ,
    .Test_en ( { BUF_net_1657 } ) ,
    .clk ( { ctsbuf_net_131995 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_69_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_212_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__75_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__75_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__75_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__75_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__75_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__75_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__75_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__75_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__75_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__75_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__75_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__75_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__75_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__75_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__75_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__75_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__68_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__68_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__68_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__68_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__68_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__68_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__68_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__68_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__68_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__68_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__68_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__68_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__68_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__68_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__68_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__68_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__63_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__63_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_75_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_75_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_75_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_75_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_75_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_75_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_75_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_75_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_75_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_75_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_75_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_75_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_75_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_75_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_75_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_75_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_75_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_75_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_75_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_75_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_75_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_75_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_75_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_75_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_75_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_75_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_75_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_75_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_75_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_75_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_75_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_75_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_75_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_75_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_75_ccff_tail ) ) ;
grid_clb grid_clb_7__5_ (
    .prog_clk ( { ctsbuf_net_3592341 } ) ,
    .Test_en ( { BUF_net_1741 } ) ,
    .clk ( { ctsbuf_net_161998 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_70_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_213_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__76_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__76_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__76_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__76_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__76_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__76_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__76_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__76_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__76_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__76_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__76_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__76_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__76_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__76_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__76_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__76_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__69_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__69_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__69_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__69_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__69_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__69_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__69_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__69_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__69_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__69_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__69_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__69_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__69_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__69_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__69_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__69_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__64_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__64_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_76_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_76_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_76_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_76_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_76_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_76_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_76_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_76_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_76_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_76_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_76_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_76_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_76_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_76_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_76_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_76_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_76_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_76_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_76_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_76_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_76_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_76_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_76_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_76_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_76_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_76_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_76_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_76_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_76_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_76_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_76_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_76_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_76_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_76_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_76_ccff_tail ) ) ;
grid_clb grid_clb_7__6_ (
    .prog_clk ( { ctsbuf_net_4032385 } ) ,
    .Test_en ( { BUF_net_506 } ) ,
    .clk ( { ctsbuf_net_182000 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_71_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_214_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__77_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__77_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__77_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__77_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__77_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__77_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__77_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__77_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__77_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__77_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__77_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__77_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__77_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__77_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__77_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__77_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__70_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__70_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__70_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__70_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__70_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__70_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__70_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__70_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__70_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__70_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__70_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__70_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__70_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__70_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__70_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__70_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__65_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__65_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_77_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_77_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_77_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_77_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_77_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_77_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_77_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_77_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_77_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_77_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_77_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_77_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_77_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_77_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_77_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_77_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_77_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_77_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_77_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_77_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_77_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_77_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_77_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_77_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_77_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_77_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_77_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_77_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_77_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_77_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_77_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_77_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_77_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_77_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_77_ccff_tail ) ) ;
grid_clb grid_clb_7__7_ (
    .prog_clk ( { ctsbuf_net_4312413 } ) ,
    .Test_en ( { BUF_net_505 } ) ,
    .clk ( { ctsbuf_net_212003 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_72_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_215_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__78_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__78_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__78_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__78_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__78_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__78_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__78_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__78_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__78_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__78_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__78_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__78_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__78_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__78_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__78_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__78_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__71_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__71_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__71_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__71_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__71_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__71_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__71_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__71_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__71_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__71_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__71_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__71_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__71_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__71_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__71_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__71_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__66_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__66_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_78_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_78_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_78_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_78_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_78_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_78_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_78_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_78_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_78_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_78_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_78_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_78_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_78_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_78_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_78_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_78_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_78_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_78_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_78_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_78_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_78_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_78_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_78_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_78_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_78_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_78_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_78_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_78_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_78_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_78_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_78_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_78_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_78_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_78_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_78_ccff_tail ) ) ;
grid_clb grid_clb_7__8_ (
    .prog_clk ( { ctsbuf_net_3852367 } ) ,
    .Test_en ( { BUF_net_1521 } ) ,
    .clk ( { ctsbuf_net_262008 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_73_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_216_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__79_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__79_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__79_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__79_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__79_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__79_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__79_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__79_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__79_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__79_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__79_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__79_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__79_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__79_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__79_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__79_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__72_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__72_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__72_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__72_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__72_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__72_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__72_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__72_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__72_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__72_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__72_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__72_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__72_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__72_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__72_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__72_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__67_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__67_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_79_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_79_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_79_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_79_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_79_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_79_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_79_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_79_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_79_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_79_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_79_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_79_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_79_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_79_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_79_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_79_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_79_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_79_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_79_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_79_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_79_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_79_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_79_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_79_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_79_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_79_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_79_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_79_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_79_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_79_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_79_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_79_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_79_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_79_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_79_ccff_tail ) ) ;
grid_clb grid_clb_7__9_ (
    .prog_clk ( { ctsbuf_net_3402322 } ) ,
    .Test_en ( { BUF_net_1729 } ) ,
    .clk ( { ctsbuf_net_262008 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_74_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_217_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__80_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__80_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__80_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__80_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__80_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__80_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__80_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__80_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__80_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__80_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__80_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__80_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__80_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__80_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__80_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__80_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__73_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__73_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__73_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__73_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__73_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__73_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__73_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__73_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__73_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__73_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__73_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__73_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__73_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__73_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__73_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__73_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__68_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__68_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_80_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_80_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_80_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_80_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_80_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_80_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_80_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_80_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_80_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_80_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_80_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_80_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_80_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_80_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_80_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_80_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_80_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_80_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_80_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_80_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_80_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_80_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_80_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_80_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_80_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_80_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_80_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_80_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_80_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_80_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_80_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_80_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_80_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_80_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_80_ccff_tail ) ) ;
grid_clb grid_clb_7__10_ (
    .prog_clk ( { ctsbuf_net_2932275 } ) ,
    .Test_en ( { BUF_net_1523 } ) ,
    .clk ( { ctsbuf_net_272009 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_75_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_218_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__81_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__81_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__81_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__81_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__81_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__81_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__81_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__81_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__81_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__81_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__81_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__81_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__81_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__81_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__81_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__81_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__74_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__74_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__74_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__74_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__74_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__74_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__74_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__74_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__74_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__74_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__74_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__74_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__74_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__74_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__74_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__74_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__69_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__69_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_81_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_81_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_81_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_81_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_81_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_81_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_81_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_81_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_81_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_81_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_81_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_81_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_81_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_81_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_81_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_81_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_81_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_81_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_81_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_81_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_81_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_81_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_81_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_81_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_81_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_81_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_81_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_81_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_81_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_81_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_81_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_81_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_81_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_81_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_81_ccff_tail ) ) ;
grid_clb grid_clb_7__11_ (
    .prog_clk ( { ctsbuf_net_2472229 } ) ,
    .Test_en ( { BUF_net_1726 } ) ,
    .clk ( { ctsbuf_net_272009 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_76_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_219_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__82_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__82_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__82_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__82_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__82_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__82_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__82_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__82_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__82_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__82_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__82_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__82_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__82_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__82_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__82_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__82_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__75_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__75_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__75_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__75_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__75_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__75_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__75_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__75_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__75_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__75_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__75_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__75_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__75_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__75_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__75_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__75_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__70_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__70_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_82_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_82_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_82_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_82_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_82_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_82_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_82_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_82_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_82_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_82_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_82_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_82_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_82_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_82_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_82_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_82_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_82_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_82_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_82_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_82_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_82_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_82_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_82_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_82_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_82_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_82_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_82_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_82_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_82_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_82_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_82_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_82_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_82_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_82_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_82_ccff_tail ) ) ;
grid_clb grid_clb_7__12_ (
    .prog_clk ( { ctsbuf_net_2002182 } ) ,
    .Test_en ( { BUF_net_500 } ) ,
    .clk ( { ctsbuf_net_292011 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_137_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_280_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__83_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__83_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__83_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__83_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__83_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__83_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__83_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__83_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__83_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__83_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__83_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__83_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__83_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__83_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__83_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__83_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__76_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__76_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__76_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__76_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__76_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__76_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__76_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__76_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__76_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__76_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__76_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__76_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__76_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__76_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__76_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__76_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__71_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__71_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_83_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_83_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_83_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_83_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_83_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_83_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_83_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_83_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_83_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_83_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_83_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_83_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_83_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_83_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_83_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_83_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_83_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_83_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_83_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_83_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_83_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_83_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_83_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_83_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_83_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_83_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_83_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_83_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_83_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_83_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_83_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_83_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_83_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_83_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_83_ccff_tail ) ) ;
grid_clb grid_clb_8__1_ (
    .prog_clk ( { ctsbuf_net_1382120 } ) ,
    .Test_en ( { BUF_net_499 } ) ,
    .clk ( { ctsbuf_net_61988 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_77_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_220_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__84_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__84_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__84_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__84_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__84_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__84_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__84_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__84_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__84_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__84_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__84_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__84_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__84_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__84_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__84_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__84_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__0__7_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__0__7_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__0__7_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__0__7_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__0__7_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__0__7_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__0__7_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__0__7_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__0__7_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__0__7_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__0__7_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__0__7_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__0__7_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__0__7_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__0__7_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__0__7_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__72_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__72_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_84_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_84_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_84_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_84_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_84_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_84_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_84_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_84_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_84_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_84_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_84_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_84_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_84_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_84_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_84_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_84_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_84_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_84_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_84_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_84_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_84_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_84_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_84_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_84_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_84_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_84_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_84_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_84_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_84_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_84_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_84_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_84_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_84_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_84_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_84_ccff_tail ) ) ;
grid_clb grid_clb_8__2_ (
    .prog_clk ( { ctsbuf_net_1782160 } ) ,
    .Test_en ( { BUF_net_1635 } ) ,
    .clk ( { ctsbuf_net_61988 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_78_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_221_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__85_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__85_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__85_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__85_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__85_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__85_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__85_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__85_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__85_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__85_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__85_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__85_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__85_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__85_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__85_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__85_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__77_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__77_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__77_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__77_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__77_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__77_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__77_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__77_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__77_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__77_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__77_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__77_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__77_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__77_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__77_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__77_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__73_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__73_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_85_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_85_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_85_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_85_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_85_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_85_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_85_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_85_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_85_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_85_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_85_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_85_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_85_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_85_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_85_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_85_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_85_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_85_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_85_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_85_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_85_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_85_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_85_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_85_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_85_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_85_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_85_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_85_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_85_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_85_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_85_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_85_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_85_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_85_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_85_ccff_tail ) ) ;
grid_clb grid_clb_8__3_ (
    .prog_clk ( { ctsbuf_net_2232205 } ) ,
    .Test_en ( { BUF_net_1380 } ) ,
    .clk ( { ctsbuf_net_111993 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_79_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_222_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__86_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__86_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__86_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__86_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__86_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__86_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__86_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__86_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__86_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__86_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__86_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__86_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__86_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__86_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__86_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__86_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__78_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__78_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__78_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__78_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__78_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__78_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__78_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__78_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__78_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__78_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__78_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__78_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__78_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__78_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__78_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__78_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__74_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__74_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_86_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_86_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_86_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_86_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_86_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_86_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_86_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_86_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_86_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_86_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_86_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_86_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_86_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_86_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_86_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_86_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_86_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_86_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_86_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_86_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_86_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_86_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_86_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_86_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_86_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_86_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_86_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_86_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_86_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_86_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_86_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_86_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_86_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_86_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_86_ccff_tail ) ) ;
grid_clb grid_clb_8__4_ (
    .prog_clk ( { ctsbuf_net_2692251 } ) ,
    .Test_en ( { BUF_net_1570 } ) ,
    .clk ( { ctsbuf_net_111993 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_80_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_223_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__87_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__87_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__87_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__87_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__87_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__87_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__87_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__87_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__87_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__87_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__87_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__87_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__87_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__87_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__87_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__87_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__79_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__79_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__79_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__79_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__79_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__79_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__79_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__79_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__79_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__79_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__79_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__79_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__79_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__79_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__79_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__79_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__75_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__75_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_87_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_87_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_87_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_87_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_87_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_87_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_87_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_87_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_87_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_87_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_87_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_87_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_87_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_87_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_87_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_87_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_87_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_87_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_87_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_87_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_87_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_87_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_87_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_87_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_87_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_87_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_87_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_87_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_87_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_87_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_87_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_87_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_87_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_87_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_87_ccff_tail ) ) ;
grid_clb grid_clb_8__5_ (
    .prog_clk ( { ctsbuf_net_3152297 } ) ,
    .Test_en ( { BUF_net_1714 } ) ,
    .clk ( { ctsbuf_net_161998 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_81_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_224_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__88_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__88_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__88_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__88_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__88_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__88_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__88_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__88_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__88_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__88_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__88_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__88_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__88_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__88_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__88_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__88_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__80_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__80_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__80_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__80_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__80_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__80_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__80_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__80_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__80_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__80_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__80_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__80_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__80_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__80_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__80_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__80_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__76_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__76_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_88_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_88_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_88_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_88_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_88_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_88_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_88_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_88_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_88_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_88_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_88_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_88_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_88_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_88_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_88_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_88_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_88_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_88_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_88_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_88_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_88_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_88_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_88_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_88_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_88_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_88_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_88_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_88_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_88_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_88_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_88_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_88_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_88_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_88_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_88_ccff_tail ) ) ;
grid_clb grid_clb_8__6_ (
    .prog_clk ( { ctsbuf_net_3602342 } ) ,
    .Test_en ( { BUF_net_494 } ) ,
    .clk ( { ctsbuf_net_161998 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_82_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_225_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__89_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__89_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__89_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__89_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__89_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__89_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__89_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__89_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__89_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__89_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__89_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__89_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__89_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__89_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__89_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__89_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__81_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__81_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__81_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__81_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__81_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__81_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__81_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__81_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__81_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__81_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__81_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__81_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__81_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__81_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__81_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__81_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__77_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__77_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_89_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_89_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_89_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_89_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_89_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_89_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_89_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_89_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_89_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_89_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_89_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_89_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_89_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_89_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_89_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_89_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_89_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_89_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_89_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_89_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_89_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_89_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_89_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_89_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_89_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_89_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_89_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_89_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_89_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_89_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_89_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_89_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_89_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_89_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_89_ccff_tail ) ) ;
grid_clb grid_clb_8__7_ (
    .prog_clk ( { ctsbuf_net_3862368 } ) ,
    .Test_en ( { BUF_net_1665 } ) ,
    .clk ( { ctsbuf_net_212003 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_83_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_226_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__90_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__90_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__90_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__90_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__90_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__90_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__90_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__90_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__90_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__90_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__90_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__90_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__90_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__90_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__90_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__90_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__82_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__82_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__82_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__82_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__82_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__82_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__82_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__82_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__82_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__82_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__82_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__82_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__82_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__82_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__82_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__82_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__78_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__78_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_90_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_90_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_90_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_90_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_90_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_90_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_90_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_90_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_90_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_90_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_90_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_90_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_90_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_90_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_90_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_90_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_90_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_90_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_90_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_90_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_90_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_90_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_90_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_90_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_90_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_90_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_90_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_90_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_90_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_90_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_90_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_90_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_90_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_90_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_90_ccff_tail ) ) ;
grid_clb grid_clb_8__8_ (
    .prog_clk ( { p_abuf15 } ) ,
    .Test_en ( { BUF_net_1381 } ) ,
    .clk ( { ctsbuf_net_212003 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_84_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_227_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__91_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__91_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__91_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__91_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__91_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__91_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__91_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__91_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__91_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__91_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__91_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__91_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__91_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__91_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__91_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__91_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__83_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__83_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__83_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__83_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__83_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__83_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__83_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__83_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__83_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__83_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__83_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__83_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__83_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__83_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__83_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__83_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__79_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__79_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_91_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_91_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_91_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_91_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_91_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_91_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_91_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_91_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_91_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_91_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_91_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_91_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_91_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_91_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_91_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_91_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_91_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_91_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_91_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_91_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_91_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_91_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_91_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_91_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_91_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_91_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_91_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_91_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_91_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_91_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_91_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_91_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_91_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_91_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_91_ccff_tail ) ) ;
grid_clb grid_clb_8__9_ (
    .prog_clk ( { ctsbuf_net_2942276 } ) ,
    .Test_en ( { BUF_net_1631 } ) ,
    .clk ( { ctsbuf_net_262008 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_85_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_228_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__92_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__92_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__92_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__92_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__92_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__92_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__92_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__92_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__92_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__92_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__92_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__92_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__92_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__92_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__92_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__92_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__84_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__84_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__84_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__84_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__84_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__84_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__84_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__84_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__84_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__84_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__84_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__84_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__84_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__84_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__84_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__84_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__80_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__80_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_92_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_92_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_92_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_92_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_92_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_92_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_92_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_92_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_92_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_92_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_92_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_92_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_92_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_92_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_92_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_92_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_92_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_92_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_92_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_92_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_92_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_92_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_92_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_92_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_92_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_92_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_92_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_92_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_92_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_92_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_92_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_92_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_92_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_92_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_92_ccff_tail ) ) ;
grid_clb grid_clb_8__10_ (
    .prog_clk ( { ctsbuf_net_2492231 } ) ,
    .Test_en ( { BUF_net_1382 } ) ,
    .clk ( { ctsbuf_net_272009 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_86_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_229_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__93_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__93_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__93_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__93_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__93_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__93_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__93_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__93_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__93_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__93_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__93_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__93_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__93_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__93_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__93_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__93_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__85_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__85_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__85_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__85_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__85_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__85_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__85_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__85_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__85_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__85_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__85_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__85_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__85_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__85_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__85_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__85_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__81_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__81_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_93_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_93_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_93_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_93_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_93_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_93_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_93_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_93_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_93_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_93_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_93_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_93_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_93_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_93_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_93_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_93_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_93_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_93_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_93_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_93_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_93_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_93_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_93_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_93_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_93_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_93_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_93_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_93_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_93_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_93_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_93_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_93_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_93_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_93_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_93_ccff_tail ) ) ;
grid_clb grid_clb_8__11_ (
    .prog_clk ( { ctsbuf_net_2012183 } ) ,
    .Test_en ( { BUF_net_1634 } ) ,
    .clk ( { ctsbuf_net_272009 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_87_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_230_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__94_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__94_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__94_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__94_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__94_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__94_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__94_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__94_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__94_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__94_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__94_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__94_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__94_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__94_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__94_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__94_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__86_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__86_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__86_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__86_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__86_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__86_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__86_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__86_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__86_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__86_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__86_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__86_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__86_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__86_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__86_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__86_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__82_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__82_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_94_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_94_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_94_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_94_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_94_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_94_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_94_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_94_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_94_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_94_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_94_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_94_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_94_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_94_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_94_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_94_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_94_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_94_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_94_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_94_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_94_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_94_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_94_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_94_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_94_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_94_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_94_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_94_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_94_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_94_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_94_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_94_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_94_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_94_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_94_ccff_tail ) ) ;
grid_clb grid_clb_8__12_ (
    .prog_clk ( { ctsbuf_net_1592141 } ) ,
    .Test_en ( { BUF_net_488 } ) ,
    .clk ( { ctsbuf_net_292011 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_138_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_281_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__95_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__95_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__95_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__95_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__95_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__95_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__95_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__95_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__95_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__95_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__95_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__95_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__95_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__95_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__95_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__95_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__87_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__87_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__87_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__87_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__87_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__87_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__87_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__87_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__87_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__87_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__87_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__87_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__87_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__87_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__87_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__87_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__83_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__83_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_95_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_95_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_95_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_95_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_95_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_95_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_95_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_95_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_95_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_95_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_95_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_95_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_95_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_95_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_95_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_95_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_95_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_95_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_95_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_95_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_95_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_95_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_95_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_95_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_95_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_95_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_95_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_95_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_95_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_95_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_95_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_95_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_95_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_95_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_95_ccff_tail ) ) ;
grid_clb grid_clb_9__1_ (
    .prog_clk ( { ctsbuf_net_1072089 } ) ,
    .Test_en ( { BUF_net_487 } ) ,
    .clk ( { ctsbuf_net_61988 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_88_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_231_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__96_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__96_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__96_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__96_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__96_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__96_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__96_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__96_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__96_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__96_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__96_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__96_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__96_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__96_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__96_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__96_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__0__8_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__0__8_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__0__8_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__0__8_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__0__8_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__0__8_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__0__8_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__0__8_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__0__8_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__0__8_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__0__8_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__0__8_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__0__8_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__0__8_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__0__8_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__0__8_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__84_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__84_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_96_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_96_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_96_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_96_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_96_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_96_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_96_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_96_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_96_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_96_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_96_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_96_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_96_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_96_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_96_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_96_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_96_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_96_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_96_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_96_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_96_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_96_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_96_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_96_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_96_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_96_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_96_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_96_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_96_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_96_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_96_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_96_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_96_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_96_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_96_ccff_tail ) ) ;
grid_clb grid_clb_9__2_ (
    .prog_clk ( { ctsbuf_net_1392121 } ) ,
    .Test_en ( { BUF_net_1445 } ) ,
    .clk ( { ctsbuf_net_31985 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_89_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_232_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__97_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__97_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__97_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__97_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__97_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__97_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__97_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__97_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__97_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__97_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__97_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__97_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__97_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__97_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__97_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__97_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__88_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__88_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__88_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__88_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__88_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__88_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__88_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__88_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__88_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__88_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__88_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__88_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__88_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__88_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__88_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__88_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__85_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__85_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_97_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_97_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_97_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_97_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_97_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_97_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_97_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_97_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_97_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_97_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_97_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_97_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_97_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_97_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_97_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_97_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_97_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_97_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_97_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_97_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_97_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_97_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_97_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_97_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_97_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_97_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_97_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_97_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_97_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_97_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_97_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_97_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_97_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_97_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_97_ccff_tail ) ) ;
grid_clb grid_clb_9__3_ (
    .prog_clk ( { ctsbuf_net_1792161 } ) ,
    .Test_en ( { BUF_net_1187 } ) ,
    .clk ( { ctsbuf_net_111993 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_90_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_233_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__98_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__98_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__98_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__98_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__98_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__98_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__98_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__98_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__98_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__98_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__98_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__98_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__98_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__98_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__98_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__98_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__89_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__89_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__89_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__89_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__89_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__89_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__89_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__89_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__89_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__89_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__89_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__89_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__89_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__89_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__89_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__89_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__86_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__86_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_98_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_98_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_98_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_98_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_98_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_98_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_98_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_98_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_98_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_98_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_98_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_98_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_98_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_98_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_98_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_98_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_98_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_98_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_98_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_98_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_98_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_98_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_98_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_98_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_98_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_98_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_98_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_98_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_98_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_98_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_98_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_98_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_98_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_98_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_98_ccff_tail ) ) ;
grid_clb grid_clb_9__4_ (
    .prog_clk ( { ctsbuf_net_2242206 } ) ,
    .Test_en ( { BUF_net_1447 } ) ,
    .clk ( { ctsbuf_net_111993 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_91_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_234_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__99_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__99_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__99_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__99_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__99_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__99_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__99_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__99_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__99_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__99_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__99_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__99_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__99_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__99_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__99_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__99_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__90_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__90_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__90_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__90_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__90_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__90_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__90_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__90_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__90_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__90_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__90_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__90_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__90_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__90_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__90_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__90_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__87_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__87_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_99_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_99_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_99_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_99_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_99_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_99_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_99_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_99_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_99_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_99_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_99_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_99_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_99_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_99_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_99_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_99_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_99_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_99_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_99_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_99_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_99_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_99_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_99_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_99_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_99_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_99_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_99_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_99_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_99_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_99_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_99_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_99_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_99_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_99_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_99_ccff_tail ) ) ;
grid_clb grid_clb_9__5_ (
    .prog_clk ( { ctsbuf_net_2702252 } ) ,
    .Test_en ( { BUF_net_1515 } ) ,
    .clk ( { ctsbuf_net_161998 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_92_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_235_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__100_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__100_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__100_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__100_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__100_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__100_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__100_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__100_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__100_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__100_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__100_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__100_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__100_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__100_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__100_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__100_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__91_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__91_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__91_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__91_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__91_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__91_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__91_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__91_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__91_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__91_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__91_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__91_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__91_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__91_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__91_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__91_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__88_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__88_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_100_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_100_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_100_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_100_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_100_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_100_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_100_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_100_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_100_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_100_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_100_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_100_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_100_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_100_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_100_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_100_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_100_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_100_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_100_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_100_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_100_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_100_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_100_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_100_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_100_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_100_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_100_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_100_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_100_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_100_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_100_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_100_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_100_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_100_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_100_ccff_tail ) ) ;
grid_clb grid_clb_9__6_ (
    .prog_clk ( { ctsbuf_net_3162298 } ) ,
    .Test_en ( { BUF_net_482 } ) ,
    .clk ( { ctsbuf_net_161998 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_93_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_236_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__101_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__101_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__101_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__101_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__101_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__101_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__101_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__101_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__101_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__101_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__101_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__101_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__101_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__101_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__101_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__101_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__92_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__92_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__92_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__92_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__92_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__92_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__92_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__92_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__92_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__92_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__92_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__92_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__92_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__92_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__92_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__92_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__89_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__89_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_101_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_101_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_101_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_101_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_101_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_101_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_101_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_101_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_101_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_101_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_101_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_101_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_101_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_101_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_101_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_101_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_101_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_101_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_101_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_101_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_101_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_101_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_101_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_101_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_101_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_101_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_101_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_101_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_101_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_101_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_101_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_101_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_101_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_101_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_101_ccff_tail ) ) ;
grid_clb grid_clb_9__7_ (
    .prog_clk ( { ctsbuf_net_3442326 } ) ,
    .Test_en ( { BUF_net_1460 } ) ,
    .clk ( { ctsbuf_net_212003 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_94_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_237_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__102_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__102_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__102_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__102_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__102_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__102_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__102_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__102_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__102_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__102_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__102_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__102_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__102_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__102_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__102_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__102_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__93_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__93_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__93_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__93_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__93_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__93_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__93_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__93_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__93_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__93_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__93_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__93_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__93_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__93_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__93_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__93_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__90_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__90_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_102_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_102_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_102_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_102_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_102_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_102_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_102_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_102_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_102_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_102_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_102_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_102_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_102_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_102_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_102_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_102_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_102_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_102_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_102_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_102_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_102_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_102_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_102_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_102_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_102_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_102_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_102_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_102_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_102_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_102_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_102_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_102_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_102_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_102_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_102_ccff_tail ) ) ;
grid_clb grid_clb_9__8_ (
    .prog_clk ( { ctsbuf_net_2962278 } ) ,
    .Test_en ( { BUF_net_1192 } ) ,
    .clk ( { ctsbuf_net_212003 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_95_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_238_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__103_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__103_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__103_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__103_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__103_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__103_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__103_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__103_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__103_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__103_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__103_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__103_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__103_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__103_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__103_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__103_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__94_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__94_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__94_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__94_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__94_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__94_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__94_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__94_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__94_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__94_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__94_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__94_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__94_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__94_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__94_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__94_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__91_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__91_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_103_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_103_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_103_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_103_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_103_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_103_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_103_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_103_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_103_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_103_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_103_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_103_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_103_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_103_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_103_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_103_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_103_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_103_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_103_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_103_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_103_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_103_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_103_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_103_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_103_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_103_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_103_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_103_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_103_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_103_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_103_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_103_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_103_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_103_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_103_ccff_tail ) ) ;
grid_clb grid_clb_9__9_ (
    .prog_clk ( { ctsbuf_net_2502232 } ) ,
    .Test_en ( { BUF_net_1462 } ) ,
    .clk ( { ctsbuf_net_222004 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_96_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_239_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__104_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__104_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__104_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__104_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__104_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__104_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__104_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__104_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__104_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__104_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__104_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__104_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__104_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__104_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__104_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__104_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__95_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__95_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__95_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__95_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__95_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__95_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__95_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__95_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__95_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__95_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__95_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__95_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__95_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__95_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__95_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__95_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__92_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__92_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_104_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_104_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_104_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_104_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_104_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_104_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_104_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_104_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_104_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_104_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_104_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_104_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_104_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_104_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_104_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_104_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_104_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_104_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_104_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_104_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_104_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_104_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_104_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_104_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_104_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_104_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_104_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_104_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_104_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_104_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_104_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_104_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_104_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_104_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_104_ccff_tail ) ) ;
grid_clb grid_clb_9__10_ (
    .prog_clk ( { ctsbuf_net_2032185 } ) ,
    .Test_en ( { BUF_net_1195 } ) ,
    .clk ( { ctsbuf_net_272009 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_97_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_240_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__105_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__105_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__105_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__105_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__105_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__105_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__105_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__105_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__105_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__105_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__105_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__105_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__105_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__105_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__105_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__105_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__96_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__96_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__96_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__96_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__96_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__96_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__96_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__96_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__96_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__96_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__96_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__96_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__96_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__96_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__96_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__96_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__93_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__93_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_105_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_105_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_105_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_105_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_105_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_105_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_105_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_105_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_105_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_105_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_105_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_105_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_105_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_105_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_105_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_105_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_105_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_105_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_105_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_105_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_105_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_105_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_105_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_105_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_105_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_105_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_105_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_105_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_105_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_105_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_105_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_105_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_105_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_105_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_105_ccff_tail ) ) ;
grid_clb grid_clb_9__11_ (
    .prog_clk ( { ctsbuf_net_1602142 } ) ,
    .Test_en ( { BUF_net_1466 } ) ,
    .clk ( { ctsbuf_net_272009 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_98_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_241_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__106_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__106_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__106_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__106_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__106_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__106_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__106_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__106_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__106_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__106_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__106_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__106_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__106_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__106_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__106_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__106_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__97_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__97_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__97_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__97_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__97_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__97_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__97_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__97_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__97_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__97_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__97_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__97_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__97_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__97_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__97_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__97_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__94_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__94_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_106_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_106_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_106_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_106_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_106_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_106_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_106_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_106_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_106_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_106_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_106_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_106_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_106_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_106_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_106_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_106_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_106_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_106_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_106_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_106_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_106_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_106_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_106_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_106_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_106_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_106_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_106_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_106_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_106_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_106_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_106_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_106_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_106_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_106_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_106_ccff_tail ) ) ;
grid_clb grid_clb_9__12_ (
    .prog_clk ( { ctsbuf_net_1252107 } ) ,
    .Test_en ( { BUF_net_476 } ) ,
    .clk ( { ctsbuf_net_292011 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_139_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_282_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__107_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__107_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__107_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__107_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__107_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__107_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__107_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__107_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__107_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__107_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__107_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__107_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__107_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__107_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__107_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__107_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__98_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__98_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__98_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__98_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__98_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__98_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__98_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__98_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__98_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__98_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__98_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__98_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__98_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__98_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__98_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__98_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__95_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__95_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_107_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_107_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_107_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_107_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_107_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_107_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_107_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_107_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_107_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_107_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_107_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_107_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_107_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_107_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_107_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_107_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_107_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_107_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_107_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_107_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_107_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_107_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_107_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_107_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_107_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_107_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_107_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_107_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_107_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_107_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_107_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_107_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_107_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_107_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_107_ccff_tail ) ) ;
grid_clb grid_clb_10__1_ (
    .prog_clk ( { ctsbuf_net_802062 } ) ,
    .Test_en ( { BUF_net_475 } ) ,
    .clk ( { ctsbuf_net_11983 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_99_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_242_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__108_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__108_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__108_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__108_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__108_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__108_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__108_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__108_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__108_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__108_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__108_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__108_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__108_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__108_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__108_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__108_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__0__9_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__0__9_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__0__9_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__0__9_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__0__9_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__0__9_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__0__9_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__0__9_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__0__9_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__0__9_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__0__9_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__0__9_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__0__9_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__0__9_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__0__9_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__0__9_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__96_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__96_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_108_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_108_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_108_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_108_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_108_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_108_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_108_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_108_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_108_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_108_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_108_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_108_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_108_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_108_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_108_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_108_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_108_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_108_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_108_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_108_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_108_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_108_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_108_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_108_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_108_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_108_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_108_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_108_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_108_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_108_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_108_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_108_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_108_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_108_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_108_ccff_tail ) ) ;
grid_clb grid_clb_10__2_ (
    .prog_clk ( { ctsbuf_net_1082090 } ) ,
    .Test_en ( { BUF_net_1197 } ) ,
    .clk ( { ctsbuf_net_31985 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_100_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_243_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__109_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__109_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__109_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__109_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__109_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__109_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__109_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__109_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__109_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__109_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__109_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__109_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__109_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__109_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__109_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__109_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__99_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__99_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__99_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__99_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__99_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__99_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__99_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__99_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__99_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__99_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__99_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__99_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__99_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__99_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__99_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__99_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__97_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__97_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_109_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_109_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_109_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_109_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_109_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_109_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_109_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_109_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_109_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_109_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_109_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_109_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_109_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_109_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_109_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_109_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_109_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_109_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_109_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_109_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_109_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_109_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_109_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_109_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_109_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_109_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_109_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_109_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_109_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_109_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_109_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_109_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_109_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_109_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_109_ccff_tail ) ) ;
grid_clb grid_clb_10__3_ (
    .prog_clk ( { ctsbuf_net_1402122 } ) ,
    .Test_en ( { BUF_net_967 } ) ,
    .clk ( { ctsbuf_net_41986 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_101_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_244_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__110_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__110_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__110_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__110_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__110_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__110_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__110_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__110_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__110_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__110_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__110_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__110_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__110_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__110_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__110_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__110_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__100_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__100_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__100_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__100_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__100_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__100_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__100_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__100_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__100_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__100_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__100_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__100_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__100_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__100_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__100_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__100_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__98_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__98_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_110_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_110_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_110_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_110_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_110_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_110_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_110_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_110_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_110_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_110_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_110_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_110_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_110_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_110_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_110_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_110_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_110_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_110_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_110_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_110_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_110_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_110_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_110_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_110_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_110_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_110_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_110_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_110_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_110_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_110_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_110_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_110_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_110_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_110_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_110_ccff_tail ) ) ;
grid_clb grid_clb_10__4_ (
    .prog_clk ( { ctsbuf_net_1802162 } ) ,
    .Test_en ( { BUF_net_1199 } ) ,
    .clk ( { ctsbuf_net_111993 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_102_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_245_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__111_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__111_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__111_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__111_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__111_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__111_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__111_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__111_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__111_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__111_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__111_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__111_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__111_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__111_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__111_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__111_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__101_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__101_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__101_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__101_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__101_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__101_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__101_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__101_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__101_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__101_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__101_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__101_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__101_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__101_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__101_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__101_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__99_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__99_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_111_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_111_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_111_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_111_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_111_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_111_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_111_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_111_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_111_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_111_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_111_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_111_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_111_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_111_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_111_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_111_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_111_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_111_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_111_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_111_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_111_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_111_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_111_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_111_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_111_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_111_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_111_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_111_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_111_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_111_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_111_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_111_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_111_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_111_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_111_ccff_tail ) ) ;
grid_clb grid_clb_10__5_ (
    .prog_clk ( { ctsbuf_net_2252207 } ) ,
    .Test_en ( { BUF_net_1189 } ) ,
    .clk ( { ctsbuf_net_91991 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_103_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_246_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__112_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__112_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__112_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__112_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__112_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__112_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__112_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__112_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__112_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__112_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__112_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__112_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__112_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__112_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__112_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__112_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__102_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__102_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__102_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__102_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__102_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__102_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__102_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__102_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__102_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__102_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__102_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__102_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__102_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__102_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__102_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__102_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__100_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__100_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_112_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_112_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_112_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_112_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_112_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_112_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_112_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_112_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_112_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_112_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_112_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_112_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_112_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_112_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_112_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_112_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_112_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_112_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_112_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_112_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_112_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_112_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_112_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_112_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_112_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_112_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_112_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_112_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_112_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_112_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_112_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_112_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_112_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_112_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_112_ccff_tail ) ) ;
grid_clb grid_clb_10__6_ (
    .prog_clk ( { ctsbuf_net_2712253 } ) ,
    .Test_en ( { BUF_net_470 } ) ,
    .clk ( { ctsbuf_net_161998 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_104_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_247_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__113_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__113_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__113_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__113_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__113_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__113_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__113_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__113_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__113_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__113_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__113_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__113_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__113_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__113_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__113_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__113_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__103_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__103_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__103_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__103_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__103_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__103_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__103_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__103_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__103_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__103_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__103_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__103_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__103_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__103_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__103_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__103_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__101_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__101_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_113_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_113_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_113_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_113_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_113_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_113_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_113_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_113_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_113_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_113_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_113_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_113_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_113_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_113_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_113_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_113_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_113_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_113_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_113_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_113_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_113_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_113_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_113_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_113_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_113_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_113_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_113_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_113_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_113_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_113_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_113_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_113_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_113_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_113_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_113_ccff_tail ) ) ;
grid_clb grid_clb_10__7_ (
    .prog_clk ( { ctsbuf_net_2982280 } ) ,
    .Test_en ( { BUF_net_1190 } ) ,
    .clk ( { ctsbuf_net_141996 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_105_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_248_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__114_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__114_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__114_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__114_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__114_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__114_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__114_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__114_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__114_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__114_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__114_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__114_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__114_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__114_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__114_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__114_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__104_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__104_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__104_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__104_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__104_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__104_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__104_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__104_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__104_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__104_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__104_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__104_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__104_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__104_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__104_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__104_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__102_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__102_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_114_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_114_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_114_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_114_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_114_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_114_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_114_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_114_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_114_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_114_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_114_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_114_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_114_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_114_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_114_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_114_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_114_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_114_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_114_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_114_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_114_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_114_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_114_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_114_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_114_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_114_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_114_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_114_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_114_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_114_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_114_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_114_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_114_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_114_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_114_ccff_tail ) ) ;
grid_clb grid_clb_10__8_ (
    .prog_clk ( { ctsbuf_net_2522234 } ) ,
    .Test_en ( { BUF_net_976 } ) ,
    .clk ( { ctsbuf_net_212003 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_106_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_249_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__115_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__115_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__115_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__115_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__115_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__115_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__115_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__115_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__115_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__115_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__115_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__115_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__115_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__115_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__115_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__115_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__105_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__105_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__105_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__105_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__105_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__105_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__105_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__105_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__105_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__105_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__105_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__105_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__105_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__105_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__105_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__105_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__103_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__103_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_115_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_115_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_115_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_115_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_115_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_115_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_115_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_115_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_115_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_115_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_115_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_115_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_115_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_115_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_115_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_115_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_115_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_115_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_115_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_115_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_115_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_115_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_115_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_115_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_115_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_115_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_115_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_115_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_115_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_115_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_115_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_115_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_115_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_115_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_115_ccff_tail ) ) ;
grid_clb grid_clb_10__9_ (
    .prog_clk ( { ctsbuf_net_2042186 } ) ,
    .Test_en ( { BUF_net_1207 } ) ,
    .clk ( { ctsbuf_net_171999 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_107_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_250_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__116_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__116_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__116_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__116_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__116_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__116_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__116_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__116_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__116_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__116_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__116_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__116_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__116_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__116_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__116_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__116_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__106_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__106_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__106_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__106_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__106_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__106_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__106_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__106_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__106_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__106_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__106_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__106_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__106_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__106_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__106_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__106_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__104_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__104_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_116_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_116_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_116_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_116_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_116_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_116_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_116_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_116_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_116_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_116_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_116_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_116_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_116_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_116_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_116_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_116_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_116_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_116_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_116_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_116_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_116_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_116_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_116_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_116_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_116_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_116_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_116_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_116_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_116_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_116_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_116_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_116_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_116_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_116_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_116_ccff_tail ) ) ;
grid_clb grid_clb_10__10_ (
    .prog_clk ( { ctsbuf_net_1622144 } ) ,
    .Test_en ( { BUF_net_980 } ) ,
    .clk ( { ctsbuf_net_222004 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_108_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_251_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__117_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__117_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__117_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__117_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__117_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__117_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__117_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__117_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__117_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__117_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__117_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__117_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__117_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__117_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__117_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__117_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__107_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__107_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__107_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__107_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__107_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__107_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__107_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__107_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__107_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__107_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__107_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__107_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__107_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__107_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__107_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__107_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__105_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__105_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_117_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_117_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_117_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_117_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_117_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_117_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_117_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_117_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_117_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_117_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_117_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_117_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_117_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_117_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_117_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_117_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_117_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_117_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_117_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_117_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_117_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_117_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_117_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_117_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_117_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_117_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_117_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_117_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_117_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_117_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_117_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_117_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_117_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_117_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_117_ccff_tail ) ) ;
grid_clb grid_clb_10__11_ (
    .prog_clk ( { ctsbuf_net_1262108 } ) ,
    .Test_en ( { BUF_net_1210 } ) ,
    .clk ( { ctsbuf_net_242006 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_109_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_252_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__118_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__118_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__118_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__118_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__118_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__118_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__118_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__118_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__118_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__118_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__118_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__118_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__118_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__118_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__118_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__118_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__108_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__108_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__108_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__108_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__108_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__108_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__108_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__108_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__108_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__108_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__108_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__108_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__108_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__108_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__108_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__108_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__106_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__106_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_118_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_118_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_118_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_118_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_118_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_118_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_118_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_118_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_118_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_118_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_118_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_118_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_118_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_118_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_118_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_118_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_118_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_118_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_118_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_118_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_118_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_118_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_118_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_118_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_118_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_118_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_118_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_118_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_118_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_118_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_118_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_118_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_118_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_118_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_118_ccff_tail ) ) ;
grid_clb grid_clb_10__12_ (
    .prog_clk ( { ctsbuf_net_972079 } ) ,
    .Test_en ( { BUF_net_464 } ) ,
    .clk ( { ctsbuf_net_292011 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_140_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_283_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__119_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__119_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__119_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__119_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__119_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__119_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__119_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__119_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__119_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__119_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__119_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__119_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__119_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__119_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__119_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__119_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__109_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__109_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__109_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__109_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__109_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__109_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__109_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__109_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__109_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__109_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__109_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__109_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__109_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__109_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__109_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__109_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__107_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__107_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_119_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_119_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_119_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_119_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_119_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_119_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_119_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_119_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_119_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_119_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_119_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_119_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_119_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_119_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_119_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_119_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_119_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_119_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_119_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_119_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_119_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_119_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_119_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_119_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_119_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_119_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_119_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_119_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_119_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_119_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_119_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_119_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_119_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_119_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_119_ccff_tail ) ) ;
grid_clb grid_clb_11__1_ (
    .prog_clk ( { ctsbuf_net_612043 } ) ,
    .Test_en ( { BUF_net_463 } ) ,
    .clk ( { ctsbuf_net_11983 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_110_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_253_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__120_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__120_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__120_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__120_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__120_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__120_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__120_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__120_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__120_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__120_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__120_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__120_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__120_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__120_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__120_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__120_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__0__10_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__0__10_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__0__10_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__0__10_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__0__10_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__0__10_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__0__10_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__0__10_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__0__10_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__0__10_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__0__10_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__0__10_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__0__10_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__0__10_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__0__10_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__0__10_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__108_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__108_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_120_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_120_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_120_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_120_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_120_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_120_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_120_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_120_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_120_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_120_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_120_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_120_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_120_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_120_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_120_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_120_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_120_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_120_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_120_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_120_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_120_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_120_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_120_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_120_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_120_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_120_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_120_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_120_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_120_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_120_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_120_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_120_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_120_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_120_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_120_ccff_tail ) ) ;
grid_clb grid_clb_11__2_ (
    .prog_clk ( { ctsbuf_net_812063 } ) ,
    .Test_en ( { BUF_net_847 } ) ,
    .clk ( { ctsbuf_net_31985 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_111_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_254_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__121_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__121_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__121_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__121_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__121_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__121_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__121_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__121_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__121_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__121_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__121_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__121_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__121_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__121_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__121_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__121_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__110_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__110_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__110_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__110_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__110_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__110_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__110_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__110_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__110_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__110_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__110_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__110_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__110_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__110_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__110_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__110_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__109_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__109_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_121_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_121_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_121_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_121_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_121_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_121_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_121_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_121_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_121_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_121_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_121_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_121_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_121_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_121_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_121_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_121_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_121_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_121_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_121_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_121_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_121_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_121_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_121_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_121_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_121_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_121_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_121_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_121_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_121_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_121_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_121_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_121_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_121_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_121_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_121_ccff_tail ) ) ;
grid_clb grid_clb_11__3_ (
    .prog_clk ( { ctsbuf_net_1092091 } ) ,
    .Test_en ( { BUF_net_719 } ) ,
    .clk ( { ctsbuf_net_31985 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_112_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_255_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__122_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__122_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__122_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__122_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__122_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__122_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__122_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__122_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__122_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__122_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__122_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__122_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__122_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__122_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__122_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__122_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__111_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__111_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__111_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__111_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__111_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__111_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__111_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__111_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__111_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__111_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__111_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__111_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__111_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__111_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__111_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__111_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__110_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__110_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_122_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_122_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_122_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_122_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_122_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_122_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_122_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_122_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_122_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_122_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_122_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_122_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_122_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_122_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_122_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_122_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_122_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_122_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_122_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_122_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_122_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_122_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_122_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_122_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_122_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_122_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_122_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_122_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_122_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_122_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_122_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_122_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_122_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_122_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_122_ccff_tail ) ) ;
grid_clb grid_clb_11__4_ (
    .prog_clk ( { ctsbuf_net_1412123 } ) ,
    .Test_en ( { BUF_net_848 } ) ,
    .clk ( { ctsbuf_net_41986 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_113_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_256_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__123_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__123_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__123_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__123_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__123_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__123_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__123_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__123_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__123_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__123_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__123_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__123_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__123_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__123_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__123_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__123_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__112_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__112_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__112_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__112_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__112_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__112_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__112_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__112_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__112_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__112_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__112_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__112_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__112_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__112_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__112_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__112_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__111_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__111_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_123_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_123_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_123_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_123_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_123_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_123_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_123_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_123_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_123_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_123_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_123_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_123_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_123_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_123_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_123_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_123_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_123_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_123_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_123_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_123_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_123_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_123_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_123_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_123_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_123_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_123_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_123_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_123_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_123_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_123_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_123_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_123_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_123_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_123_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_123_ccff_tail ) ) ;
grid_clb grid_clb_11__5_ (
    .prog_clk ( { ctsbuf_net_1812163 } ) ,
    .Test_en ( { BUF_net_850 } ) ,
    .clk ( { ctsbuf_net_91991 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_114_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_257_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__124_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__124_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__124_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__124_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__124_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__124_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__124_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__124_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__124_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__124_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__124_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__124_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__124_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__124_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__124_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__124_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__113_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__113_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__113_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__113_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__113_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__113_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__113_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__113_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__113_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__113_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__113_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__113_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__113_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__113_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__113_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__113_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__112_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__112_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_124_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_124_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_124_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_124_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_124_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_124_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_124_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_124_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_124_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_124_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_124_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_124_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_124_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_124_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_124_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_124_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_124_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_124_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_124_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_124_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_124_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_124_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_124_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_124_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_124_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_124_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_124_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_124_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_124_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_124_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_124_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_124_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_124_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_124_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_124_ccff_tail ) ) ;
grid_clb grid_clb_11__6_ (
    .prog_clk ( { ctsbuf_net_2262208 } ) ,
    .Test_en ( { BUF_net_458 } ) ,
    .clk ( { ctsbuf_net_91991 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_115_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_258_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__125_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__125_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__125_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__125_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__125_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__125_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__125_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__125_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__125_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__125_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__125_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__125_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__125_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__125_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__125_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__125_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__114_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__114_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__114_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__114_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__114_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__114_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__114_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__114_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__114_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__114_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__114_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__114_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__114_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__114_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__114_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__114_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__113_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__113_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_125_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_125_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_125_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_125_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_125_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_125_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_125_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_125_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_125_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_125_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_125_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_125_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_125_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_125_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_125_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_125_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_125_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_125_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_125_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_125_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_125_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_125_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_125_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_125_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_125_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_125_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_125_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_125_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_125_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_125_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_125_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_125_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_125_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_125_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_125_ccff_tail ) ) ;
grid_clb grid_clb_11__7_ (
    .prog_clk ( { ctsbuf_net_2542236 } ) ,
    .Test_en ( { BUF_net_852 } ) ,
    .clk ( { ctsbuf_net_141996 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_116_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_259_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__126_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__126_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__126_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__126_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__126_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__126_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__126_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__126_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__126_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__126_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__126_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__126_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__126_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__126_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__126_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__126_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__115_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__115_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__115_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__115_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__115_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__115_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__115_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__115_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__115_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__115_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__115_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__115_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__115_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__115_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__115_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__115_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__114_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__114_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_126_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_126_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_126_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_126_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_126_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_126_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_126_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_126_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_126_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_126_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_126_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_126_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_126_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_126_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_126_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_126_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_126_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_126_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_126_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_126_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_126_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_126_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_126_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_126_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_126_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_126_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_126_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_126_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_126_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_126_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_126_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_126_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_126_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_126_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_126_ccff_tail ) ) ;
grid_clb grid_clb_11__8_ (
    .prog_clk ( { ctsbuf_net_2062188 } ) ,
    .Test_en ( { BUF_net_727 } ) ,
    .clk ( { ctsbuf_net_141996 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_117_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_260_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__127_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__127_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__127_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__127_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__127_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__127_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__127_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__127_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__127_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__127_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__127_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__127_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__127_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__127_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__127_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__127_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__116_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__116_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__116_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__116_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__116_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__116_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__116_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__116_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__116_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__116_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__116_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__116_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__116_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__116_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__116_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__116_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__115_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__115_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_127_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_127_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_127_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_127_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_127_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_127_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_127_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_127_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_127_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_127_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_127_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_127_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_127_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_127_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_127_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_127_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_127_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_127_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_127_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_127_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_127_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_127_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_127_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_127_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_127_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_127_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_127_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_127_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_127_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_127_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_127_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_127_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_127_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_127_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_127_ccff_tail ) ) ;
grid_clb grid_clb_11__9_ (
    .prog_clk ( { ctsbuf_net_1632145 } ) ,
    .Test_en ( { BUF_net_854 } ) ,
    .clk ( { ctsbuf_net_171999 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_118_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_261_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__128_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__128_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__128_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__128_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__128_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__128_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__128_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__128_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__128_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__128_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__128_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__128_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__128_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__128_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__128_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__128_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__117_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__117_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__117_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__117_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__117_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__117_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__117_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__117_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__117_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__117_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__117_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__117_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__117_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__117_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__117_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__117_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__116_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__116_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_128_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_128_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_128_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_128_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_128_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_128_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_128_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_128_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_128_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_128_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_128_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_128_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_128_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_128_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_128_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_128_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_128_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_128_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_128_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_128_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_128_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_128_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_128_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_128_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_128_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_128_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_128_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_128_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_128_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_128_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_128_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_128_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_128_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_128_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_128_ccff_tail ) ) ;
grid_clb grid_clb_11__10_ (
    .prog_clk ( { ctsbuf_net_1282110 } ) ,
    .Test_en ( { BUF_net_731 } ) ,
    .clk ( { ctsbuf_net_171999 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_119_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_262_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__129_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__129_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__129_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__129_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__129_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__129_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__129_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__129_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__129_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__129_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__129_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__129_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__129_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__129_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__129_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__129_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__118_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__118_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__118_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__118_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__118_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__118_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__118_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__118_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__118_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__118_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__118_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__118_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__118_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__118_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__118_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__118_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__117_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__117_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_129_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_129_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_129_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_129_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_129_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_129_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_129_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_129_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_129_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_129_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_129_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_129_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_129_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_129_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_129_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_129_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_129_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_129_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_129_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_129_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_129_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_129_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_129_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_129_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_129_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_129_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_129_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_129_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_129_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_129_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_129_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_129_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_129_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_129_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_129_ccff_tail ) ) ;
grid_clb grid_clb_11__11_ (
    .prog_clk ( { ctsbuf_net_992081 } ) ,
    .Test_en ( { BUF_net_858 } ) ,
    .clk ( { ctsbuf_net_242006 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_120_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_263_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__130_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__130_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__130_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__130_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__130_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__130_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__130_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__130_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__130_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__130_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__130_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__130_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__130_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__130_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__130_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__130_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__119_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__119_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__119_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__119_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__119_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__119_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__119_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__119_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__119_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__119_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__119_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__119_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__119_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__119_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__119_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__119_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__118_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__118_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_130_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_130_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_130_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_130_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_130_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_130_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_130_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_130_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_130_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_130_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_130_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_130_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_130_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_130_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_130_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_130_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_130_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_130_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_130_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_130_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_130_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_130_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_130_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_130_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_130_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_130_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_130_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_130_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_130_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_130_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_130_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_130_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_130_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_130_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_130_ccff_tail ) ) ;
grid_clb grid_clb_11__12_ (
    .prog_clk ( { p_abuf0 } ) ,
    .Test_en ( { BUF_net_452 } ) ,
    .clk ( { ctsbuf_net_242006 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_141_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_284_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__131_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__131_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__131_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__131_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__131_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__131_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__131_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__131_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__131_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__131_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__131_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__131_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__131_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__131_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__131_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__131_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__120_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__120_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__120_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__120_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__120_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__120_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__120_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__120_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__120_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__120_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__120_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__120_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__120_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__120_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__120_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__120_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__119_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__119_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_131_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_131_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_131_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_131_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_131_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_131_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_131_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_131_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_131_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_131_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_131_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_131_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_131_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_131_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_131_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_131_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_131_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_131_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_131_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_131_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_131_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_131_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_131_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_131_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_131_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_131_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_131_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_131_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_131_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_131_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_131_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_131_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_131_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_131_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_131_ccff_tail ) ) ;
grid_clb grid_clb_12__1_ (
    .prog_clk ( { ctsbuf_net_492031 } ) ,
    .Test_en ( { BUF_net_451 } ) ,
    .clk ( { ctsbuf_net_11983 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_121_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_264_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__132_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__132_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__132_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__132_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__132_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__132_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__132_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__132_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__132_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__132_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__132_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__132_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__132_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__132_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__132_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__132_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__0__11_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__0__11_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__0__11_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__0__11_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__0__11_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__0__11_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__0__11_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__0__11_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__0__11_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__0__11_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__0__11_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__0__11_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__0__11_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__0__11_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__0__11_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__0__11_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__120_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__120_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_132_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_132_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_132_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_132_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_132_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_132_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_132_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_132_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_132_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_132_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_132_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_132_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_132_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_132_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_132_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_132_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_132_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_132_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_132_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_132_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_132_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_132_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_132_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_132_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_132_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_132_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_132_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_132_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_132_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_132_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_132_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_132_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_12__1__undriven_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_12__1__undriven_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_132_ccff_tail ) ) ;
grid_clb grid_clb_12__2_ (
    .prog_clk ( { ctsbuf_net_622044 } ) ,
    .Test_en ( { BUF_net_450 } ) ,
    .clk ( { ctsbuf_net_11983 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_122_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_265_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__133_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__133_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__133_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__133_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__133_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__133_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__133_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__133_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__133_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__133_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__133_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__133_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__133_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__133_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__133_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__133_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__121_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__121_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__121_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__121_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__121_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__121_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__121_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__121_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__121_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__121_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__121_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__121_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__121_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__121_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__121_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__121_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__121_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__121_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_133_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_133_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_133_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_133_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_133_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_133_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_133_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_133_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_133_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_133_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_133_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_133_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_133_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_133_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_133_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_133_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_133_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_133_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_133_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_133_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_133_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_133_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_133_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_133_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_133_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_133_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_133_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_133_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_133_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_133_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_133_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_133_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_133_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_133_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_133_ccff_tail ) ) ;
grid_clb grid_clb_12__3_ (
    .prog_clk ( { ctsbuf_net_822064 } ) ,
    .Test_en ( { BUF_net_449 } ) ,
    .clk ( { ctsbuf_net_41986 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_123_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_266_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__134_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__134_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__134_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__134_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__134_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__134_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__134_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__134_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__134_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__134_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__134_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__134_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__134_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__134_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__134_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__134_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__122_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__122_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__122_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__122_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__122_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__122_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__122_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__122_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__122_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__122_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__122_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__122_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__122_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__122_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__122_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__122_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__122_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__122_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_134_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_134_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_134_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_134_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_134_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_134_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_134_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_134_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_134_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_134_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_134_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_134_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_134_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_134_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_134_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_134_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_134_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_134_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_134_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_134_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_134_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_134_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_134_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_134_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_134_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_134_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_134_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_134_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_134_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_134_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_134_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_134_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_134_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_134_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_134_ccff_tail ) ) ;
grid_clb grid_clb_12__4_ (
    .prog_clk ( { ctsbuf_net_1102092 } ) ,
    .Test_en ( { BUF_net_448 } ) ,
    .clk ( { ctsbuf_net_41986 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_124_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_267_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__135_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__135_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__135_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__135_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__135_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__135_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__135_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__135_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__135_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__135_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__135_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__135_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__135_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__135_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__135_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__135_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__123_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__123_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__123_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__123_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__123_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__123_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__123_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__123_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__123_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__123_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__123_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__123_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__123_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__123_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__123_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__123_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__123_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__123_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_135_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_135_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_135_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_135_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_135_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_135_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_135_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_135_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_135_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_135_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_135_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_135_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_135_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_135_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_135_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_135_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_135_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_135_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_135_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_135_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_135_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_135_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_135_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_135_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_135_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_135_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_135_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_135_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_135_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_135_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_135_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_135_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_135_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_135_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_135_ccff_tail ) ) ;
grid_clb grid_clb_12__5_ (
    .prog_clk ( { ctsbuf_net_1422124 } ) ,
    .Test_en ( { BUF_net_447 } ) ,
    .clk ( { ctsbuf_net_91991 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_125_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_268_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__136_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__136_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__136_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__136_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__136_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__136_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__136_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__136_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__136_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__136_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__136_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__136_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__136_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__136_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__136_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__136_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__124_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__124_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__124_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__124_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__124_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__124_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__124_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__124_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__124_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__124_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__124_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__124_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__124_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__124_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__124_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__124_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__124_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__124_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_136_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_136_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_136_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_136_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_136_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_136_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_136_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_136_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_136_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_136_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_136_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_136_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_136_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_136_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_136_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_136_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_136_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_136_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_136_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_136_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_136_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_136_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_136_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_136_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_136_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_136_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_136_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_136_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_136_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_136_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_136_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_136_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_136_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_136_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_136_ccff_tail ) ) ;
grid_clb grid_clb_12__6_ (
    .prog_clk ( { ctsbuf_net_1822164 } ) ,
    .Test_en ( { BUF_net_446 } ) ,
    .clk ( { ctsbuf_net_91991 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_126_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_269_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__137_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__137_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__137_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__137_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__137_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__137_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__137_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__137_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__137_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__137_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__137_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__137_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__137_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__137_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__137_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__137_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__125_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__125_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__125_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__125_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__125_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__125_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__125_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__125_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__125_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__125_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__125_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__125_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__125_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__125_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__125_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__125_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__125_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__125_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_137_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_137_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_137_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_137_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_137_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_137_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_137_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_137_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_137_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_137_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_137_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_137_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_137_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_137_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_137_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_137_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_137_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_137_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_137_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_137_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_137_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_137_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_137_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_137_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_137_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_137_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_137_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_137_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_137_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_137_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_137_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_137_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_137_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_137_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_137_ccff_tail ) ) ;
grid_clb grid_clb_12__7_ (
    .prog_clk ( { ctsbuf_net_2082190 } ) ,
    .Test_en ( { BUF_net_445 } ) ,
    .clk ( { ctsbuf_net_141996 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_127_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_270_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__138_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__138_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__138_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__138_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__138_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__138_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__138_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__138_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__138_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__138_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__138_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__138_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__138_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__138_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__138_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__138_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__126_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__126_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__126_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__126_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__126_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__126_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__126_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__126_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__126_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__126_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__126_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__126_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__126_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__126_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__126_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__126_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__126_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__126_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_138_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_138_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_138_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_138_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_138_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_138_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_138_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_138_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_138_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_138_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_138_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_138_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_138_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_138_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_138_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_138_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_138_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_138_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_138_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_138_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_138_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_138_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_138_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_138_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_138_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_138_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_138_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_138_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_138_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_138_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_138_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_138_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_138_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_138_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_138_ccff_tail ) ) ;
grid_clb grid_clb_12__8_ (
    .prog_clk ( { ctsbuf_net_1652147 } ) ,
    .Test_en ( { BUF_net_444 } ) ,
    .clk ( { ctsbuf_net_141996 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_128_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_271_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__139_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__139_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__139_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__139_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__139_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__139_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__139_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__139_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__139_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__139_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__139_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__139_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__139_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__139_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__139_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__139_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__127_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__127_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__127_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__127_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__127_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__127_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__127_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__127_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__127_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__127_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__127_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__127_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__127_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__127_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__127_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__127_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__127_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__127_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_139_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_139_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_139_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_139_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_139_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_139_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_139_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_139_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_139_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_139_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_139_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_139_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_139_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_139_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_139_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_139_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_139_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_139_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_139_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_139_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_139_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_139_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_139_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_139_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_139_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_139_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_139_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_139_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_139_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_139_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_139_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_139_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_139_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_139_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_139_ccff_tail ) ) ;
grid_clb grid_clb_12__9_ (
    .prog_clk ( { ctsbuf_net_1292111 } ) ,
    .Test_en ( { BUF_net_443 } ) ,
    .clk ( { ctsbuf_net_171999 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_129_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_272_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__140_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__140_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__140_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__140_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__140_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__140_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__140_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__140_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__140_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__140_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__140_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__140_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__140_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__140_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__140_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__140_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__128_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__128_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__128_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__128_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__128_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__128_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__128_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__128_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__128_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__128_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__128_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__128_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__128_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__128_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__128_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__128_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__128_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__128_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_140_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_140_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_140_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_140_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_140_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_140_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_140_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_140_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_140_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_140_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_140_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_140_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_140_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_140_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_140_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_140_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_140_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_140_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_140_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_140_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_140_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_140_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_140_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_140_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_140_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_140_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_140_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_140_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_140_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_140_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_140_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_140_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_140_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_140_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_140_ccff_tail ) ) ;
grid_clb grid_clb_12__10_ (
    .prog_clk ( { ctsbuf_net_1012083 } ) ,
    .Test_en ( { BUF_net_442 } ) ,
    .clk ( { ctsbuf_net_171999 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_130_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_273_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__141_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__141_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__141_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__141_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__141_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__141_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__141_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__141_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__141_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__141_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__141_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__141_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__141_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__141_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__141_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__141_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__129_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__129_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__129_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__129_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__129_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__129_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__129_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__129_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__129_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__129_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__129_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__129_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__129_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__129_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__129_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__129_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__129_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__129_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_141_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_141_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_141_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_141_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_141_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_141_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_141_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_141_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_141_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_141_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_141_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_141_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_141_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_141_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_141_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_141_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_141_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_141_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_141_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_141_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_141_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_141_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_141_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_141_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_141_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_141_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_141_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_141_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_141_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_141_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_141_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_141_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_141_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_141_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_141_ccff_tail ) ) ;
grid_clb grid_clb_12__11_ (
    .prog_clk ( { ctsbuf_net_742056 } ) ,
    .Test_en ( { BUF_net_441 } ) ,
    .clk ( { ctsbuf_net_242006 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_131_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_274_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__142_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__142_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__142_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__142_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__142_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__142_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__142_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__142_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__142_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__142_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__142_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__142_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__142_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__142_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__142_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__142_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__130_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__130_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__130_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__130_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__130_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__130_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__130_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__130_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__130_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__130_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__130_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__130_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__130_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__130_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__130_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__130_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__130_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__130_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_142_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_142_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_142_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_142_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_142_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_142_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_142_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_142_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_142_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_142_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_142_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_142_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_142_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_142_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_142_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_142_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_142_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_142_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_142_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_142_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_142_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_142_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_142_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_142_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_142_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_142_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_142_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_142_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_142_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_142_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_142_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_142_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_142_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_142_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_142_ccff_tail ) ) ;
grid_clb grid_clb_12__12_ (
    .prog_clk ( { ctsbuf_net_562038 } ) ,
    .Test_en ( { BUF_net_440 } ) ,
    .clk ( { ctsbuf_net_242006 } ) ,
    .top_width_0_height_0__pin_32_ ( direct_interc_142_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_285_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__143_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__143_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__143_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__143_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__143_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__143_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__143_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__143_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__143_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__143_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__143_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__143_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__143_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__143_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__143_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__143_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__131_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__131_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__131_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__131_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__131_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__131_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__131_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__131_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__131_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__131_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__131_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__131_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__131_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__131_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__131_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__131_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__131_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__131_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_143_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_143_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_143_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_143_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_143_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_143_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_143_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_143_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_143_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_143_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_143_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_143_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_143_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_143_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_143_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_143_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_143_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_143_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_143_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_143_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_143_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_143_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_143_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_143_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_143_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_143_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_143_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_143_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_143_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_143_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_143_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_143_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_143_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_143_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_143_ccff_tail ) ) ;
grid_io_top grid_io_top_1__13_ (
    .prog_clk ( { ctsbuf_net_4162398 } ) ,
    .gfpga_pad_GPIO_A ( gfpga_pad_GPIO_A[0] ) , 
    .gfpga_pad_GPIO_IE ( gfpga_pad_GPIO_IE[0] ) , 
    .gfpga_pad_GPIO_OE ( gfpga_pad_GPIO_OE[0] ) , 
    .gfpga_pad_GPIO_Y ( gfpga_pad_GPIO_Y[0] ) , 
    .bottom_width_0_height_0__pin_0_ ( cbx_1__12__0_top_grid_pin_0_ ) , 
    .ccff_head ( cbx_1__12__0_ccff_tail ) , 
    .bottom_width_0_height_0__pin_1_upper ( grid_io_top_0_bottom_width_0_height_0__pin_1_upper ) , 
    .bottom_width_0_height_0__pin_1_lower ( grid_io_top_0_bottom_width_0_height_0__pin_1_lower ) , 
    .ccff_tail ( grid_io_top_0_ccff_tail ) ) ;
grid_io_top grid_io_top_2__13_ (
    .prog_clk ( { ctsbuf_net_3292311 } ) ,
    .gfpga_pad_GPIO_A ( gfpga_pad_GPIO_A[1] ) , 
    .gfpga_pad_GPIO_IE ( gfpga_pad_GPIO_IE[1] ) , 
    .gfpga_pad_GPIO_OE ( gfpga_pad_GPIO_OE[1] ) , 
    .gfpga_pad_GPIO_Y ( gfpga_pad_GPIO_Y[1] ) , 
    .bottom_width_0_height_0__pin_0_ ( cbx_1__12__1_top_grid_pin_0_ ) , 
    .ccff_head ( cbx_1__12__1_ccff_tail ) , 
    .bottom_width_0_height_0__pin_1_upper ( grid_io_top_1_bottom_width_0_height_0__pin_1_upper ) , 
    .bottom_width_0_height_0__pin_1_lower ( grid_io_top_1_bottom_width_0_height_0__pin_1_lower ) , 
    .ccff_tail ( grid_io_top_1_ccff_tail ) ) ;
grid_io_top grid_io_top_3__13_ (
    .prog_clk ( { ctsbuf_net_3292311 } ) ,
    .gfpga_pad_GPIO_A ( gfpga_pad_GPIO_A[2] ) , 
    .gfpga_pad_GPIO_IE ( gfpga_pad_GPIO_IE[2] ) , 
    .gfpga_pad_GPIO_OE ( gfpga_pad_GPIO_OE[2] ) , 
    .gfpga_pad_GPIO_Y ( gfpga_pad_GPIO_Y[2] ) , 
    .bottom_width_0_height_0__pin_0_ ( cbx_1__12__2_top_grid_pin_0_ ) , 
    .ccff_head ( cbx_1__12__2_ccff_tail ) , 
    .bottom_width_0_height_0__pin_1_upper ( grid_io_top_2_bottom_width_0_height_0__pin_1_upper ) , 
    .bottom_width_0_height_0__pin_1_lower ( grid_io_top_2_bottom_width_0_height_0__pin_1_lower ) , 
    .ccff_tail ( grid_io_top_2_ccff_tail ) ) ;
grid_io_top grid_io_top_4__13_ (
    .prog_clk ( { ctsbuf_net_2392221 } ) ,
    .gfpga_pad_GPIO_A ( gfpga_pad_GPIO_A[3] ) , 
    .gfpga_pad_GPIO_IE ( gfpga_pad_GPIO_IE[3] ) , 
    .gfpga_pad_GPIO_OE ( gfpga_pad_GPIO_OE[3] ) , 
    .gfpga_pad_GPIO_Y ( gfpga_pad_GPIO_Y[3] ) , 
    .bottom_width_0_height_0__pin_0_ ( cbx_1__12__3_top_grid_pin_0_ ) , 
    .ccff_head ( cbx_1__12__3_ccff_tail ) , 
    .bottom_width_0_height_0__pin_1_upper ( grid_io_top_3_bottom_width_0_height_0__pin_1_upper ) , 
    .bottom_width_0_height_0__pin_1_lower ( grid_io_top_3_bottom_width_0_height_0__pin_1_lower ) , 
    .ccff_tail ( grid_io_top_3_ccff_tail ) ) ;
grid_io_top grid_io_top_5__13_ (
    .prog_clk ( { ctsbuf_net_2392221 } ) ,
    .gfpga_pad_GPIO_A ( gfpga_pad_GPIO_A[4] ) , 
    .gfpga_pad_GPIO_IE ( gfpga_pad_GPIO_IE[4] ) , 
    .gfpga_pad_GPIO_OE ( gfpga_pad_GPIO_OE[4] ) , 
    .gfpga_pad_GPIO_Y ( gfpga_pad_GPIO_Y[4] ) , 
    .bottom_width_0_height_0__pin_0_ ( cbx_1__12__4_top_grid_pin_0_ ) , 
    .ccff_head ( cbx_1__12__4_ccff_tail ) , 
    .bottom_width_0_height_0__pin_1_upper ( grid_io_top_4_bottom_width_0_height_0__pin_1_upper ) , 
    .bottom_width_0_height_0__pin_1_lower ( grid_io_top_4_bottom_width_0_height_0__pin_1_lower ) , 
    .ccff_tail ( grid_io_top_4_ccff_tail ) ) ;
grid_io_top grid_io_top_6__13_ (
    .prog_clk ( { ctsbuf_net_1532135 } ) ,
    .gfpga_pad_GPIO_A ( gfpga_pad_GPIO_A[5] ) , 
    .gfpga_pad_GPIO_IE ( gfpga_pad_GPIO_IE[5] ) , 
    .gfpga_pad_GPIO_OE ( gfpga_pad_GPIO_OE[5] ) , 
    .gfpga_pad_GPIO_Y ( gfpga_pad_GPIO_Y[5] ) , 
    .bottom_width_0_height_0__pin_0_ ( cbx_1__12__5_top_grid_pin_0_ ) , 
    .ccff_head ( cbx_1__12__5_ccff_tail ) , 
    .bottom_width_0_height_0__pin_1_upper ( grid_io_top_5_bottom_width_0_height_0__pin_1_upper ) , 
    .bottom_width_0_height_0__pin_1_lower ( grid_io_top_5_bottom_width_0_height_0__pin_1_lower ) , 
    .ccff_tail ( grid_io_top_5_ccff_tail ) ) ;
grid_io_top grid_io_top_7__13_ (
    .prog_clk ( { ctsbuf_net_1532135 } ) ,
    .gfpga_pad_GPIO_A ( gfpga_pad_GPIO_A[6] ) , 
    .gfpga_pad_GPIO_IE ( gfpga_pad_GPIO_IE[6] ) , 
    .gfpga_pad_GPIO_OE ( gfpga_pad_GPIO_OE[6] ) , 
    .gfpga_pad_GPIO_Y ( gfpga_pad_GPIO_Y[6] ) , 
    .bottom_width_0_height_0__pin_0_ ( cbx_1__12__6_top_grid_pin_0_ ) , 
    .ccff_head ( cbx_1__12__6_ccff_tail ) , 
    .bottom_width_0_height_0__pin_1_upper ( grid_io_top_6_bottom_width_0_height_0__pin_1_upper ) , 
    .bottom_width_0_height_0__pin_1_lower ( grid_io_top_6_bottom_width_0_height_0__pin_1_lower ) , 
    .ccff_tail ( grid_io_top_6_ccff_tail ) ) ;
grid_io_top grid_io_top_8__13_ (
    .prog_clk ( { p_abuf3 } ) ,
    .gfpga_pad_GPIO_A ( gfpga_pad_GPIO_A[7] ) , 
    .gfpga_pad_GPIO_IE ( gfpga_pad_GPIO_IE[7] ) , 
    .gfpga_pad_GPIO_OE ( gfpga_pad_GPIO_OE[7] ) , 
    .gfpga_pad_GPIO_Y ( gfpga_pad_GPIO_Y[7] ) , 
    .bottom_width_0_height_0__pin_0_ ( cbx_1__12__7_top_grid_pin_0_ ) , 
    .ccff_head ( cbx_1__12__7_ccff_tail ) , 
    .bottom_width_0_height_0__pin_1_upper ( grid_io_top_7_bottom_width_0_height_0__pin_1_upper ) , 
    .bottom_width_0_height_0__pin_1_lower ( grid_io_top_7_bottom_width_0_height_0__pin_1_lower ) , 
    .ccff_tail ( grid_io_top_7_ccff_tail ) ) ;
grid_io_top grid_io_top_9__13_ (
    .prog_clk ( { p_abuf4 } ) ,
    .gfpga_pad_GPIO_A ( gfpga_pad_GPIO_A[8] ) , 
    .gfpga_pad_GPIO_IE ( gfpga_pad_GPIO_IE[8] ) , 
    .gfpga_pad_GPIO_OE ( gfpga_pad_GPIO_OE[8] ) , 
    .gfpga_pad_GPIO_Y ( gfpga_pad_GPIO_Y[8] ) , 
    .bottom_width_0_height_0__pin_0_ ( cbx_1__12__8_top_grid_pin_0_ ) , 
    .ccff_head ( cbx_1__12__8_ccff_tail ) , 
    .bottom_width_0_height_0__pin_1_upper ( grid_io_top_8_bottom_width_0_height_0__pin_1_upper ) , 
    .bottom_width_0_height_0__pin_1_lower ( grid_io_top_8_bottom_width_0_height_0__pin_1_lower ) , 
    .ccff_tail ( grid_io_top_8_ccff_tail ) ) ;
grid_io_top grid_io_top_10__13_ (
    .prog_clk ( { ctsbuf_net_532035 } ) ,
    .gfpga_pad_GPIO_A ( gfpga_pad_GPIO_A[9] ) , 
    .gfpga_pad_GPIO_IE ( gfpga_pad_GPIO_IE[9] ) , 
    .gfpga_pad_GPIO_OE ( gfpga_pad_GPIO_OE[9] ) , 
    .gfpga_pad_GPIO_Y ( gfpga_pad_GPIO_Y[9] ) , 
    .bottom_width_0_height_0__pin_0_ ( cbx_1__12__9_top_grid_pin_0_ ) , 
    .ccff_head ( cbx_1__12__9_ccff_tail ) , 
    .bottom_width_0_height_0__pin_1_upper ( grid_io_top_9_bottom_width_0_height_0__pin_1_upper ) , 
    .bottom_width_0_height_0__pin_1_lower ( grid_io_top_9_bottom_width_0_height_0__pin_1_lower ) , 
    .ccff_tail ( grid_io_top_9_ccff_tail ) ) ;
grid_io_top grid_io_top_11__13_ (
    .prog_clk ( { ctsbuf_net_532035 } ) ,
    .gfpga_pad_GPIO_A ( gfpga_pad_GPIO_A[10] ) , 
    .gfpga_pad_GPIO_IE ( gfpga_pad_GPIO_IE[10] ) , 
    .gfpga_pad_GPIO_OE ( gfpga_pad_GPIO_OE[10] ) , 
    .gfpga_pad_GPIO_Y ( gfpga_pad_GPIO_Y[10] ) , 
    .bottom_width_0_height_0__pin_0_ ( cbx_1__12__10_top_grid_pin_0_ ) , 
    .ccff_head ( cbx_1__12__10_ccff_tail ) , 
    .bottom_width_0_height_0__pin_1_upper ( grid_io_top_10_bottom_width_0_height_0__pin_1_upper ) , 
    .bottom_width_0_height_0__pin_1_lower ( grid_io_top_10_bottom_width_0_height_0__pin_1_lower ) , 
    .ccff_tail ( grid_io_top_10_ccff_tail ) ) ;
grid_io_top grid_io_top_12__13_ (
    .prog_clk ( { ctsbuf_net_462028 } ) ,
    .gfpga_pad_GPIO_A ( gfpga_pad_GPIO_A[11] ) , 
    .gfpga_pad_GPIO_IE ( gfpga_pad_GPIO_IE[11] ) , 
    .gfpga_pad_GPIO_OE ( gfpga_pad_GPIO_OE[11] ) , 
    .gfpga_pad_GPIO_Y ( gfpga_pad_GPIO_Y[11] ) , 
    .bottom_width_0_height_0__pin_0_ ( cbx_1__12__11_top_grid_pin_0_ ) , 
    .ccff_head ( cbx_1__12__11_ccff_tail ) , 
    .bottom_width_0_height_0__pin_1_upper ( grid_io_top_11_bottom_width_0_height_0__pin_1_upper ) , 
    .bottom_width_0_height_0__pin_1_lower ( grid_io_top_11_bottom_width_0_height_0__pin_1_lower ) , 
    .ccff_tail ( grid_io_top_11_ccff_tail ) ) ;
grid_io_right grid_io_right_13__1_ (
    .prog_clk ( { ctsbuf_net_452027 } ) ,
    .gfpga_pad_GPIO_A ( gfpga_pad_GPIO_A[12] ) , 
    .gfpga_pad_GPIO_IE ( gfpga_pad_GPIO_IE[12] ) , 
    .gfpga_pad_GPIO_OE ( gfpga_pad_GPIO_OE[12] ) , 
    .gfpga_pad_GPIO_Y ( gfpga_pad_GPIO_Y[12] ) , 
    .left_width_0_height_0__pin_0_ ( cby_1__1__132_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__132_ccff_tail ) , 
    .left_width_0_height_0__pin_1_upper ( grid_io_right_0_left_width_0_height_0__pin_1_upper ) , 
    .left_width_0_height_0__pin_1_lower ( grid_io_right_0_left_width_0_height_0__pin_1_lower ) , 
    .ccff_tail ( grid_io_right_0_ccff_tail ) ) ;
grid_io_right grid_io_right_13__2_ (
    .prog_clk ( { ctsbuf_net_502032 } ) ,
    .gfpga_pad_GPIO_A ( gfpga_pad_GPIO_A[13] ) , 
    .gfpga_pad_GPIO_IE ( gfpga_pad_GPIO_IE[13] ) , 
    .gfpga_pad_GPIO_OE ( gfpga_pad_GPIO_OE[13] ) , 
    .gfpga_pad_GPIO_Y ( gfpga_pad_GPIO_Y[13] ) , 
    .left_width_0_height_0__pin_0_ ( cby_1__1__133_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__133_ccff_tail ) , 
    .left_width_0_height_0__pin_1_upper ( grid_io_right_1_left_width_0_height_0__pin_1_upper ) , 
    .left_width_0_height_0__pin_1_lower ( grid_io_right_1_left_width_0_height_0__pin_1_lower ) , 
    .ccff_tail ( grid_io_right_1_ccff_tail ) ) ;
grid_io_right grid_io_right_13__3_ (
    .prog_clk ( { ctsbuf_net_632045 } ) ,
    .gfpga_pad_GPIO_A ( gfpga_pad_GPIO_A[14] ) , 
    .gfpga_pad_GPIO_IE ( gfpga_pad_GPIO_IE[14] ) , 
    .gfpga_pad_GPIO_OE ( gfpga_pad_GPIO_OE[14] ) , 
    .gfpga_pad_GPIO_Y ( gfpga_pad_GPIO_Y[14] ) , 
    .left_width_0_height_0__pin_0_ ( cby_1__1__134_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__134_ccff_tail ) , 
    .left_width_0_height_0__pin_1_upper ( grid_io_right_2_left_width_0_height_0__pin_1_upper ) , 
    .left_width_0_height_0__pin_1_lower ( grid_io_right_2_left_width_0_height_0__pin_1_lower ) , 
    .ccff_tail ( grid_io_right_2_ccff_tail ) ) ;
grid_io_right grid_io_right_13__4_ (
    .prog_clk ( { ctsbuf_net_832065 } ) ,
    .gfpga_pad_GPIO_A ( gfpga_pad_GPIO_A[15] ) , 
    .gfpga_pad_GPIO_IE ( gfpga_pad_GPIO_IE[15] ) , 
    .gfpga_pad_GPIO_OE ( gfpga_pad_GPIO_OE[15] ) , 
    .gfpga_pad_GPIO_Y ( gfpga_pad_GPIO_Y[15] ) , 
    .left_width_0_height_0__pin_0_ ( cby_1__1__135_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__135_ccff_tail ) , 
    .left_width_0_height_0__pin_1_upper ( grid_io_right_3_left_width_0_height_0__pin_1_upper ) , 
    .left_width_0_height_0__pin_1_lower ( grid_io_right_3_left_width_0_height_0__pin_1_lower ) , 
    .ccff_tail ( grid_io_right_3_ccff_tail ) ) ;
grid_io_right grid_io_right_13__5_ (
    .prog_clk ( { ctsbuf_net_1112093 } ) ,
    .gfpga_pad_GPIO_A ( gfpga_pad_GPIO_A[16] ) , 
    .gfpga_pad_GPIO_IE ( gfpga_pad_GPIO_IE[16] ) , 
    .gfpga_pad_GPIO_OE ( gfpga_pad_GPIO_OE[16] ) , 
    .gfpga_pad_GPIO_Y ( gfpga_pad_GPIO_Y[16] ) , 
    .left_width_0_height_0__pin_0_ ( cby_1__1__136_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__136_ccff_tail ) , 
    .left_width_0_height_0__pin_1_upper ( grid_io_right_4_left_width_0_height_0__pin_1_upper ) , 
    .left_width_0_height_0__pin_1_lower ( grid_io_right_4_left_width_0_height_0__pin_1_lower ) , 
    .ccff_tail ( grid_io_right_4_ccff_tail ) ) ;
grid_io_right grid_io_right_13__6_ (
    .prog_clk ( { ctsbuf_net_1432125 } ) ,
    .gfpga_pad_GPIO_A ( gfpga_pad_GPIO_A[17] ) , 
    .gfpga_pad_GPIO_IE ( gfpga_pad_GPIO_IE[17] ) , 
    .gfpga_pad_GPIO_OE ( gfpga_pad_GPIO_OE[17] ) , 
    .gfpga_pad_GPIO_Y ( gfpga_pad_GPIO_Y[17] ) , 
    .left_width_0_height_0__pin_0_ ( cby_1__1__137_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__137_ccff_tail ) , 
    .left_width_0_height_0__pin_1_upper ( grid_io_right_5_left_width_0_height_0__pin_1_upper ) , 
    .left_width_0_height_0__pin_1_lower ( grid_io_right_5_left_width_0_height_0__pin_1_lower ) , 
    .ccff_tail ( grid_io_right_5_ccff_tail ) ) ;
grid_io_right grid_io_right_13__7_ (
    .prog_clk ( { ctsbuf_net_1202102 } ) ,
    .gfpga_pad_GPIO_A ( gfpga_pad_GPIO_A[18] ) , 
    .gfpga_pad_GPIO_IE ( gfpga_pad_GPIO_IE[18] ) , 
    .gfpga_pad_GPIO_OE ( gfpga_pad_GPIO_OE[18] ) , 
    .gfpga_pad_GPIO_Y ( gfpga_pad_GPIO_Y[18] ) , 
    .left_width_0_height_0__pin_0_ ( cby_1__1__138_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__138_ccff_tail ) , 
    .left_width_0_height_0__pin_1_upper ( grid_io_right_6_left_width_0_height_0__pin_1_upper ) , 
    .left_width_0_height_0__pin_1_lower ( grid_io_right_6_left_width_0_height_0__pin_1_lower ) , 
    .ccff_tail ( grid_io_right_6_ccff_tail ) ) ;
grid_io_right grid_io_right_13__8_ (
    .prog_clk ( { ctsbuf_net_1202102 } ) ,
    .gfpga_pad_GPIO_A ( gfpga_pad_GPIO_A[19] ) , 
    .gfpga_pad_GPIO_IE ( gfpga_pad_GPIO_IE[19] ) , 
    .gfpga_pad_GPIO_OE ( gfpga_pad_GPIO_OE[19] ) , 
    .gfpga_pad_GPIO_Y ( gfpga_pad_GPIO_Y[19] ) , 
    .left_width_0_height_0__pin_0_ ( cby_1__1__139_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__139_ccff_tail ) , 
    .left_width_0_height_0__pin_1_upper ( grid_io_right_7_left_width_0_height_0__pin_1_upper ) , 
    .left_width_0_height_0__pin_1_lower ( grid_io_right_7_left_width_0_height_0__pin_1_lower ) , 
    .ccff_tail ( grid_io_right_7_ccff_tail ) ) ;
grid_io_right grid_io_right_13__9_ (
    .prog_clk ( { ctsbuf_net_912073 } ) ,
    .gfpga_pad_GPIO_A ( gfpga_pad_GPIO_A[20] ) , 
    .gfpga_pad_GPIO_IE ( gfpga_pad_GPIO_IE[20] ) , 
    .gfpga_pad_GPIO_OE ( gfpga_pad_GPIO_OE[20] ) , 
    .gfpga_pad_GPIO_Y ( gfpga_pad_GPIO_Y[20] ) , 
    .left_width_0_height_0__pin_0_ ( cby_1__1__140_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__140_ccff_tail ) , 
    .left_width_0_height_0__pin_1_upper ( grid_io_right_8_left_width_0_height_0__pin_1_upper ) , 
    .left_width_0_height_0__pin_1_lower ( grid_io_right_8_left_width_0_height_0__pin_1_lower ) , 
    .ccff_tail ( grid_io_right_8_ccff_tail ) ) ;
grid_io_right grid_io_right_13__10_ (
    .prog_clk ( { ctsbuf_net_682050 } ) ,
    .gfpga_pad_GPIO_A ( gfpga_pad_GPIO_A[21] ) , 
    .gfpga_pad_GPIO_IE ( gfpga_pad_GPIO_IE[21] ) , 
    .gfpga_pad_GPIO_OE ( gfpga_pad_GPIO_OE[21] ) , 
    .gfpga_pad_GPIO_Y ( gfpga_pad_GPIO_Y[21] ) , 
    .left_width_0_height_0__pin_0_ ( cby_1__1__141_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__141_ccff_tail ) , 
    .left_width_0_height_0__pin_1_upper ( grid_io_right_9_left_width_0_height_0__pin_1_upper ) , 
    .left_width_0_height_0__pin_1_lower ( grid_io_right_9_left_width_0_height_0__pin_1_lower ) , 
    .ccff_tail ( grid_io_right_9_ccff_tail ) ) ;
grid_io_right grid_io_right_13__11_ (
    .prog_clk ( { ctsbuf_net_472029 } ) ,
    .gfpga_pad_GPIO_A ( gfpga_pad_GPIO_A[22] ) , 
    .gfpga_pad_GPIO_IE ( gfpga_pad_GPIO_IE[22] ) , 
    .gfpga_pad_GPIO_OE ( gfpga_pad_GPIO_OE[22] ) , 
    .gfpga_pad_GPIO_Y ( gfpga_pad_GPIO_Y[22] ) , 
    .left_width_0_height_0__pin_0_ ( cby_1__1__142_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__142_ccff_tail ) , 
    .left_width_0_height_0__pin_1_upper ( grid_io_right_10_left_width_0_height_0__pin_1_upper ) , 
    .left_width_0_height_0__pin_1_lower ( grid_io_right_10_left_width_0_height_0__pin_1_lower ) , 
    .ccff_tail ( grid_io_right_10_ccff_tail ) ) ;
grid_io_right grid_io_right_13__12_ (
    .prog_clk ( { ctsbuf_net_472029 } ) ,
    .gfpga_pad_GPIO_A ( gfpga_pad_GPIO_A[23] ) , 
    .gfpga_pad_GPIO_IE ( gfpga_pad_GPIO_IE[23] ) , 
    .gfpga_pad_GPIO_OE ( gfpga_pad_GPIO_OE[23] ) , 
    .gfpga_pad_GPIO_Y ( gfpga_pad_GPIO_Y[23] ) , 
    .left_width_0_height_0__pin_0_ ( cby_1__1__143_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__143_ccff_tail ) , 
    .left_width_0_height_0__pin_1_upper ( grid_io_right_11_left_width_0_height_0__pin_1_upper ) , 
    .left_width_0_height_0__pin_1_lower ( grid_io_right_11_left_width_0_height_0__pin_1_lower ) , 
    .ccff_tail ( grid_io_right_11_ccff_tail ) ) ;
grid_io_bottom grid_io_bottom_1__0_ (
    .prog_clk ( { ctsbuf_net_4172399 } ) ,
    .gfpga_pad_GPIO_A ( gfpga_pad_GPIO_A[24] ) , 
    .gfpga_pad_GPIO_IE ( gfpga_pad_GPIO_IE[24] ) , 
    .gfpga_pad_GPIO_OE ( gfpga_pad_GPIO_OE[24] ) , 
    .gfpga_pad_GPIO_Y ( gfpga_pad_GPIO_Y[24] ) , 
    .top_width_0_height_0__pin_0_ ( cbx_1__0__0_bottom_grid_pin_0_ ) , 
    .ccff_head ( cbx_1__0__0_ccff_tail ) , 
    .top_width_0_height_0__pin_1_upper ( grid_io_bottom_0_top_width_0_height_0__pin_1_upper ) , 
    .top_width_0_height_0__pin_1_lower ( grid_io_bottom_0_top_width_0_height_0__pin_1_lower ) , 
    .ccff_tail ( grid_io_bottom_0_ccff_tail ) ) ;
grid_io_bottom grid_io_bottom_2__0_ (
    .prog_clk ( { ctsbuf_net_3732355 } ) ,
    .gfpga_pad_GPIO_A ( gfpga_pad_GPIO_A[25] ) , 
    .gfpga_pad_GPIO_IE ( gfpga_pad_GPIO_IE[25] ) , 
    .gfpga_pad_GPIO_OE ( gfpga_pad_GPIO_OE[25] ) , 
    .gfpga_pad_GPIO_Y ( gfpga_pad_GPIO_Y[25] ) , 
    .top_width_0_height_0__pin_0_ ( cbx_1__0__1_bottom_grid_pin_0_ ) , 
    .ccff_head ( cbx_1__0__1_ccff_tail ) , 
    .top_width_0_height_0__pin_1_upper ( grid_io_bottom_1_top_width_0_height_0__pin_1_upper ) , 
    .top_width_0_height_0__pin_1_lower ( grid_io_bottom_1_top_width_0_height_0__pin_1_lower ) , 
    .ccff_tail ( grid_io_bottom_1_ccff_tail ) ) ;
grid_io_bottom grid_io_bottom_3__0_ (
    .prog_clk ( { ctsbuf_net_3302312 } ) ,
    .gfpga_pad_GPIO_A ( gfpga_pad_GPIO_A[26] ) , 
    .gfpga_pad_GPIO_IE ( gfpga_pad_GPIO_IE[26] ) , 
    .gfpga_pad_GPIO_OE ( gfpga_pad_GPIO_OE[26] ) , 
    .gfpga_pad_GPIO_Y ( gfpga_pad_GPIO_Y[26] ) , 
    .top_width_0_height_0__pin_0_ ( cbx_1__0__2_bottom_grid_pin_0_ ) , 
    .ccff_head ( cbx_1__0__2_ccff_tail ) , 
    .top_width_0_height_0__pin_1_upper ( grid_io_bottom_2_top_width_0_height_0__pin_1_upper ) , 
    .top_width_0_height_0__pin_1_lower ( grid_io_bottom_2_top_width_0_height_0__pin_1_lower ) , 
    .ccff_tail ( grid_io_bottom_2_ccff_tail ) ) ;
grid_io_bottom grid_io_bottom_4__0_ (
    .prog_clk ( { ctsbuf_net_2842266 } ) ,
    .gfpga_pad_GPIO_A ( gfpga_pad_GPIO_A[27] ) , 
    .gfpga_pad_GPIO_IE ( gfpga_pad_GPIO_IE[27] ) , 
    .gfpga_pad_GPIO_OE ( gfpga_pad_GPIO_OE[27] ) , 
    .gfpga_pad_GPIO_Y ( gfpga_pad_GPIO_Y[27] ) , 
    .top_width_0_height_0__pin_0_ ( cbx_1__0__3_bottom_grid_pin_0_ ) , 
    .ccff_head ( cbx_1__0__3_ccff_tail ) , 
    .top_width_0_height_0__pin_1_upper ( grid_io_bottom_3_top_width_0_height_0__pin_1_upper ) , 
    .top_width_0_height_0__pin_1_lower ( grid_io_bottom_3_top_width_0_height_0__pin_1_lower ) , 
    .ccff_tail ( grid_io_bottom_3_ccff_tail ) ) ;
grid_io_bottom grid_io_bottom_5__0_ (
    .prog_clk ( { ctsbuf_net_2402222 } ) ,
    .gfpga_pad_GPIO_A ( gfpga_pad_GPIO_A[28] ) , 
    .gfpga_pad_GPIO_IE ( gfpga_pad_GPIO_IE[28] ) , 
    .gfpga_pad_GPIO_OE ( gfpga_pad_GPIO_OE[28] ) , 
    .gfpga_pad_GPIO_Y ( gfpga_pad_GPIO_Y[28] ) , 
    .top_width_0_height_0__pin_0_ ( cbx_1__0__4_bottom_grid_pin_0_ ) , 
    .ccff_head ( cbx_1__0__4_ccff_tail ) , 
    .top_width_0_height_0__pin_1_upper ( grid_io_bottom_4_top_width_0_height_0__pin_1_upper ) , 
    .top_width_0_height_0__pin_1_lower ( grid_io_bottom_4_top_width_0_height_0__pin_1_lower ) , 
    .ccff_tail ( grid_io_bottom_4_ccff_tail ) ) ;
grid_io_bottom grid_io_bottom_6__0_ (
    .prog_clk ( { ctsbuf_net_1942176 } ) ,
    .gfpga_pad_GPIO_A ( gfpga_pad_GPIO_A[29] ) , 
    .gfpga_pad_GPIO_IE ( gfpga_pad_GPIO_IE[29] ) , 
    .gfpga_pad_GPIO_OE ( gfpga_pad_GPIO_OE[29] ) , 
    .gfpga_pad_GPIO_Y ( gfpga_pad_GPIO_Y[29] ) , 
    .top_width_0_height_0__pin_0_ ( cbx_1__0__5_bottom_grid_pin_0_ ) , 
    .ccff_head ( cbx_1__0__5_ccff_tail ) , 
    .top_width_0_height_0__pin_1_upper ( grid_io_bottom_5_top_width_0_height_0__pin_1_upper ) , 
    .top_width_0_height_0__pin_1_lower ( grid_io_bottom_5_top_width_0_height_0__pin_1_lower ) , 
    .ccff_tail ( grid_io_bottom_5_ccff_tail ) ) ;
grid_io_bottom grid_io_bottom_7__0_ (
    .prog_clk ( { ctsbuf_net_1542136 } ) ,
    .gfpga_pad_GPIO_A ( gfpga_pad_GPIO_A[30] ) , 
    .gfpga_pad_GPIO_IE ( gfpga_pad_GPIO_IE[30] ) , 
    .gfpga_pad_GPIO_OE ( gfpga_pad_GPIO_OE[30] ) , 
    .gfpga_pad_GPIO_Y ( gfpga_pad_GPIO_Y[30] ) , 
    .top_width_0_height_0__pin_0_ ( cbx_1__0__6_bottom_grid_pin_0_ ) , 
    .ccff_head ( cbx_1__0__6_ccff_tail ) , 
    .top_width_0_height_0__pin_1_upper ( grid_io_bottom_6_top_width_0_height_0__pin_1_upper ) , 
    .top_width_0_height_0__pin_1_lower ( grid_io_bottom_6_top_width_0_height_0__pin_1_lower ) , 
    .ccff_tail ( grid_io_bottom_6_ccff_tail ) ) ;
grid_io_bottom grid_io_bottom_8__0_ (
    .prog_clk ( { ctsbuf_net_1212103 } ) ,
    .gfpga_pad_GPIO_A ( gfpga_pad_GPIO_A[31] ) , 
    .gfpga_pad_GPIO_IE ( gfpga_pad_GPIO_IE[31] ) , 
    .gfpga_pad_GPIO_OE ( gfpga_pad_GPIO_OE[31] ) , 
    .gfpga_pad_GPIO_Y ( gfpga_pad_GPIO_Y[31] ) , 
    .top_width_0_height_0__pin_0_ ( cbx_1__0__7_bottom_grid_pin_0_ ) , 
    .ccff_head ( cbx_1__0__7_ccff_tail ) , 
    .top_width_0_height_0__pin_1_upper ( grid_io_bottom_7_top_width_0_height_0__pin_1_upper ) , 
    .top_width_0_height_0__pin_1_lower ( grid_io_bottom_7_top_width_0_height_0__pin_1_lower ) , 
    .ccff_tail ( grid_io_bottom_7_ccff_tail ) ) ;
grid_io_bottom grid_io_bottom_9__0_ (
    .prog_clk ( { ctsbuf_net_932075 } ) ,
    .gfpga_pad_GPIO_A ( gfpga_pad_GPIO_A[32] ) , 
    .gfpga_pad_GPIO_IE ( gfpga_pad_GPIO_IE[32] ) , 
    .gfpga_pad_GPIO_OE ( gfpga_pad_GPIO_OE[32] ) , 
    .gfpga_pad_GPIO_Y ( gfpga_pad_GPIO_Y[32] ) , 
    .top_width_0_height_0__pin_0_ ( cbx_1__0__8_bottom_grid_pin_0_ ) , 
    .ccff_head ( cbx_1__0__8_ccff_tail ) , 
    .top_width_0_height_0__pin_1_upper ( grid_io_bottom_8_top_width_0_height_0__pin_1_upper ) , 
    .top_width_0_height_0__pin_1_lower ( grid_io_bottom_8_top_width_0_height_0__pin_1_lower ) , 
    .ccff_tail ( grid_io_bottom_8_ccff_tail ) ) ;
grid_io_bottom grid_io_bottom_10__0_ (
    .prog_clk ( { ctsbuf_net_692051 } ) ,
    .gfpga_pad_GPIO_A ( gfpga_pad_GPIO_A[33] ) , 
    .gfpga_pad_GPIO_IE ( gfpga_pad_GPIO_IE[33] ) , 
    .gfpga_pad_GPIO_OE ( gfpga_pad_GPIO_OE[33] ) , 
    .gfpga_pad_GPIO_Y ( gfpga_pad_GPIO_Y[33] ) , 
    .top_width_0_height_0__pin_0_ ( cbx_1__0__9_bottom_grid_pin_0_ ) , 
    .ccff_head ( cbx_1__0__9_ccff_tail ) , 
    .top_width_0_height_0__pin_1_upper ( grid_io_bottom_9_top_width_0_height_0__pin_1_upper ) , 
    .top_width_0_height_0__pin_1_lower ( grid_io_bottom_9_top_width_0_height_0__pin_1_lower ) , 
    .ccff_tail ( grid_io_bottom_9_ccff_tail ) ) ;
grid_io_bottom grid_io_bottom_11__0_ (
    .prog_clk ( { ctsbuf_net_542036 } ) ,
    .gfpga_pad_GPIO_A ( gfpga_pad_GPIO_A[34] ) , 
    .gfpga_pad_GPIO_IE ( gfpga_pad_GPIO_IE[34] ) , 
    .gfpga_pad_GPIO_OE ( gfpga_pad_GPIO_OE[34] ) , 
    .gfpga_pad_GPIO_Y ( gfpga_pad_GPIO_Y[34] ) , 
    .top_width_0_height_0__pin_0_ ( cbx_1__0__10_bottom_grid_pin_0_ ) , 
    .ccff_head ( cbx_1__0__10_ccff_tail ) , 
    .top_width_0_height_0__pin_1_upper ( grid_io_bottom_10_top_width_0_height_0__pin_1_upper ) , 
    .top_width_0_height_0__pin_1_lower ( grid_io_bottom_10_top_width_0_height_0__pin_1_lower ) , 
    .ccff_tail ( grid_io_bottom_10_ccff_tail ) ) ;
grid_io_bottom grid_io_bottom_12__0_ (
    .prog_clk ( { ctsbuf_net_482030 } ) ,
    .gfpga_pad_GPIO_A ( gfpga_pad_GPIO_A[35] ) , 
    .gfpga_pad_GPIO_IE ( gfpga_pad_GPIO_IE[35] ) , 
    .gfpga_pad_GPIO_OE ( gfpga_pad_GPIO_OE[35] ) , 
    .gfpga_pad_GPIO_Y ( gfpga_pad_GPIO_Y[35] ) , 
    .top_width_0_height_0__pin_0_ ( cbx_1__0__11_bottom_grid_pin_0_ ) , 
    .ccff_head ( cbx_1__0__11_ccff_tail ) , 
    .top_width_0_height_0__pin_1_upper ( grid_io_bottom_11_top_width_0_height_0__pin_1_upper ) , 
    .top_width_0_height_0__pin_1_lower ( grid_io_bottom_11_top_width_0_height_0__pin_1_lower ) , 
    .ccff_tail ( grid_io_bottom_11_ccff_tail ) ) ;
grid_io_left grid_io_left_0__1_ (
    .prog_clk ( { ctsbuf_net_4542436 } ) ,
    .gfpga_pad_GPIO_A ( gfpga_pad_GPIO_A[36] ) , 
    .gfpga_pad_GPIO_IE ( gfpga_pad_GPIO_IE[36] ) , 
    .gfpga_pad_GPIO_OE ( gfpga_pad_GPIO_OE[36] ) , 
    .gfpga_pad_GPIO_Y ( gfpga_pad_GPIO_Y[36] ) , 
    .right_width_0_height_0__pin_0_ ( cby_0__1__0_left_grid_pin_0_ ) , 
    .ccff_head ( cby_0__1__0_ccff_tail ) , 
    .right_width_0_height_0__pin_1_upper ( grid_io_left_0_right_width_0_height_0__pin_1_upper ) , 
    .right_width_0_height_0__pin_1_lower ( grid_io_left_0_right_width_0_height_0__pin_1_lower ) , 
    .ccff_tail ( grid_io_left_0_ccff_tail ) ) ;
grid_io_left grid_io_left_0__2_ (
    .prog_clk ( { ctsbuf_net_4942476 } ) ,
    .gfpga_pad_GPIO_A ( gfpga_pad_GPIO_A[37] ) , 
    .gfpga_pad_GPIO_IE ( gfpga_pad_GPIO_IE[37] ) , 
    .gfpga_pad_GPIO_OE ( gfpga_pad_GPIO_OE[37] ) , 
    .gfpga_pad_GPIO_Y ( gfpga_pad_GPIO_Y[37] ) , 
    .right_width_0_height_0__pin_0_ ( cby_0__1__1_left_grid_pin_0_ ) , 
    .ccff_head ( cby_0__1__1_ccff_tail ) , 
    .right_width_0_height_0__pin_1_upper ( grid_io_left_1_right_width_0_height_0__pin_1_upper ) , 
    .right_width_0_height_0__pin_1_lower ( grid_io_left_1_right_width_0_height_0__pin_1_lower ) , 
    .ccff_tail ( grid_io_left_1_ccff_tail ) ) ;
grid_io_left grid_io_left_0__3_ (
    .prog_clk ( { ctsbuf_net_5252507 } ) ,
    .gfpga_pad_GPIO_A ( gfpga_pad_GPIO_A[38] ) , 
    .gfpga_pad_GPIO_IE ( gfpga_pad_GPIO_IE[38] ) , 
    .gfpga_pad_GPIO_OE ( gfpga_pad_GPIO_OE[38] ) , 
    .gfpga_pad_GPIO_Y ( gfpga_pad_GPIO_Y[38] ) , 
    .right_width_0_height_0__pin_0_ ( cby_0__1__2_left_grid_pin_0_ ) , 
    .ccff_head ( cby_0__1__2_ccff_tail ) , 
    .right_width_0_height_0__pin_1_upper ( grid_io_left_2_right_width_0_height_0__pin_1_upper ) , 
    .right_width_0_height_0__pin_1_lower ( grid_io_left_2_right_width_0_height_0__pin_1_lower ) , 
    .ccff_tail ( grid_io_left_2_ccff_tail ) ) ;
grid_io_left grid_io_left_0__4_ (
    .prog_clk ( { ctsbuf_net_5512533 } ) ,
    .gfpga_pad_GPIO_A ( gfpga_pad_GPIO_A[39] ) , 
    .gfpga_pad_GPIO_IE ( gfpga_pad_GPIO_IE[39] ) , 
    .gfpga_pad_GPIO_OE ( gfpga_pad_GPIO_OE[39] ) , 
    .gfpga_pad_GPIO_Y ( gfpga_pad_GPIO_Y[39] ) , 
    .right_width_0_height_0__pin_0_ ( cby_0__1__3_left_grid_pin_0_ ) , 
    .ccff_head ( cby_0__1__3_ccff_tail ) , 
    .right_width_0_height_0__pin_1_upper ( grid_io_left_3_right_width_0_height_0__pin_1_upper ) , 
    .right_width_0_height_0__pin_1_lower ( grid_io_left_3_right_width_0_height_0__pin_1_lower ) , 
    .ccff_tail ( grid_io_left_3_ccff_tail ) ) ;
grid_io_left grid_io_left_0__5_ (
    .prog_clk ( { ctsbuf_net_5692551 } ) ,
    .gfpga_pad_GPIO_A ( gfpga_pad_GPIO_A[40] ) , 
    .gfpga_pad_GPIO_IE ( gfpga_pad_GPIO_IE[40] ) , 
    .gfpga_pad_GPIO_OE ( gfpga_pad_GPIO_OE[40] ) , 
    .gfpga_pad_GPIO_Y ( gfpga_pad_GPIO_Y[40] ) , 
    .right_width_0_height_0__pin_0_ ( cby_0__1__4_left_grid_pin_0_ ) , 
    .ccff_head ( cby_0__1__4_ccff_tail ) , 
    .right_width_0_height_0__pin_1_upper ( grid_io_left_4_right_width_0_height_0__pin_1_upper ) , 
    .right_width_0_height_0__pin_1_lower ( grid_io_left_4_right_width_0_height_0__pin_1_lower ) , 
    .ccff_tail ( grid_io_left_4_ccff_tail ) ) ;
grid_io_left grid_io_left_0__6_ (
    .prog_clk ( { ctsbuf_net_5802562 } ) ,
    .gfpga_pad_GPIO_A ( gfpga_pad_GPIO_A[41] ) , 
    .gfpga_pad_GPIO_IE ( gfpga_pad_GPIO_IE[41] ) , 
    .gfpga_pad_GPIO_OE ( gfpga_pad_GPIO_OE[41] ) , 
    .gfpga_pad_GPIO_Y ( gfpga_pad_GPIO_Y[41] ) , 
    .right_width_0_height_0__pin_0_ ( cby_0__1__5_left_grid_pin_0_ ) , 
    .ccff_head ( cby_0__1__5_ccff_tail ) , 
    .right_width_0_height_0__pin_1_upper ( grid_io_left_5_right_width_0_height_0__pin_1_upper ) , 
    .right_width_0_height_0__pin_1_lower ( grid_io_left_5_right_width_0_height_0__pin_1_lower ) , 
    .ccff_tail ( grid_io_left_5_ccff_tail ) ) ;
grid_io_left grid_io_left_0__7_ (
    .prog_clk ( { ctsbuf_net_5772559 } ) ,
    .gfpga_pad_GPIO_A ( gfpga_pad_GPIO_A[42] ) , 
    .gfpga_pad_GPIO_IE ( gfpga_pad_GPIO_IE[42] ) , 
    .gfpga_pad_GPIO_OE ( gfpga_pad_GPIO_OE[42] ) , 
    .gfpga_pad_GPIO_Y ( gfpga_pad_GPIO_Y[42] ) , 
    .right_width_0_height_0__pin_0_ ( cby_0__1__6_left_grid_pin_0_ ) , 
    .ccff_head ( cby_0__1__6_ccff_tail ) , 
    .right_width_0_height_0__pin_1_upper ( grid_io_left_6_right_width_0_height_0__pin_1_upper ) , 
    .right_width_0_height_0__pin_1_lower ( grid_io_left_6_right_width_0_height_0__pin_1_lower ) , 
    .ccff_tail ( grid_io_left_6_ccff_tail ) ) ;
grid_io_left grid_io_left_0__8_ (
    .prog_clk ( { ctsbuf_net_5772559 } ) ,
    .gfpga_pad_GPIO_A ( gfpga_pad_GPIO_A[43] ) , 
    .gfpga_pad_GPIO_IE ( gfpga_pad_GPIO_IE[43] ) , 
    .gfpga_pad_GPIO_OE ( gfpga_pad_GPIO_OE[43] ) , 
    .gfpga_pad_GPIO_Y ( gfpga_pad_GPIO_Y[43] ) , 
    .right_width_0_height_0__pin_0_ ( cby_0__1__7_left_grid_pin_0_ ) , 
    .ccff_head ( cby_0__1__7_ccff_tail ) , 
    .right_width_0_height_0__pin_1_upper ( grid_io_left_7_right_width_0_height_0__pin_1_upper ) , 
    .right_width_0_height_0__pin_1_lower ( grid_io_left_7_right_width_0_height_0__pin_1_lower ) , 
    .ccff_tail ( grid_io_left_7_ccff_tail ) ) ;
grid_io_left grid_io_left_0__9_ (
    .prog_clk ( { ctsbuf_net_5442526 } ) ,
    .gfpga_pad_GPIO_A ( gfpga_pad_GPIO_A[44] ) , 
    .gfpga_pad_GPIO_IE ( gfpga_pad_GPIO_IE[44] ) , 
    .gfpga_pad_GPIO_OE ( gfpga_pad_GPIO_OE[44] ) , 
    .gfpga_pad_GPIO_Y ( gfpga_pad_GPIO_Y[44] ) , 
    .right_width_0_height_0__pin_0_ ( cby_0__1__8_left_grid_pin_0_ ) , 
    .ccff_head ( cby_0__1__8_ccff_tail ) , 
    .right_width_0_height_0__pin_1_upper ( grid_io_left_8_right_width_0_height_0__pin_1_upper ) , 
    .right_width_0_height_0__pin_1_lower ( grid_io_left_8_right_width_0_height_0__pin_1_lower ) , 
    .ccff_tail ( grid_io_left_8_ccff_tail ) ) ;
grid_io_left grid_io_left_0__10_ (
    .prog_clk ( { ctsbuf_net_5442526 } ) ,
    .gfpga_pad_GPIO_A ( gfpga_pad_GPIO_A[45] ) , 
    .gfpga_pad_GPIO_IE ( gfpga_pad_GPIO_IE[45] ) , 
    .gfpga_pad_GPIO_OE ( gfpga_pad_GPIO_OE[45] ) , 
    .gfpga_pad_GPIO_Y ( gfpga_pad_GPIO_Y[45] ) , 
    .right_width_0_height_0__pin_0_ ( cby_0__1__9_left_grid_pin_0_ ) , 
    .ccff_head ( cby_0__1__9_ccff_tail ) , 
    .right_width_0_height_0__pin_1_upper ( grid_io_left_9_right_width_0_height_0__pin_1_upper ) , 
    .right_width_0_height_0__pin_1_lower ( grid_io_left_9_right_width_0_height_0__pin_1_lower ) , 
    .ccff_tail ( grid_io_left_9_ccff_tail ) ) ;
grid_io_left grid_io_left_0__11_ (
    .prog_clk ( { ctsbuf_net_4832465 } ) ,
    .gfpga_pad_GPIO_A ( gfpga_pad_GPIO_A[46] ) , 
    .gfpga_pad_GPIO_IE ( gfpga_pad_GPIO_IE[46] ) , 
    .gfpga_pad_GPIO_OE ( gfpga_pad_GPIO_OE[46] ) , 
    .gfpga_pad_GPIO_Y ( gfpga_pad_GPIO_Y[46] ) , 
    .right_width_0_height_0__pin_0_ ( cby_0__1__10_left_grid_pin_0_ ) , 
    .ccff_head ( cby_0__1__10_ccff_tail ) , 
    .right_width_0_height_0__pin_1_upper ( grid_io_left_10_right_width_0_height_0__pin_1_upper ) , 
    .right_width_0_height_0__pin_1_lower ( grid_io_left_10_right_width_0_height_0__pin_1_lower ) , 
    .ccff_tail ( grid_io_left_10_ccff_tail ) ) ;
grid_io_left grid_io_left_0__12_ (
    .prog_clk ( { ctsbuf_net_4832465 } ) ,
    .gfpga_pad_GPIO_A ( gfpga_pad_GPIO_A[47] ) , 
    .gfpga_pad_GPIO_IE ( gfpga_pad_GPIO_IE[47] ) , 
    .gfpga_pad_GPIO_OE ( gfpga_pad_GPIO_OE[47] ) , 
    .gfpga_pad_GPIO_Y ( gfpga_pad_GPIO_Y[47] ) , 
    .right_width_0_height_0__pin_0_ ( cby_0__1__11_left_grid_pin_0_ ) , 
    .ccff_head ( cby_0__1__11_ccff_tail ) , 
    .right_width_0_height_0__pin_1_upper ( grid_io_left_11_right_width_0_height_0__pin_1_upper ) , 
    .right_width_0_height_0__pin_1_lower ( grid_io_left_11_right_width_0_height_0__pin_1_lower ) , 
    .ccff_tail ( grid_io_left_11_ccff_tail ) ) ;
sb_0__0_ sb_0__0_ (
    .prog_clk ( { ctsbuf_net_4172399 } ) ,
    .chany_top_in ( cby_0__1__0_chany_bottom_out ) , 
    .top_left_grid_pin_1_ ( grid_io_left_0_right_width_0_height_0__pin_1_lower ) , 
    .chanx_right_in ( cbx_1__0__0_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_0_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_0_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_0_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_0_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_0_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_0_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_0_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_0_bottom_width_0_height_0__pin_49_upper ) , 
    .right_bottom_grid_pin_1_ ( grid_io_bottom_0_top_width_0_height_0__pin_1_upper ) , 
    .ccff_head ( grid_io_bottom_0_ccff_tail ) , 
    .chany_top_out ( sb_0__0__0_chany_top_out ) , 
    .chanx_right_out ( sb_0__0__0_chanx_right_out ) , 
    .ccff_tail ( ccff_tail ) ) ;
sb_0__1_ sb_0__1_ (
    .prog_clk ( { ctsbuf_net_4542436 } ) ,
    .chany_top_in ( cby_0__1__1_chany_bottom_out ) , 
    .top_left_grid_pin_1_ ( grid_io_left_1_right_width_0_height_0__pin_1_lower ) , 
    .chanx_right_in ( cbx_1__1__0_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_1_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_1_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_1_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_1_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_1_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_1_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_1_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_1_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_0__1__0_chany_top_out ) , 
    .bottom_left_grid_pin_1_ ( grid_io_left_0_right_width_0_height_0__pin_1_upper ) , 
    .ccff_head ( cbx_1__1__0_ccff_tail ) , 
    .chany_top_out ( sb_0__1__0_chany_top_out ) , 
    .chanx_right_out ( sb_0__1__0_chanx_right_out ) , 
    .chany_bottom_out ( sb_0__1__0_chany_bottom_out ) , 
    .ccff_tail ( sb_0__1__0_ccff_tail ) ) ;
sb_0__1_ sb_0__2_ (
    .prog_clk ( { ctsbuf_net_4942476 } ) ,
    .chany_top_in ( cby_0__1__2_chany_bottom_out ) , 
    .top_left_grid_pin_1_ ( grid_io_left_2_right_width_0_height_0__pin_1_lower ) , 
    .chanx_right_in ( cbx_1__1__1_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_2_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_2_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_2_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_2_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_2_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_2_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_2_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_2_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_0__1__1_chany_top_out ) , 
    .bottom_left_grid_pin_1_ ( grid_io_left_1_right_width_0_height_0__pin_1_upper ) , 
    .ccff_head ( cbx_1__1__1_ccff_tail ) , 
    .chany_top_out ( sb_0__1__1_chany_top_out ) , 
    .chanx_right_out ( sb_0__1__1_chanx_right_out ) , 
    .chany_bottom_out ( sb_0__1__1_chany_bottom_out ) , 
    .ccff_tail ( sb_0__1__1_ccff_tail ) ) ;
sb_0__1_ sb_0__3_ (
    .prog_clk ( { ctsbuf_net_5252507 } ) ,
    .chany_top_in ( cby_0__1__3_chany_bottom_out ) , 
    .top_left_grid_pin_1_ ( grid_io_left_3_right_width_0_height_0__pin_1_lower ) , 
    .chanx_right_in ( cbx_1__1__2_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_3_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_3_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_3_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_3_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_3_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_3_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_3_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_3_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_0__1__2_chany_top_out ) , 
    .bottom_left_grid_pin_1_ ( grid_io_left_2_right_width_0_height_0__pin_1_upper ) , 
    .ccff_head ( cbx_1__1__2_ccff_tail ) , 
    .chany_top_out ( sb_0__1__2_chany_top_out ) , 
    .chanx_right_out ( sb_0__1__2_chanx_right_out ) , 
    .chany_bottom_out ( sb_0__1__2_chany_bottom_out ) , 
    .ccff_tail ( sb_0__1__2_ccff_tail ) ) ;
sb_0__1_ sb_0__4_ (
    .prog_clk ( { ctsbuf_net_5512533 } ) ,
    .chany_top_in ( cby_0__1__4_chany_bottom_out ) , 
    .top_left_grid_pin_1_ ( grid_io_left_4_right_width_0_height_0__pin_1_lower ) , 
    .chanx_right_in ( cbx_1__1__3_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_4_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_4_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_4_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_4_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_4_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_4_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_4_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_4_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_0__1__3_chany_top_out ) , 
    .bottom_left_grid_pin_1_ ( grid_io_left_3_right_width_0_height_0__pin_1_upper ) , 
    .ccff_head ( cbx_1__1__3_ccff_tail ) , 
    .chany_top_out ( sb_0__1__3_chany_top_out ) , 
    .chanx_right_out ( sb_0__1__3_chanx_right_out ) , 
    .chany_bottom_out ( sb_0__1__3_chany_bottom_out ) , 
    .ccff_tail ( sb_0__1__3_ccff_tail ) ) ;
sb_0__1_ sb_0__5_ (
    .prog_clk ( { ctsbuf_net_5692551 } ) ,
    .chany_top_in ( cby_0__1__5_chany_bottom_out ) , 
    .top_left_grid_pin_1_ ( grid_io_left_5_right_width_0_height_0__pin_1_lower ) , 
    .chanx_right_in ( cbx_1__1__4_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_5_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_5_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_5_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_5_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_5_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_5_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_5_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_5_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_0__1__4_chany_top_out ) , 
    .bottom_left_grid_pin_1_ ( grid_io_left_4_right_width_0_height_0__pin_1_upper ) , 
    .ccff_head ( cbx_1__1__4_ccff_tail ) , 
    .chany_top_out ( sb_0__1__4_chany_top_out ) , 
    .chanx_right_out ( sb_0__1__4_chanx_right_out ) , 
    .chany_bottom_out ( sb_0__1__4_chany_bottom_out ) , 
    .ccff_tail ( sb_0__1__4_ccff_tail ) ) ;
sb_0__1_ sb_0__6_ (
    .prog_clk ( { ctsbuf_net_5802562 } ) ,
    .chany_top_in ( cby_0__1__6_chany_bottom_out ) , 
    .top_left_grid_pin_1_ ( grid_io_left_6_right_width_0_height_0__pin_1_lower ) , 
    .chanx_right_in ( cbx_1__1__5_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_6_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_6_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_6_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_6_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_6_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_6_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_6_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_6_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_0__1__5_chany_top_out ) , 
    .bottom_left_grid_pin_1_ ( grid_io_left_5_right_width_0_height_0__pin_1_upper ) , 
    .ccff_head ( cbx_1__1__5_ccff_tail ) , 
    .chany_top_out ( sb_0__1__5_chany_top_out ) , 
    .chanx_right_out ( sb_0__1__5_chanx_right_out ) , 
    .chany_bottom_out ( sb_0__1__5_chany_bottom_out ) , 
    .ccff_tail ( sb_0__1__5_ccff_tail ) ) ;
sb_0__1_ sb_0__7_ (
    .prog_clk ( { ctsbuf_net_5752557 } ) ,
    .chany_top_in ( cby_0__1__7_chany_bottom_out ) , 
    .top_left_grid_pin_1_ ( grid_io_left_7_right_width_0_height_0__pin_1_lower ) , 
    .chanx_right_in ( cbx_1__1__6_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_7_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_7_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_7_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_7_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_7_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_7_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_7_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_7_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_0__1__6_chany_top_out ) , 
    .bottom_left_grid_pin_1_ ( grid_io_left_6_right_width_0_height_0__pin_1_upper ) , 
    .ccff_head ( cbx_1__1__6_ccff_tail ) , 
    .chany_top_out ( sb_0__1__6_chany_top_out ) , 
    .chanx_right_out ( sb_0__1__6_chanx_right_out ) , 
    .chany_bottom_out ( sb_0__1__6_chany_bottom_out ) , 
    .ccff_tail ( sb_0__1__6_ccff_tail ) ) ;
sb_0__1_ sb_0__8_ (
    .prog_clk ( { ctsbuf_net_5642546 } ) ,
    .chany_top_in ( cby_0__1__8_chany_bottom_out ) , 
    .top_left_grid_pin_1_ ( grid_io_left_8_right_width_0_height_0__pin_1_lower ) , 
    .chanx_right_in ( cbx_1__1__7_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_8_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_8_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_8_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_8_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_8_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_8_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_8_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_8_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_0__1__7_chany_top_out ) , 
    .bottom_left_grid_pin_1_ ( grid_io_left_7_right_width_0_height_0__pin_1_upper ) , 
    .ccff_head ( cbx_1__1__7_ccff_tail ) , 
    .chany_top_out ( sb_0__1__7_chany_top_out ) , 
    .chanx_right_out ( sb_0__1__7_chanx_right_out ) , 
    .chany_bottom_out ( sb_0__1__7_chany_bottom_out ) , 
    .ccff_tail ( sb_0__1__7_ccff_tail ) ) ;
sb_0__1_ sb_0__9_ (
    .prog_clk ( { ctsbuf_net_5392521 } ) ,
    .chany_top_in ( cby_0__1__9_chany_bottom_out ) , 
    .top_left_grid_pin_1_ ( grid_io_left_9_right_width_0_height_0__pin_1_lower ) , 
    .chanx_right_in ( cbx_1__1__8_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_9_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_9_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_9_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_9_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_9_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_9_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_9_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_9_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_0__1__8_chany_top_out ) , 
    .bottom_left_grid_pin_1_ ( grid_io_left_8_right_width_0_height_0__pin_1_upper ) , 
    .ccff_head ( cbx_1__1__8_ccff_tail ) , 
    .chany_top_out ( sb_0__1__8_chany_top_out ) , 
    .chanx_right_out ( sb_0__1__8_chanx_right_out ) , 
    .chany_bottom_out ( sb_0__1__8_chany_bottom_out ) , 
    .ccff_tail ( sb_0__1__8_ccff_tail ) ) ;
sb_0__1_ sb_0__10_ (
    .prog_clk ( { ctsbuf_net_5162498 } ) ,
    .chany_top_in ( cby_0__1__10_chany_bottom_out ) , 
    .top_left_grid_pin_1_ ( grid_io_left_10_right_width_0_height_0__pin_1_lower ) , 
    .chanx_right_in ( cbx_1__1__9_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_10_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_10_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_10_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_10_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_10_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_10_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_10_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_10_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_0__1__9_chany_top_out ) , 
    .bottom_left_grid_pin_1_ ( grid_io_left_9_right_width_0_height_0__pin_1_upper ) , 
    .ccff_head ( cbx_1__1__9_ccff_tail ) , 
    .chany_top_out ( sb_0__1__9_chany_top_out ) , 
    .chanx_right_out ( sb_0__1__9_chanx_right_out ) , 
    .chany_bottom_out ( sb_0__1__9_chany_bottom_out ) , 
    .ccff_tail ( sb_0__1__9_ccff_tail ) ) ;
sb_0__1_ sb_0__11_ (
    .prog_clk ( { ctsbuf_net_4752457 } ) ,
    .chany_top_in ( cby_0__1__11_chany_bottom_out ) , 
    .top_left_grid_pin_1_ ( grid_io_left_11_right_width_0_height_0__pin_1_lower ) , 
    .chanx_right_in ( cbx_1__1__10_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_11_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_11_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_11_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_11_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_11_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_11_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_11_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_11_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_0__1__10_chany_top_out ) , 
    .bottom_left_grid_pin_1_ ( grid_io_left_10_right_width_0_height_0__pin_1_upper ) , 
    .ccff_head ( cbx_1__1__10_ccff_tail ) , 
    .chany_top_out ( sb_0__1__10_chany_top_out ) , 
    .chanx_right_out ( sb_0__1__10_chanx_right_out ) , 
    .chany_bottom_out ( sb_0__1__10_chany_bottom_out ) , 
    .ccff_tail ( sb_0__1__10_ccff_tail ) ) ;
sb_0__2_ sb_0__12_ (
    .prog_clk ( { ctsbuf_net_4162398 } ) ,
    .chanx_right_in ( cbx_1__12__0_chanx_left_out ) , 
    .right_top_grid_pin_1_ ( grid_io_top_0_bottom_width_0_height_0__pin_1_upper ) , 
    .chany_bottom_in ( cby_0__1__11_chany_top_out ) , 
    .bottom_left_grid_pin_1_ ( grid_io_left_11_right_width_0_height_0__pin_1_upper ) , 
    .ccff_head ( grid_io_top_0_ccff_tail ) , 
    .chanx_right_out ( sb_0__12__0_chanx_right_out ) , 
    .chany_bottom_out ( sb_0__12__0_chany_bottom_out ) , 
    .ccff_tail ( sb_0__12__0_ccff_tail ) ) ;
sb_1__0_ sb_1__0_ (
    .prog_clk ( { ctsbuf_net_4112393 } ) ,
    .chany_top_in ( cby_1__1__0_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_0_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_0_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_0_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_0_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_0_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_0_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_0_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_0_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__0__1_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_12_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_12_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_12_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_12_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_12_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_12_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_12_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_12_bottom_width_0_height_0__pin_49_upper ) , 
    .right_bottom_grid_pin_1_ ( grid_io_bottom_1_top_width_0_height_0__pin_1_upper ) , 
    .chanx_left_in ( cbx_1__0__0_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_0_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_0_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_0_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_0_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_0_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_0_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_0_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_0_bottom_width_0_height_0__pin_49_lower ) , 
    .left_bottom_grid_pin_1_ ( grid_io_bottom_0_top_width_0_height_0__pin_1_lower ) , 
    .ccff_head ( grid_io_bottom_1_ccff_tail ) , 
    .chany_top_out ( sb_1__0__0_chany_top_out ) , 
    .chanx_right_out ( sb_1__0__0_chanx_right_out ) , 
    .chanx_left_out ( sb_1__0__0_chanx_left_out ) , 
    .ccff_tail ( sb_1__0__0_ccff_tail ) ) ;
sb_1__0_ sb_2__0_ (
    .prog_clk ( { ctsbuf_net_3682350 } ) ,
    .chany_top_in ( cby_1__1__12_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_12_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_12_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_12_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_12_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_12_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_12_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_12_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_12_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__0__2_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_24_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_24_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_24_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_24_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_24_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_24_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_24_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_24_bottom_width_0_height_0__pin_49_upper ) , 
    .right_bottom_grid_pin_1_ ( grid_io_bottom_2_top_width_0_height_0__pin_1_upper ) , 
    .chanx_left_in ( cbx_1__0__1_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_12_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_12_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_12_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_12_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_12_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_12_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_12_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_12_bottom_width_0_height_0__pin_49_lower ) , 
    .left_bottom_grid_pin_1_ ( grid_io_bottom_1_top_width_0_height_0__pin_1_lower ) , 
    .ccff_head ( grid_io_bottom_2_ccff_tail ) , 
    .chany_top_out ( sb_1__0__1_chany_top_out ) , 
    .chanx_right_out ( sb_1__0__1_chanx_right_out ) , 
    .chanx_left_out ( sb_1__0__1_chanx_left_out ) , 
    .ccff_tail ( sb_1__0__1_ccff_tail ) ) ;
sb_1__0_ sb_3__0_ (
    .prog_clk ( { ctsbuf_net_3242306 } ) ,
    .chany_top_in ( cby_1__1__24_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_24_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_24_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_24_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_24_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_24_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_24_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_24_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_24_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__0__3_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_36_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_36_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_36_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_36_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_36_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_36_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_36_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_36_bottom_width_0_height_0__pin_49_upper ) , 
    .right_bottom_grid_pin_1_ ( grid_io_bottom_3_top_width_0_height_0__pin_1_upper ) , 
    .chanx_left_in ( cbx_1__0__2_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_24_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_24_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_24_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_24_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_24_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_24_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_24_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_24_bottom_width_0_height_0__pin_49_lower ) , 
    .left_bottom_grid_pin_1_ ( grid_io_bottom_2_top_width_0_height_0__pin_1_lower ) , 
    .ccff_head ( grid_io_bottom_3_ccff_tail ) , 
    .chany_top_out ( sb_1__0__2_chany_top_out ) , 
    .chanx_right_out ( sb_1__0__2_chanx_right_out ) , 
    .chanx_left_out ( sb_1__0__2_chanx_left_out ) , 
    .ccff_tail ( sb_1__0__2_ccff_tail ) ) ;
sb_1__0_ sb_4__0_ (
    .prog_clk ( { ctsbuf_net_2792261 } ) ,
    .chany_top_in ( cby_1__1__36_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_36_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_36_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_36_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_36_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_36_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_36_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_36_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_36_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__0__4_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_48_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_48_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_48_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_48_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_48_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_48_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_48_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_48_bottom_width_0_height_0__pin_49_upper ) , 
    .right_bottom_grid_pin_1_ ( grid_io_bottom_4_top_width_0_height_0__pin_1_upper ) , 
    .chanx_left_in ( cbx_1__0__3_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_36_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_36_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_36_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_36_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_36_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_36_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_36_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_36_bottom_width_0_height_0__pin_49_lower ) , 
    .left_bottom_grid_pin_1_ ( grid_io_bottom_3_top_width_0_height_0__pin_1_lower ) , 
    .ccff_head ( grid_io_bottom_4_ccff_tail ) , 
    .chany_top_out ( sb_1__0__3_chany_top_out ) , 
    .chanx_right_out ( sb_1__0__3_chanx_right_out ) , 
    .chanx_left_out ( sb_1__0__3_chanx_left_out ) , 
    .ccff_tail ( sb_1__0__3_ccff_tail ) ) ;
sb_1__0_ sb_5__0_ (
    .prog_clk ( { ctsbuf_net_2342216 } ) ,
    .chany_top_in ( cby_1__1__48_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_48_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_48_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_48_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_48_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_48_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_48_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_48_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_48_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__0__5_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_60_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_60_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_60_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_60_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_60_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_60_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_60_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_60_bottom_width_0_height_0__pin_49_upper ) , 
    .right_bottom_grid_pin_1_ ( grid_io_bottom_5_top_width_0_height_0__pin_1_upper ) , 
    .chanx_left_in ( cbx_1__0__4_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_48_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_48_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_48_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_48_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_48_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_48_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_48_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_48_bottom_width_0_height_0__pin_49_lower ) , 
    .left_bottom_grid_pin_1_ ( grid_io_bottom_4_top_width_0_height_0__pin_1_lower ) , 
    .ccff_head ( grid_io_bottom_5_ccff_tail ) , 
    .chany_top_out ( sb_1__0__4_chany_top_out ) , 
    .chanx_right_out ( sb_1__0__4_chanx_right_out ) , 
    .chanx_left_out ( sb_1__0__4_chanx_left_out ) , 
    .ccff_tail ( sb_1__0__4_ccff_tail ) ) ;
sb_1__0_ sb_6__0_ (
    .prog_clk ( { ctsbuf_net_1892171 } ) ,
    .chany_top_in ( cby_1__1__60_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_60_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_60_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_60_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_60_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_60_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_60_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_60_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_60_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__0__6_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_72_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_72_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_72_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_72_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_72_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_72_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_72_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_72_bottom_width_0_height_0__pin_49_upper ) , 
    .right_bottom_grid_pin_1_ ( grid_io_bottom_6_top_width_0_height_0__pin_1_upper ) , 
    .chanx_left_in ( cbx_1__0__5_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_60_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_60_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_60_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_60_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_60_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_60_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_60_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_60_bottom_width_0_height_0__pin_49_lower ) , 
    .left_bottom_grid_pin_1_ ( grid_io_bottom_5_top_width_0_height_0__pin_1_lower ) , 
    .ccff_head ( grid_io_bottom_6_ccff_tail ) , 
    .chany_top_out ( sb_1__0__5_chany_top_out ) , 
    .chanx_right_out ( sb_1__0__5_chanx_right_out ) , 
    .chanx_left_out ( sb_1__0__5_chanx_left_out ) , 
    .ccff_tail ( sb_1__0__5_ccff_tail ) ) ;
sb_1__0_ sb_7__0_ (
    .prog_clk ( { ctsbuf_net_1492131 } ) ,
    .chany_top_in ( cby_1__1__72_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_72_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_72_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_72_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_72_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_72_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_72_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_72_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_72_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__0__7_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_84_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_84_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_84_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_84_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_84_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_84_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_84_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_84_bottom_width_0_height_0__pin_49_upper ) , 
    .right_bottom_grid_pin_1_ ( grid_io_bottom_7_top_width_0_height_0__pin_1_upper ) , 
    .chanx_left_in ( cbx_1__0__6_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_72_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_72_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_72_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_72_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_72_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_72_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_72_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_72_bottom_width_0_height_0__pin_49_lower ) , 
    .left_bottom_grid_pin_1_ ( grid_io_bottom_6_top_width_0_height_0__pin_1_lower ) , 
    .ccff_head ( grid_io_bottom_7_ccff_tail ) , 
    .chany_top_out ( sb_1__0__6_chany_top_out ) , 
    .chanx_right_out ( sb_1__0__6_chanx_right_out ) , 
    .chanx_left_out ( sb_1__0__6_chanx_left_out ) , 
    .ccff_tail ( sb_1__0__6_ccff_tail ) ) ;
sb_1__0_ sb_8__0_ (
    .prog_clk ( { ctsbuf_net_1162098 } ) ,
    .chany_top_in ( cby_1__1__84_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_84_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_84_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_84_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_84_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_84_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_84_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_84_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_84_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__0__8_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_96_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_96_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_96_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_96_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_96_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_96_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_96_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_96_bottom_width_0_height_0__pin_49_upper ) , 
    .right_bottom_grid_pin_1_ ( grid_io_bottom_8_top_width_0_height_0__pin_1_upper ) , 
    .chanx_left_in ( cbx_1__0__7_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_84_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_84_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_84_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_84_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_84_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_84_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_84_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_84_bottom_width_0_height_0__pin_49_lower ) , 
    .left_bottom_grid_pin_1_ ( grid_io_bottom_7_top_width_0_height_0__pin_1_lower ) , 
    .ccff_head ( grid_io_bottom_8_ccff_tail ) , 
    .chany_top_out ( sb_1__0__7_chany_top_out ) , 
    .chanx_right_out ( sb_1__0__7_chanx_right_out ) , 
    .chanx_left_out ( sb_1__0__7_chanx_left_out ) , 
    .ccff_tail ( sb_1__0__7_ccff_tail ) ) ;
sb_1__0_ sb_9__0_ (
    .prog_clk ( { ctsbuf_net_882070 } ) ,
    .chany_top_in ( cby_1__1__96_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_96_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_96_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_96_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_96_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_96_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_96_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_96_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_96_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__0__9_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_108_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_108_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_108_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_108_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_108_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_108_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_108_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_108_bottom_width_0_height_0__pin_49_upper ) , 
    .right_bottom_grid_pin_1_ ( grid_io_bottom_9_top_width_0_height_0__pin_1_upper ) , 
    .chanx_left_in ( cbx_1__0__8_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_96_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_96_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_96_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_96_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_96_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_96_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_96_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_96_bottom_width_0_height_0__pin_49_lower ) , 
    .left_bottom_grid_pin_1_ ( grid_io_bottom_8_top_width_0_height_0__pin_1_lower ) , 
    .ccff_head ( grid_io_bottom_9_ccff_tail ) , 
    .chany_top_out ( sb_1__0__8_chany_top_out ) , 
    .chanx_right_out ( sb_1__0__8_chanx_right_out ) , 
    .chanx_left_out ( sb_1__0__8_chanx_left_out ) , 
    .ccff_tail ( sb_1__0__8_ccff_tail ) ) ;
sb_1__0_ sb_10__0_ (
    .prog_clk ( { ctsbuf_net_672049 } ) ,
    .chany_top_in ( cby_1__1__108_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_108_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_108_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_108_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_108_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_108_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_108_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_108_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_108_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__0__10_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_120_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_120_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_120_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_120_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_120_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_120_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_120_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_120_bottom_width_0_height_0__pin_49_upper ) , 
    .right_bottom_grid_pin_1_ ( grid_io_bottom_10_top_width_0_height_0__pin_1_upper ) , 
    .chanx_left_in ( cbx_1__0__9_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_108_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_108_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_108_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_108_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_108_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_108_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_108_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_108_bottom_width_0_height_0__pin_49_lower ) , 
    .left_bottom_grid_pin_1_ ( grid_io_bottom_9_top_width_0_height_0__pin_1_lower ) , 
    .ccff_head ( grid_io_bottom_10_ccff_tail ) , 
    .chany_top_out ( sb_1__0__9_chany_top_out ) , 
    .chanx_right_out ( sb_1__0__9_chanx_right_out ) , 
    .chanx_left_out ( sb_1__0__9_chanx_left_out ) , 
    .ccff_tail ( sb_1__0__9_ccff_tail ) ) ;
sb_1__0_ sb_11__0_ (
    .prog_clk ( { ctsbuf_net_522034 } ) ,
    .chany_top_in ( cby_1__1__120_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_120_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_120_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_120_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_120_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_120_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_120_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_120_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_120_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__0__11_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_132_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_132_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_132_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_132_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_132_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_132_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_132_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_132_bottom_width_0_height_0__pin_49_upper ) , 
    .right_bottom_grid_pin_1_ ( grid_io_bottom_11_top_width_0_height_0__pin_1_upper ) , 
    .chanx_left_in ( cbx_1__0__10_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_120_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_120_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_120_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_120_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_120_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_120_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_120_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_120_bottom_width_0_height_0__pin_49_lower ) , 
    .left_bottom_grid_pin_1_ ( grid_io_bottom_10_top_width_0_height_0__pin_1_lower ) , 
    .ccff_head ( grid_io_bottom_11_ccff_tail ) , 
    .chany_top_out ( sb_1__0__10_chany_top_out ) , 
    .chanx_right_out ( sb_1__0__10_chanx_right_out ) , 
    .chanx_left_out ( sb_1__0__10_chanx_left_out ) , 
    .ccff_tail ( sb_1__0__10_ccff_tail ) ) ;
sb_1__1_ sb_1__1_ (
    .prog_clk ( { ctsbuf_net_4482430 } ) ,
    .chany_top_in ( cby_1__1__1_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_1_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_1_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_1_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_1_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_1_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_1_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_1_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_1_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__1__11_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_13_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_13_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_13_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_13_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_13_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_13_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_13_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_13_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_1__1__0_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_0_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_0_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_0_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_0_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_0_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_0_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_0_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_0_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__0_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_1_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_1_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_1_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_1_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_1_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_1_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_1_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_1_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( cbx_1__1__11_ccff_tail ) , 
    .chany_top_out ( sb_1__1__0_chany_top_out ) , 
    .chanx_right_out ( sb_1__1__0_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__1__0_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__1__0_chanx_left_out ) , 
    .ccff_tail ( sb_1__1__0_ccff_tail ) ) ;
sb_1__1_ sb_1__2_ (
    .prog_clk ( { ctsbuf_net_4892471 } ) ,
    .chany_top_in ( cby_1__1__2_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_2_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_2_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_2_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_2_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_2_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_2_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_2_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_2_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__1__12_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_14_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_14_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_14_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_14_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_14_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_14_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_14_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_14_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_1__1__1_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_1_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_1_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_1_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_1_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_1_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_1_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_1_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_1_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__1_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_2_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_2_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_2_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_2_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_2_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_2_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_2_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_2_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( cbx_1__1__12_ccff_tail ) , 
    .chany_top_out ( sb_1__1__1_chany_top_out ) , 
    .chanx_right_out ( sb_1__1__1_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__1__1_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__1__1_chanx_left_out ) , 
    .ccff_tail ( sb_1__1__1_ccff_tail ) ) ;
sb_1__1_ sb_1__3_ (
    .prog_clk ( { ctsbuf_net_5212503 } ) ,
    .chany_top_in ( cby_1__1__3_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_3_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_3_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_3_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_3_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_3_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_3_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_3_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_3_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__1__13_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_15_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_15_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_15_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_15_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_15_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_15_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_15_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_15_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_1__1__2_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_2_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_2_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_2_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_2_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_2_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_2_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_2_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_2_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__2_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_3_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_3_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_3_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_3_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_3_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_3_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_3_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_3_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( cbx_1__1__13_ccff_tail ) , 
    .chany_top_out ( sb_1__1__2_chany_top_out ) , 
    .chanx_right_out ( sb_1__1__2_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__1__2_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__1__2_chanx_left_out ) , 
    .ccff_tail ( sb_1__1__2_ccff_tail ) ) ;
sb_1__1_ sb_1__4_ (
    .prog_clk ( { ctsbuf_net_5482530 } ) ,
    .chany_top_in ( cby_1__1__4_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_4_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_4_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_4_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_4_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_4_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_4_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_4_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_4_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__1__14_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_16_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_16_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_16_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_16_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_16_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_16_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_16_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_16_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_1__1__3_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_3_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_3_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_3_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_3_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_3_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_3_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_3_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_3_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__3_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_4_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_4_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_4_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_4_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_4_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_4_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_4_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_4_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( cbx_1__1__14_ccff_tail ) , 
    .chany_top_out ( sb_1__1__3_chany_top_out ) , 
    .chanx_right_out ( sb_1__1__3_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__1__3_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__1__3_chanx_left_out ) , 
    .ccff_tail ( sb_1__1__3_ccff_tail ) ) ;
sb_1__1_ sb_1__5_ (
    .prog_clk ( { ctsbuf_net_5672549 } ) ,
    .chany_top_in ( cby_1__1__5_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_5_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_5_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_5_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_5_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_5_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_5_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_5_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_5_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__1__15_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_17_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_17_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_17_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_17_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_17_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_17_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_17_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_17_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_1__1__4_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_4_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_4_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_4_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_4_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_4_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_4_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_4_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_4_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__4_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_5_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_5_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_5_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_5_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_5_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_5_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_5_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_5_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( cbx_1__1__15_ccff_tail ) , 
    .chany_top_out ( sb_1__1__4_chany_top_out ) , 
    .chanx_right_out ( sb_1__1__4_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__1__4_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__1__4_chanx_left_out ) , 
    .ccff_tail ( sb_1__1__4_ccff_tail ) ) ;
sb_1__1_ sb_1__6_ (
    .prog_clk ( { ctsbuf_net_5792561 } ) ,
    .chany_top_in ( cby_1__1__6_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_6_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_6_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_6_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_6_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_6_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_6_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_6_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_6_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__1__16_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_18_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_18_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_18_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_18_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_18_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_18_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_18_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_18_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_1__1__5_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_5_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_5_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_5_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_5_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_5_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_5_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_5_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_5_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__5_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_6_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_6_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_6_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_6_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_6_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_6_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_6_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_6_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( cbx_1__1__16_ccff_tail ) , 
    .chany_top_out ( sb_1__1__5_chany_top_out ) , 
    .chanx_right_out ( sb_1__1__5_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__1__5_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__1__5_chanx_left_out ) , 
    .ccff_tail ( sb_1__1__5_ccff_tail ) ) ;
sb_1__1_ sb_1__7_ (
    .prog_clk ( { ctsbuf_net_5702552 } ) ,
    .chany_top_in ( cby_1__1__7_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_7_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_7_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_7_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_7_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_7_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_7_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_7_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_7_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__1__17_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_19_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_19_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_19_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_19_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_19_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_19_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_19_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_19_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_1__1__6_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_6_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_6_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_6_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_6_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_6_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_6_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_6_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_6_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__6_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_7_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_7_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_7_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_7_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_7_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_7_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_7_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_7_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( cbx_1__1__17_ccff_tail ) , 
    .chany_top_out ( sb_1__1__6_chany_top_out ) , 
    .chanx_right_out ( sb_1__1__6_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__1__6_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__1__6_chanx_left_out ) , 
    .ccff_tail ( sb_1__1__6_ccff_tail ) ) ;
sb_1__1_ sb_1__8_ (
    .prog_clk ( { ctsbuf_net_5522534 } ) ,
    .chany_top_in ( cby_1__1__8_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_8_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_8_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_8_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_8_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_8_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_8_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_8_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_8_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__1__18_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_20_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_20_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_20_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_20_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_20_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_20_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_20_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_20_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_1__1__7_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_7_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_7_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_7_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_7_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_7_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_7_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_7_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_7_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__7_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_8_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_8_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_8_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_8_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_8_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_8_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_8_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_8_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( cbx_1__1__18_ccff_tail ) , 
    .chany_top_out ( sb_1__1__7_chany_top_out ) , 
    .chanx_right_out ( sb_1__1__7_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__1__7_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__1__7_chanx_left_out ) , 
    .ccff_tail ( sb_1__1__7_ccff_tail ) ) ;
sb_1__1_ sb_1__9_ (
    .prog_clk ( { ctsbuf_net_5262508 } ) ,
    .chany_top_in ( cby_1__1__9_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_9_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_9_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_9_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_9_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_9_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_9_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_9_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_9_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__1__19_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_21_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_21_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_21_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_21_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_21_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_21_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_21_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_21_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_1__1__8_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_8_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_8_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_8_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_8_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_8_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_8_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_8_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_8_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__8_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_9_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_9_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_9_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_9_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_9_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_9_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_9_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_9_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( cbx_1__1__19_ccff_tail ) , 
    .chany_top_out ( sb_1__1__8_chany_top_out ) , 
    .chanx_right_out ( sb_1__1__8_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__1__8_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__1__8_chanx_left_out ) , 
    .ccff_tail ( sb_1__1__8_ccff_tail ) ) ;
sb_1__1_ sb_1__10_ (
    .prog_clk ( { ctsbuf_net_4952477 } ) ,
    .chany_top_in ( cby_1__1__10_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_10_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_10_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_10_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_10_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_10_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_10_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_10_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_10_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__1__20_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_22_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_22_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_22_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_22_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_22_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_22_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_22_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_22_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_1__1__9_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_9_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_9_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_9_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_9_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_9_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_9_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_9_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_9_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__9_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_10_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_10_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_10_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_10_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_10_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_10_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_10_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_10_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( cbx_1__1__20_ccff_tail ) , 
    .chany_top_out ( sb_1__1__9_chany_top_out ) , 
    .chanx_right_out ( sb_1__1__9_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__1__9_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__1__9_chanx_left_out ) , 
    .ccff_tail ( sb_1__1__9_ccff_tail ) ) ;
sb_1__1_ sb_1__11_ (
    .prog_clk ( { p_abuf19 } ) ,
    .chany_top_in ( cby_1__1__11_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_11_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_11_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_11_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_11_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_11_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_11_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_11_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_11_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__1__21_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_23_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_23_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_23_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_23_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_23_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_23_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_23_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_23_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_1__1__10_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_10_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_10_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_10_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_10_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_10_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_10_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_10_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_10_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__10_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_11_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_11_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_11_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_11_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_11_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_11_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_11_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_11_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( cbx_1__1__21_ccff_tail ) , 
    .chany_top_out ( sb_1__1__10_chany_top_out ) , 
    .chanx_right_out ( sb_1__1__10_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__1__10_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__1__10_chanx_left_out ) , 
    .ccff_tail ( sb_1__1__10_ccff_tail ) ) ;
sb_1__1_ sb_2__1_ (
    .prog_clk ( { ctsbuf_net_4042386 } ) ,
    .chany_top_in ( cby_1__1__13_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_13_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_13_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_13_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_13_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_13_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_13_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_13_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_13_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__1__22_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_25_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_25_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_25_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_25_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_25_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_25_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_25_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_25_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_1__1__12_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_12_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_12_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_12_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_12_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_12_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_12_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_12_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_12_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__11_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_13_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_13_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_13_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_13_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_13_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_13_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_13_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_13_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( cbx_1__1__22_ccff_tail ) , 
    .chany_top_out ( sb_1__1__11_chany_top_out ) , 
    .chanx_right_out ( sb_1__1__11_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__1__11_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__1__11_chanx_left_out ) , 
    .ccff_tail ( sb_1__1__11_ccff_tail ) ) ;
sb_1__1_ sb_2__2_ (
    .prog_clk ( { ctsbuf_net_4492431 } ) ,
    .chany_top_in ( cby_1__1__14_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_14_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_14_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_14_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_14_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_14_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_14_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_14_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_14_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__1__23_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_26_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_26_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_26_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_26_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_26_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_26_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_26_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_26_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_1__1__13_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_13_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_13_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_13_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_13_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_13_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_13_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_13_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_13_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__12_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_14_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_14_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_14_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_14_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_14_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_14_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_14_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_14_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( cbx_1__1__23_ccff_tail ) , 
    .chany_top_out ( sb_1__1__12_chany_top_out ) , 
    .chanx_right_out ( sb_1__1__12_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__1__12_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__1__12_chanx_left_out ) , 
    .ccff_tail ( sb_1__1__12_ccff_tail ) ) ;
sb_1__1_ sb_2__3_ (
    .prog_clk ( { ctsbuf_net_4902472 } ) ,
    .chany_top_in ( cby_1__1__15_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_15_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_15_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_15_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_15_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_15_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_15_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_15_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_15_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__1__24_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_27_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_27_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_27_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_27_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_27_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_27_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_27_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_27_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_1__1__14_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_14_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_14_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_14_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_14_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_14_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_14_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_14_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_14_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__13_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_15_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_15_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_15_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_15_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_15_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_15_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_15_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_15_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( cbx_1__1__24_ccff_tail ) , 
    .chany_top_out ( sb_1__1__13_chany_top_out ) , 
    .chanx_right_out ( sb_1__1__13_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__1__13_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__1__13_chanx_left_out ) , 
    .ccff_tail ( sb_1__1__13_ccff_tail ) ) ;
sb_1__1_ sb_2__4_ (
    .prog_clk ( { ctsbuf_net_5222504 } ) ,
    .chany_top_in ( cby_1__1__16_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_16_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_16_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_16_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_16_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_16_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_16_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_16_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_16_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__1__25_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_28_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_28_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_28_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_28_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_28_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_28_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_28_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_28_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_1__1__15_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_15_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_15_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_15_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_15_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_15_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_15_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_15_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_15_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__14_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_16_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_16_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_16_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_16_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_16_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_16_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_16_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_16_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( cbx_1__1__25_ccff_tail ) , 
    .chany_top_out ( sb_1__1__14_chany_top_out ) , 
    .chanx_right_out ( sb_1__1__14_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__1__14_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__1__14_chanx_left_out ) , 
    .ccff_tail ( sb_1__1__14_ccff_tail ) ) ;
sb_1__1_ sb_2__5_ (
    .prog_clk ( { ctsbuf_net_5492531 } ) ,
    .chany_top_in ( cby_1__1__17_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_17_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_17_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_17_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_17_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_17_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_17_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_17_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_17_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__1__26_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_29_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_29_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_29_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_29_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_29_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_29_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_29_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_29_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_1__1__16_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_16_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_16_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_16_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_16_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_16_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_16_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_16_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_16_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__15_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_17_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_17_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_17_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_17_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_17_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_17_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_17_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_17_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( cbx_1__1__26_ccff_tail ) , 
    .chany_top_out ( sb_1__1__15_chany_top_out ) , 
    .chanx_right_out ( sb_1__1__15_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__1__15_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__1__15_chanx_left_out ) , 
    .ccff_tail ( sb_1__1__15_ccff_tail ) ) ;
sb_1__1_ sb_2__6_ (
    .prog_clk ( { ctsbuf_net_5682550 } ) ,
    .chany_top_in ( cby_1__1__18_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_18_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_18_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_18_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_18_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_18_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_18_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_18_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_18_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__1__27_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_30_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_30_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_30_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_30_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_30_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_30_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_30_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_30_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_1__1__17_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_17_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_17_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_17_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_17_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_17_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_17_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_17_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_17_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__16_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_18_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_18_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_18_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_18_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_18_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_18_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_18_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_18_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( cbx_1__1__27_ccff_tail ) , 
    .chany_top_out ( sb_1__1__16_chany_top_out ) , 
    .chanx_right_out ( sb_1__1__16_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__1__16_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__1__16_chanx_left_out ) , 
    .ccff_tail ( sb_1__1__16_ccff_tail ) ) ;
sb_1__1_ sb_2__7_ (
    .prog_clk ( { ctsbuf_net_5532535 } ) ,
    .chany_top_in ( cby_1__1__19_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_19_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_19_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_19_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_19_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_19_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_19_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_19_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_19_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__1__28_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_31_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_31_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_31_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_31_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_31_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_31_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_31_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_31_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_1__1__18_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_18_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_18_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_18_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_18_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_18_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_18_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_18_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_18_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__17_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_19_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_19_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_19_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_19_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_19_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_19_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_19_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_19_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( cbx_1__1__28_ccff_tail ) , 
    .chany_top_out ( sb_1__1__17_chany_top_out ) , 
    .chanx_right_out ( sb_1__1__17_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__1__17_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__1__17_chanx_left_out ) , 
    .ccff_tail ( sb_1__1__17_ccff_tail ) ) ;
sb_1__1_ sb_2__8_ (
    .prog_clk ( { ctsbuf_net_5272509 } ) ,
    .chany_top_in ( cby_1__1__20_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_20_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_20_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_20_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_20_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_20_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_20_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_20_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_20_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__1__29_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_32_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_32_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_32_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_32_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_32_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_32_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_32_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_32_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_1__1__19_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_19_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_19_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_19_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_19_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_19_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_19_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_19_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_19_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__18_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_20_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_20_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_20_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_20_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_20_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_20_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_20_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_20_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( cbx_1__1__29_ccff_tail ) , 
    .chany_top_out ( sb_1__1__18_chany_top_out ) , 
    .chanx_right_out ( sb_1__1__18_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__1__18_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__1__18_chanx_left_out ) , 
    .ccff_tail ( sb_1__1__18_ccff_tail ) ) ;
sb_1__1_ sb_2__9_ (
    .prog_clk ( { ctsbuf_net_4962478 } ) ,
    .chany_top_in ( cby_1__1__21_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_21_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_21_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_21_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_21_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_21_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_21_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_21_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_21_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__1__30_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_33_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_33_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_33_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_33_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_33_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_33_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_33_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_33_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_1__1__20_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_20_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_20_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_20_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_20_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_20_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_20_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_20_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_20_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__19_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_21_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_21_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_21_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_21_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_21_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_21_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_21_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_21_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( cbx_1__1__30_ccff_tail ) , 
    .chany_top_out ( sb_1__1__19_chany_top_out ) , 
    .chanx_right_out ( sb_1__1__19_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__1__19_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__1__19_chanx_left_out ) , 
    .ccff_tail ( sb_1__1__19_ccff_tail ) ) ;
sb_1__1_ sb_2__10_ (
    .prog_clk ( { ctsbuf_net_4562438 } ) ,
    .chany_top_in ( cby_1__1__22_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_22_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_22_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_22_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_22_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_22_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_22_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_22_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_22_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__1__31_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_34_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_34_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_34_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_34_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_34_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_34_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_34_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_34_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_1__1__21_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_21_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_21_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_21_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_21_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_21_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_21_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_21_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_21_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__20_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_22_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_22_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_22_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_22_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_22_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_22_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_22_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_22_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( cbx_1__1__31_ccff_tail ) , 
    .chany_top_out ( sb_1__1__20_chany_top_out ) , 
    .chanx_right_out ( sb_1__1__20_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__1__20_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__1__20_chanx_left_out ) , 
    .ccff_tail ( sb_1__1__20_ccff_tail ) ) ;
sb_1__1_ sb_2__11_ (
    .prog_clk ( { ctsbuf_net_4102392 } ) ,
    .chany_top_in ( cby_1__1__23_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_23_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_23_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_23_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_23_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_23_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_23_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_23_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_23_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__1__32_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_35_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_35_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_35_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_35_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_35_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_35_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_35_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_35_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_1__1__22_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_22_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_22_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_22_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_22_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_22_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_22_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_22_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_22_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__21_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_23_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_23_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_23_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_23_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_23_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_23_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_23_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_23_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( cbx_1__1__32_ccff_tail ) , 
    .chany_top_out ( sb_1__1__21_chany_top_out ) , 
    .chanx_right_out ( sb_1__1__21_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__1__21_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__1__21_chanx_left_out ) , 
    .ccff_tail ( sb_1__1__21_ccff_tail ) ) ;
sb_1__1_ sb_3__1_ (
    .prog_clk ( { ctsbuf_net_3612343 } ) ,
    .chany_top_in ( cby_1__1__25_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_25_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_25_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_25_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_25_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_25_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_25_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_25_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_25_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__1__33_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_37_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_37_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_37_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_37_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_37_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_37_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_37_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_37_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_1__1__24_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_24_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_24_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_24_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_24_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_24_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_24_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_24_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_24_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__22_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_25_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_25_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_25_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_25_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_25_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_25_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_25_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_25_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( cbx_1__1__33_ccff_tail ) , 
    .chany_top_out ( sb_1__1__22_chany_top_out ) , 
    .chanx_right_out ( sb_1__1__22_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__1__22_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__1__22_chanx_left_out ) , 
    .ccff_tail ( sb_1__1__22_ccff_tail ) ) ;
sb_1__1_ sb_3__2_ (
    .prog_clk ( { ctsbuf_net_4052387 } ) ,
    .chany_top_in ( cby_1__1__26_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_26_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_26_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_26_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_26_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_26_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_26_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_26_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_26_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__1__34_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_38_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_38_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_38_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_38_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_38_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_38_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_38_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_38_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_1__1__25_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_25_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_25_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_25_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_25_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_25_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_25_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_25_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_25_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__23_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_26_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_26_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_26_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_26_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_26_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_26_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_26_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_26_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( cbx_1__1__34_ccff_tail ) , 
    .chany_top_out ( sb_1__1__23_chany_top_out ) , 
    .chanx_right_out ( sb_1__1__23_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__1__23_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__1__23_chanx_left_out ) , 
    .ccff_tail ( sb_1__1__23_ccff_tail ) ) ;
sb_1__1_ sb_3__3_ (
    .prog_clk ( { p_abuf18 } ) ,
    .chany_top_in ( cby_1__1__27_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_27_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_27_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_27_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_27_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_27_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_27_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_27_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_27_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__1__35_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_39_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_39_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_39_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_39_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_39_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_39_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_39_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_39_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_1__1__26_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_26_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_26_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_26_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_26_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_26_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_26_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_26_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_26_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__24_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_27_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_27_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_27_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_27_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_27_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_27_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_27_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_27_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( cbx_1__1__35_ccff_tail ) , 
    .chany_top_out ( sb_1__1__24_chany_top_out ) , 
    .chanx_right_out ( sb_1__1__24_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__1__24_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__1__24_chanx_left_out ) , 
    .ccff_tail ( sb_1__1__24_ccff_tail ) ) ;
sb_1__1_ sb_3__4_ (
    .prog_clk ( { ctsbuf_net_4912473 } ) ,
    .chany_top_in ( cby_1__1__28_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_28_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_28_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_28_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_28_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_28_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_28_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_28_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_28_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__1__36_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_40_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_40_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_40_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_40_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_40_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_40_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_40_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_40_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_1__1__27_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_27_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_27_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_27_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_27_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_27_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_27_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_27_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_27_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__25_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_28_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_28_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_28_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_28_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_28_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_28_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_28_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_28_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( cbx_1__1__36_ccff_tail ) , 
    .chany_top_out ( sb_1__1__25_chany_top_out ) , 
    .chanx_right_out ( sb_1__1__25_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__1__25_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__1__25_chanx_left_out ) , 
    .ccff_tail ( sb_1__1__25_ccff_tail ) ) ;
sb_1__1_ sb_3__5_ (
    .prog_clk ( { ctsbuf_net_5232505 } ) ,
    .chany_top_in ( cby_1__1__29_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_29_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_29_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_29_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_29_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_29_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_29_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_29_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_29_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__1__37_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_41_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_41_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_41_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_41_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_41_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_41_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_41_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_41_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_1__1__28_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_28_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_28_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_28_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_28_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_28_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_28_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_28_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_28_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__26_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_29_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_29_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_29_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_29_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_29_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_29_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_29_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_29_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( cbx_1__1__37_ccff_tail ) , 
    .chany_top_out ( sb_1__1__26_chany_top_out ) , 
    .chanx_right_out ( sb_1__1__26_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__1__26_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__1__26_chanx_left_out ) , 
    .ccff_tail ( sb_1__1__26_ccff_tail ) ) ;
sb_1__1_ sb_3__6_ (
    .prog_clk ( { ctsbuf_net_5502532 } ) ,
    .chany_top_in ( cby_1__1__30_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_30_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_30_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_30_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_30_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_30_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_30_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_30_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_30_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__1__38_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_42_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_42_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_42_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_42_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_42_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_42_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_42_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_42_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_1__1__29_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_29_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_29_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_29_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_29_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_29_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_29_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_29_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_29_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__27_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_30_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_30_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_30_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_30_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_30_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_30_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_30_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_30_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( cbx_1__1__38_ccff_tail ) , 
    .chany_top_out ( sb_1__1__27_chany_top_out ) , 
    .chanx_right_out ( sb_1__1__27_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__1__27_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__1__27_chanx_left_out ) , 
    .ccff_tail ( sb_1__1__27_ccff_tail ) ) ;
sb_1__1_ sb_3__7_ (
    .prog_clk ( { ctsbuf_net_5282510 } ) ,
    .chany_top_in ( cby_1__1__31_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_31_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_31_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_31_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_31_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_31_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_31_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_31_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_31_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__1__39_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_43_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_43_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_43_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_43_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_43_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_43_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_43_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_43_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_1__1__30_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_30_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_30_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_30_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_30_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_30_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_30_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_30_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_30_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__28_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_31_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_31_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_31_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_31_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_31_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_31_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_31_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_31_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( cbx_1__1__39_ccff_tail ) , 
    .chany_top_out ( sb_1__1__28_chany_top_out ) , 
    .chanx_right_out ( sb_1__1__28_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__1__28_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__1__28_chanx_left_out ) , 
    .ccff_tail ( sb_1__1__28_ccff_tail ) ) ;
sb_1__1_ sb_3__8_ (
    .prog_clk ( { ctsbuf_net_4972479 } ) ,
    .chany_top_in ( cby_1__1__32_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_32_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_32_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_32_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_32_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_32_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_32_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_32_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_32_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__1__40_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_44_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_44_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_44_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_44_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_44_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_44_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_44_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_44_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_1__1__31_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_31_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_31_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_31_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_31_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_31_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_31_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_31_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_31_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__29_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_32_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_32_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_32_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_32_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_32_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_32_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_32_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_32_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( cbx_1__1__40_ccff_tail ) , 
    .chany_top_out ( sb_1__1__29_chany_top_out ) , 
    .chanx_right_out ( sb_1__1__29_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__1__29_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__1__29_chanx_left_out ) , 
    .ccff_tail ( sb_1__1__29_ccff_tail ) ) ;
sb_1__1_ sb_3__9_ (
    .prog_clk ( { ctsbuf_net_4572439 } ) ,
    .chany_top_in ( cby_1__1__33_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_33_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_33_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_33_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_33_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_33_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_33_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_33_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_33_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__1__41_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_45_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_45_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_45_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_45_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_45_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_45_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_45_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_45_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_1__1__32_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_32_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_32_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_32_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_32_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_32_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_32_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_32_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_32_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__30_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_33_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_33_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_33_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_33_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_33_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_33_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_33_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_33_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( cbx_1__1__41_ccff_tail ) , 
    .chany_top_out ( sb_1__1__30_chany_top_out ) , 
    .chanx_right_out ( sb_1__1__30_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__1__30_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__1__30_chanx_left_out ) , 
    .ccff_tail ( sb_1__1__30_ccff_tail ) ) ;
sb_1__1_ sb_3__10_ (
    .prog_clk ( { ctsbuf_net_4122394 } ) ,
    .chany_top_in ( cby_1__1__34_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_34_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_34_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_34_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_34_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_34_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_34_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_34_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_34_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__1__42_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_46_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_46_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_46_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_46_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_46_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_46_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_46_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_46_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_1__1__33_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_33_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_33_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_33_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_33_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_33_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_33_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_33_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_33_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__31_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_34_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_34_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_34_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_34_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_34_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_34_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_34_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_34_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( cbx_1__1__42_ccff_tail ) , 
    .chany_top_out ( sb_1__1__31_chany_top_out ) , 
    .chanx_right_out ( sb_1__1__31_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__1__31_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__1__31_chanx_left_out ) , 
    .ccff_tail ( sb_1__1__31_ccff_tail ) ) ;
sb_1__1_ sb_3__11_ (
    .prog_clk ( { ctsbuf_net_3672349 } ) ,
    .chany_top_in ( cby_1__1__35_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_35_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_35_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_35_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_35_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_35_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_35_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_35_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_35_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__1__43_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_47_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_47_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_47_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_47_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_47_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_47_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_47_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_47_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_1__1__34_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_34_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_34_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_34_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_34_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_34_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_34_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_34_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_34_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__32_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_35_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_35_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_35_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_35_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_35_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_35_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_35_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_35_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( cbx_1__1__43_ccff_tail ) , 
    .chany_top_out ( sb_1__1__32_chany_top_out ) , 
    .chanx_right_out ( sb_1__1__32_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__1__32_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__1__32_chanx_left_out ) , 
    .ccff_tail ( sb_1__1__32_ccff_tail ) ) ;
sb_1__1_ sb_4__1_ (
    .prog_clk ( { ctsbuf_net_3172299 } ) ,
    .chany_top_in ( cby_1__1__37_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_37_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_37_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_37_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_37_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_37_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_37_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_37_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_37_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__1__44_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_49_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_49_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_49_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_49_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_49_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_49_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_49_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_49_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_1__1__36_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_36_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_36_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_36_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_36_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_36_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_36_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_36_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_36_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__33_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_37_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_37_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_37_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_37_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_37_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_37_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_37_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_37_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( cbx_1__1__44_ccff_tail ) , 
    .chany_top_out ( sb_1__1__33_chany_top_out ) , 
    .chanx_right_out ( sb_1__1__33_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__1__33_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__1__33_chanx_left_out ) , 
    .ccff_tail ( sb_1__1__33_ccff_tail ) ) ;
sb_1__1_ sb_4__2_ (
    .prog_clk ( { ctsbuf_net_3622344 } ) ,
    .chany_top_in ( cby_1__1__38_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_38_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_38_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_38_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_38_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_38_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_38_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_38_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_38_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__1__45_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_50_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_50_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_50_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_50_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_50_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_50_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_50_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_50_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_1__1__37_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_37_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_37_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_37_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_37_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_37_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_37_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_37_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_37_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__34_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_38_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_38_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_38_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_38_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_38_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_38_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_38_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_38_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( cbx_1__1__45_ccff_tail ) , 
    .chany_top_out ( sb_1__1__34_chany_top_out ) , 
    .chanx_right_out ( sb_1__1__34_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__1__34_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__1__34_chanx_left_out ) , 
    .ccff_tail ( sb_1__1__34_ccff_tail ) ) ;
sb_1__1_ sb_4__3_ (
    .prog_clk ( { ctsbuf_net_4062388 } ) ,
    .chany_top_in ( cby_1__1__39_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_39_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_39_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_39_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_39_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_39_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_39_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_39_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_39_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__1__46_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_51_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_51_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_51_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_51_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_51_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_51_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_51_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_51_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_1__1__38_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_38_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_38_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_38_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_38_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_38_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_38_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_38_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_38_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__35_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_39_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_39_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_39_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_39_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_39_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_39_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_39_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_39_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( cbx_1__1__46_ccff_tail ) , 
    .chany_top_out ( sb_1__1__35_chany_top_out ) , 
    .chanx_right_out ( sb_1__1__35_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__1__35_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__1__35_chanx_left_out ) , 
    .ccff_tail ( sb_1__1__35_ccff_tail ) ) ;
sb_1__1_ sb_4__4_ (
    .prog_clk ( { ctsbuf_net_4512433 } ) ,
    .chany_top_in ( cby_1__1__40_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_40_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_40_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_40_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_40_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_40_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_40_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_40_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_40_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__1__47_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_52_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_52_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_52_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_52_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_52_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_52_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_52_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_52_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_1__1__39_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_39_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_39_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_39_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_39_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_39_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_39_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_39_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_39_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__36_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_40_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_40_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_40_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_40_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_40_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_40_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_40_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_40_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( cbx_1__1__47_ccff_tail ) , 
    .chany_top_out ( sb_1__1__36_chany_top_out ) , 
    .chanx_right_out ( sb_1__1__36_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__1__36_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__1__36_chanx_left_out ) , 
    .ccff_tail ( sb_1__1__36_ccff_tail ) ) ;
sb_1__1_ sb_4__5_ (
    .prog_clk ( { ctsbuf_net_4922474 } ) ,
    .chany_top_in ( cby_1__1__41_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_41_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_41_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_41_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_41_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_41_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_41_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_41_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_41_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__1__48_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_53_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_53_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_53_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_53_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_53_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_53_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_53_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_53_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_1__1__40_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_40_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_40_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_40_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_40_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_40_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_40_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_40_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_40_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__37_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_41_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_41_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_41_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_41_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_41_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_41_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_41_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_41_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( cbx_1__1__48_ccff_tail ) , 
    .chany_top_out ( sb_1__1__37_chany_top_out ) , 
    .chanx_right_out ( sb_1__1__37_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__1__37_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__1__37_chanx_left_out ) , 
    .ccff_tail ( sb_1__1__37_ccff_tail ) ) ;
sb_1__1_ sb_4__6_ (
    .prog_clk ( { ctsbuf_net_5242506 } ) ,
    .chany_top_in ( cby_1__1__42_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_42_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_42_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_42_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_42_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_42_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_42_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_42_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_42_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__1__49_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_54_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_54_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_54_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_54_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_54_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_54_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_54_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_54_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_1__1__41_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_41_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_41_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_41_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_41_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_41_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_41_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_41_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_41_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__38_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_42_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_42_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_42_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_42_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_42_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_42_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_42_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_42_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( cbx_1__1__49_ccff_tail ) , 
    .chany_top_out ( sb_1__1__38_chany_top_out ) , 
    .chanx_right_out ( sb_1__1__38_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__1__38_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__1__38_chanx_left_out ) , 
    .ccff_tail ( sb_1__1__38_ccff_tail ) ) ;
sb_1__1_ sb_4__7_ (
    .prog_clk ( { ctsbuf_net_4982480 } ) ,
    .chany_top_in ( cby_1__1__43_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_43_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_43_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_43_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_43_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_43_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_43_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_43_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_43_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__1__50_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_55_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_55_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_55_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_55_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_55_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_55_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_55_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_55_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_1__1__42_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_42_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_42_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_42_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_42_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_42_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_42_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_42_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_42_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__39_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_43_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_43_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_43_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_43_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_43_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_43_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_43_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_43_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( cbx_1__1__50_ccff_tail ) , 
    .chany_top_out ( sb_1__1__39_chany_top_out ) , 
    .chanx_right_out ( sb_1__1__39_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__1__39_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__1__39_chanx_left_out ) , 
    .ccff_tail ( sb_1__1__39_ccff_tail ) ) ;
sb_1__1_ sb_4__8_ (
    .prog_clk ( { ctsbuf_net_4582440 } ) ,
    .chany_top_in ( cby_1__1__44_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_44_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_44_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_44_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_44_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_44_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_44_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_44_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_44_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__1__51_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_56_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_56_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_56_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_56_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_56_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_56_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_56_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_56_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_1__1__43_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_43_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_43_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_43_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_43_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_43_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_43_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_43_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_43_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__40_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_44_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_44_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_44_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_44_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_44_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_44_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_44_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_44_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( cbx_1__1__51_ccff_tail ) , 
    .chany_top_out ( sb_1__1__40_chany_top_out ) , 
    .chanx_right_out ( sb_1__1__40_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__1__40_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__1__40_chanx_left_out ) , 
    .ccff_tail ( sb_1__1__40_ccff_tail ) ) ;
sb_1__1_ sb_4__9_ (
    .prog_clk ( { ctsbuf_net_4132395 } ) ,
    .chany_top_in ( cby_1__1__45_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_45_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_45_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_45_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_45_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_45_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_45_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_45_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_45_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__1__52_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_57_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_57_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_57_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_57_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_57_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_57_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_57_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_57_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_1__1__44_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_44_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_44_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_44_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_44_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_44_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_44_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_44_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_44_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__41_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_45_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_45_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_45_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_45_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_45_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_45_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_45_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_45_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( cbx_1__1__52_ccff_tail ) , 
    .chany_top_out ( sb_1__1__41_chany_top_out ) , 
    .chanx_right_out ( sb_1__1__41_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__1__41_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__1__41_chanx_left_out ) , 
    .ccff_tail ( sb_1__1__41_ccff_tail ) ) ;
sb_1__1_ sb_4__10_ (
    .prog_clk ( { ctsbuf_net_3692351 } ) ,
    .chany_top_in ( cby_1__1__46_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_46_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_46_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_46_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_46_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_46_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_46_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_46_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_46_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__1__53_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_58_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_58_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_58_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_58_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_58_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_58_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_58_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_58_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_1__1__45_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_45_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_45_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_45_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_45_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_45_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_45_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_45_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_45_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__42_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_46_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_46_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_46_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_46_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_46_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_46_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_46_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_46_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( cbx_1__1__53_ccff_tail ) , 
    .chany_top_out ( sb_1__1__42_chany_top_out ) , 
    .chanx_right_out ( sb_1__1__42_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__1__42_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__1__42_chanx_left_out ) , 
    .ccff_tail ( sb_1__1__42_ccff_tail ) ) ;
sb_1__1_ sb_4__11_ (
    .prog_clk ( { ctsbuf_net_3232305 } ) ,
    .chany_top_in ( cby_1__1__47_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_47_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_47_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_47_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_47_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_47_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_47_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_47_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_47_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__1__54_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_59_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_59_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_59_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_59_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_59_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_59_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_59_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_59_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_1__1__46_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_46_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_46_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_46_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_46_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_46_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_46_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_46_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_46_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__43_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_47_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_47_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_47_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_47_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_47_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_47_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_47_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_47_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( cbx_1__1__54_ccff_tail ) , 
    .chany_top_out ( sb_1__1__43_chany_top_out ) , 
    .chanx_right_out ( sb_1__1__43_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__1__43_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__1__43_chanx_left_out ) , 
    .ccff_tail ( sb_1__1__43_ccff_tail ) ) ;
sb_1__1_ sb_5__1_ (
    .prog_clk ( { ctsbuf_net_2722254 } ) ,
    .chany_top_in ( cby_1__1__49_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_49_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_49_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_49_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_49_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_49_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_49_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_49_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_49_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__1__55_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_61_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_61_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_61_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_61_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_61_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_61_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_61_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_61_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_1__1__48_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_48_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_48_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_48_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_48_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_48_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_48_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_48_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_48_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__44_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_49_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_49_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_49_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_49_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_49_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_49_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_49_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_49_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( cbx_1__1__55_ccff_tail ) , 
    .chany_top_out ( sb_1__1__44_chany_top_out ) , 
    .chanx_right_out ( sb_1__1__44_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__1__44_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__1__44_chanx_left_out ) , 
    .ccff_tail ( sb_1__1__44_ccff_tail ) ) ;
sb_1__1_ sb_5__2_ (
    .prog_clk ( { ctsbuf_net_3182300 } ) ,
    .chany_top_in ( cby_1__1__50_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_50_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_50_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_50_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_50_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_50_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_50_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_50_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_50_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__1__56_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_62_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_62_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_62_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_62_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_62_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_62_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_62_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_62_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_1__1__49_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_49_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_49_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_49_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_49_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_49_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_49_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_49_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_49_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__45_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_50_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_50_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_50_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_50_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_50_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_50_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_50_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_50_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( cbx_1__1__56_ccff_tail ) , 
    .chany_top_out ( sb_1__1__45_chany_top_out ) , 
    .chanx_right_out ( sb_1__1__45_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__1__45_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__1__45_chanx_left_out ) , 
    .ccff_tail ( sb_1__1__45_ccff_tail ) ) ;
sb_1__1_ sb_5__3_ (
    .prog_clk ( { ctsbuf_net_3632345 } ) ,
    .chany_top_in ( cby_1__1__51_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_51_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_51_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_51_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_51_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_51_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_51_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_51_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_51_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__1__57_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_63_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_63_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_63_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_63_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_63_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_63_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_63_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_63_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_1__1__50_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_50_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_50_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_50_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_50_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_50_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_50_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_50_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_50_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__46_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_51_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_51_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_51_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_51_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_51_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_51_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_51_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_51_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( cbx_1__1__57_ccff_tail ) , 
    .chany_top_out ( sb_1__1__46_chany_top_out ) , 
    .chanx_right_out ( sb_1__1__46_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__1__46_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__1__46_chanx_left_out ) , 
    .ccff_tail ( sb_1__1__46_ccff_tail ) ) ;
sb_1__1_ sb_5__4_ (
    .prog_clk ( { ctsbuf_net_4072389 } ) ,
    .chany_top_in ( cby_1__1__52_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_52_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_52_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_52_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_52_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_52_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_52_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_52_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_52_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__1__58_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_64_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_64_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_64_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_64_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_64_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_64_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_64_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_64_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_1__1__51_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_51_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_51_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_51_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_51_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_51_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_51_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_51_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_51_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__47_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_52_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_52_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_52_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_52_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_52_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_52_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_52_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_52_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( cbx_1__1__58_ccff_tail ) , 
    .chany_top_out ( sb_1__1__47_chany_top_out ) , 
    .chanx_right_out ( sb_1__1__47_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__1__47_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__1__47_chanx_left_out ) , 
    .ccff_tail ( sb_1__1__47_ccff_tail ) ) ;
sb_1__1_ sb_5__5_ (
    .prog_clk ( { ctsbuf_net_4522434 } ) ,
    .chany_top_in ( cby_1__1__53_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_53_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_53_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_53_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_53_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_53_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_53_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_53_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_53_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__1__59_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_65_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_65_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_65_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_65_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_65_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_65_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_65_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_65_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_1__1__52_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_52_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_52_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_52_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_52_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_52_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_52_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_52_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_52_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__48_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_53_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_53_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_53_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_53_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_53_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_53_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_53_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_53_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( cbx_1__1__59_ccff_tail ) , 
    .chany_top_out ( sb_1__1__48_chany_top_out ) , 
    .chanx_right_out ( sb_1__1__48_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__1__48_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__1__48_chanx_left_out ) , 
    .ccff_tail ( sb_1__1__48_ccff_tail ) ) ;
sb_1__1_ sb_5__6_ (
    .prog_clk ( { ctsbuf_net_4932475 } ) ,
    .chany_top_in ( cby_1__1__54_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_54_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_54_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_54_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_54_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_54_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_54_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_54_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_54_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__1__60_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_66_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_66_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_66_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_66_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_66_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_66_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_66_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_66_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_1__1__53_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_53_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_53_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_53_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_53_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_53_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_53_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_53_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_53_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__49_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_54_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_54_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_54_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_54_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_54_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_54_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_54_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_54_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( cbx_1__1__60_ccff_tail ) , 
    .chany_top_out ( sb_1__1__49_chany_top_out ) , 
    .chanx_right_out ( sb_1__1__49_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__1__49_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__1__49_chanx_left_out ) , 
    .ccff_tail ( sb_1__1__49_ccff_tail ) ) ;
sb_1__1_ sb_5__7_ (
    .prog_clk ( { ctsbuf_net_4592441 } ) ,
    .chany_top_in ( cby_1__1__55_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_55_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_55_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_55_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_55_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_55_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_55_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_55_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_55_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__1__61_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_67_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_67_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_67_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_67_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_67_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_67_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_67_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_67_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_1__1__54_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_54_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_54_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_54_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_54_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_54_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_54_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_54_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_54_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__50_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_55_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_55_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_55_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_55_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_55_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_55_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_55_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_55_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( cbx_1__1__61_ccff_tail ) , 
    .chany_top_out ( sb_1__1__50_chany_top_out ) , 
    .chanx_right_out ( sb_1__1__50_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__1__50_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__1__50_chanx_left_out ) , 
    .ccff_tail ( sb_1__1__50_ccff_tail ) ) ;
sb_1__1_ sb_5__8_ (
    .prog_clk ( { ctsbuf_net_4142396 } ) ,
    .chany_top_in ( cby_1__1__56_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_56_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_56_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_56_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_56_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_56_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_56_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_56_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_56_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__1__62_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_68_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_68_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_68_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_68_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_68_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_68_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_68_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_68_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_1__1__55_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_55_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_55_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_55_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_55_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_55_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_55_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_55_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_55_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__51_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_56_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_56_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_56_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_56_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_56_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_56_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_56_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_56_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( cbx_1__1__62_ccff_tail ) , 
    .chany_top_out ( sb_1__1__51_chany_top_out ) , 
    .chanx_right_out ( sb_1__1__51_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__1__51_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__1__51_chanx_left_out ) , 
    .ccff_tail ( sb_1__1__51_ccff_tail ) ) ;
sb_1__1_ sb_5__9_ (
    .prog_clk ( { ctsbuf_net_3702352 } ) ,
    .chany_top_in ( cby_1__1__57_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_57_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_57_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_57_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_57_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_57_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_57_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_57_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_57_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__1__63_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_69_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_69_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_69_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_69_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_69_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_69_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_69_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_69_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_1__1__56_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_56_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_56_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_56_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_56_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_56_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_56_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_56_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_56_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__52_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_57_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_57_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_57_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_57_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_57_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_57_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_57_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_57_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( cbx_1__1__63_ccff_tail ) , 
    .chany_top_out ( sb_1__1__52_chany_top_out ) , 
    .chanx_right_out ( sb_1__1__52_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__1__52_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__1__52_chanx_left_out ) , 
    .ccff_tail ( sb_1__1__52_ccff_tail ) ) ;
sb_1__1_ sb_5__10_ (
    .prog_clk ( { ctsbuf_net_3252307 } ) ,
    .chany_top_in ( cby_1__1__58_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_58_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_58_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_58_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_58_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_58_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_58_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_58_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_58_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__1__64_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_70_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_70_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_70_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_70_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_70_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_70_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_70_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_70_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_1__1__57_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_57_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_57_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_57_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_57_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_57_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_57_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_57_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_57_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__53_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_58_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_58_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_58_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_58_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_58_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_58_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_58_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_58_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( cbx_1__1__64_ccff_tail ) , 
    .chany_top_out ( sb_1__1__53_chany_top_out ) , 
    .chanx_right_out ( sb_1__1__53_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__1__53_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__1__53_chanx_left_out ) , 
    .ccff_tail ( sb_1__1__53_ccff_tail ) ) ;
sb_1__1_ sb_5__11_ (
    .prog_clk ( { ctsbuf_net_2782260 } ) ,
    .chany_top_in ( cby_1__1__59_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_59_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_59_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_59_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_59_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_59_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_59_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_59_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_59_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__1__65_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_71_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_71_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_71_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_71_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_71_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_71_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_71_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_71_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_1__1__58_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_58_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_58_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_58_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_58_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_58_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_58_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_58_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_58_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__54_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_59_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_59_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_59_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_59_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_59_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_59_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_59_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_59_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( cbx_1__1__65_ccff_tail ) , 
    .chany_top_out ( sb_1__1__54_chany_top_out ) , 
    .chanx_right_out ( sb_1__1__54_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__1__54_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__1__54_chanx_left_out ) , 
    .ccff_tail ( sb_1__1__54_ccff_tail ) ) ;
sb_1__1_ sb_6__1_ (
    .prog_clk ( { ctsbuf_net_2272209 } ) ,
    .chany_top_in ( cby_1__1__61_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_61_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_61_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_61_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_61_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_61_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_61_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_61_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_61_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__1__66_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_73_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_73_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_73_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_73_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_73_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_73_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_73_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_73_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_1__1__60_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_60_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_60_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_60_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_60_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_60_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_60_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_60_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_60_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__55_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_61_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_61_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_61_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_61_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_61_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_61_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_61_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_61_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( cbx_1__1__66_ccff_tail ) , 
    .chany_top_out ( sb_1__1__55_chany_top_out ) , 
    .chanx_right_out ( sb_1__1__55_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__1__55_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__1__55_chanx_left_out ) , 
    .ccff_tail ( sb_1__1__55_ccff_tail ) ) ;
sb_1__1_ sb_6__2_ (
    .prog_clk ( { ctsbuf_net_2732255 } ) ,
    .chany_top_in ( cby_1__1__62_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_62_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_62_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_62_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_62_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_62_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_62_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_62_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_62_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__1__67_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_74_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_74_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_74_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_74_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_74_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_74_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_74_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_74_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_1__1__61_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_61_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_61_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_61_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_61_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_61_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_61_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_61_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_61_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__56_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_62_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_62_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_62_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_62_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_62_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_62_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_62_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_62_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( cbx_1__1__67_ccff_tail ) , 
    .chany_top_out ( sb_1__1__56_chany_top_out ) , 
    .chanx_right_out ( sb_1__1__56_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__1__56_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__1__56_chanx_left_out ) , 
    .ccff_tail ( sb_1__1__56_ccff_tail ) ) ;
sb_1__1_ sb_6__3_ (
    .prog_clk ( { ctsbuf_net_3192301 } ) ,
    .chany_top_in ( cby_1__1__63_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_63_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_63_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_63_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_63_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_63_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_63_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_63_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_63_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__1__68_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_75_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_75_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_75_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_75_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_75_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_75_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_75_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_75_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_1__1__62_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_62_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_62_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_62_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_62_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_62_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_62_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_62_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_62_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__57_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_63_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_63_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_63_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_63_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_63_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_63_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_63_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_63_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( cbx_1__1__68_ccff_tail ) , 
    .chany_top_out ( sb_1__1__57_chany_top_out ) , 
    .chanx_right_out ( sb_1__1__57_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__1__57_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__1__57_chanx_left_out ) , 
    .ccff_tail ( sb_1__1__57_ccff_tail ) ) ;
sb_1__1_ sb_6__4_ (
    .prog_clk ( { ctsbuf_net_3642346 } ) ,
    .chany_top_in ( cby_1__1__64_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_64_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_64_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_64_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_64_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_64_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_64_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_64_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_64_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__1__69_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_76_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_76_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_76_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_76_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_76_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_76_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_76_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_76_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_1__1__63_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_63_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_63_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_63_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_63_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_63_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_63_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_63_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_63_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__58_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_64_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_64_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_64_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_64_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_64_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_64_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_64_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_64_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( cbx_1__1__69_ccff_tail ) , 
    .chany_top_out ( sb_1__1__58_chany_top_out ) , 
    .chanx_right_out ( sb_1__1__58_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__1__58_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__1__58_chanx_left_out ) , 
    .ccff_tail ( sb_1__1__58_ccff_tail ) ) ;
sb_1__1_ sb_6__5_ (
    .prog_clk ( { ctsbuf_net_4082390 } ) ,
    .chany_top_in ( cby_1__1__65_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_65_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_65_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_65_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_65_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_65_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_65_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_65_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_65_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__1__70_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_77_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_77_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_77_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_77_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_77_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_77_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_77_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_77_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_1__1__64_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_64_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_64_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_64_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_64_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_64_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_64_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_64_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_64_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__59_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_65_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_65_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_65_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_65_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_65_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_65_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_65_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_65_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( cbx_1__1__70_ccff_tail ) , 
    .chany_top_out ( sb_1__1__59_chany_top_out ) , 
    .chanx_right_out ( sb_1__1__59_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__1__59_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__1__59_chanx_left_out ) , 
    .ccff_tail ( sb_1__1__59_ccff_tail ) ) ;
sb_1__1_ sb_6__6_ (
    .prog_clk ( { ctsbuf_net_4532435 } ) ,
    .chany_top_in ( cby_1__1__66_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_66_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_66_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_66_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_66_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_66_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_66_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_66_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_66_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__1__71_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_78_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_78_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_78_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_78_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_78_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_78_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_78_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_78_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_1__1__65_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_65_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_65_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_65_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_65_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_65_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_65_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_65_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_65_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__60_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_66_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_66_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_66_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_66_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_66_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_66_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_66_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_66_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( cbx_1__1__71_ccff_tail ) , 
    .chany_top_out ( sb_1__1__60_chany_top_out ) , 
    .chanx_right_out ( sb_1__1__60_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__1__60_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__1__60_chanx_left_out ) , 
    .ccff_tail ( sb_1__1__60_ccff_tail ) ) ;
sb_1__1_ sb_6__7_ (
    .prog_clk ( { ctsbuf_net_4152397 } ) ,
    .chany_top_in ( cby_1__1__67_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_67_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_67_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_67_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_67_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_67_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_67_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_67_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_67_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__1__72_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_79_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_79_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_79_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_79_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_79_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_79_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_79_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_79_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_1__1__66_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_66_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_66_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_66_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_66_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_66_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_66_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_66_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_66_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__61_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_67_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_67_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_67_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_67_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_67_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_67_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_67_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_67_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( cbx_1__1__72_ccff_tail ) , 
    .chany_top_out ( sb_1__1__61_chany_top_out ) , 
    .chanx_right_out ( sb_1__1__61_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__1__61_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__1__61_chanx_left_out ) , 
    .ccff_tail ( sb_1__1__61_ccff_tail ) ) ;
sb_1__1_ sb_6__8_ (
    .prog_clk ( { ctsbuf_net_3712353 } ) ,
    .chany_top_in ( cby_1__1__68_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_68_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_68_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_68_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_68_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_68_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_68_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_68_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_68_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__1__73_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_80_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_80_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_80_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_80_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_80_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_80_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_80_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_80_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_1__1__67_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_67_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_67_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_67_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_67_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_67_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_67_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_67_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_67_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__62_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_68_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_68_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_68_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_68_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_68_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_68_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_68_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_68_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( cbx_1__1__73_ccff_tail ) , 
    .chany_top_out ( sb_1__1__62_chany_top_out ) , 
    .chanx_right_out ( sb_1__1__62_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__1__62_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__1__62_chanx_left_out ) , 
    .ccff_tail ( sb_1__1__62_ccff_tail ) ) ;
sb_1__1_ sb_6__9_ (
    .prog_clk ( { ctsbuf_net_3262308 } ) ,
    .chany_top_in ( cby_1__1__69_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_69_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_69_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_69_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_69_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_69_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_69_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_69_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_69_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__1__74_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_81_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_81_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_81_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_81_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_81_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_81_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_81_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_81_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_1__1__68_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_68_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_68_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_68_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_68_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_68_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_68_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_68_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_68_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__63_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_69_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_69_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_69_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_69_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_69_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_69_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_69_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_69_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( cbx_1__1__74_ccff_tail ) , 
    .chany_top_out ( sb_1__1__63_chany_top_out ) , 
    .chanx_right_out ( sb_1__1__63_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__1__63_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__1__63_chanx_left_out ) , 
    .ccff_tail ( sb_1__1__63_ccff_tail ) ) ;
sb_1__1_ sb_6__10_ (
    .prog_clk ( { ctsbuf_net_2802262 } ) ,
    .chany_top_in ( cby_1__1__70_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_70_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_70_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_70_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_70_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_70_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_70_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_70_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_70_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__1__75_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_82_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_82_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_82_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_82_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_82_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_82_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_82_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_82_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_1__1__69_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_69_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_69_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_69_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_69_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_69_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_69_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_69_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_69_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__64_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_70_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_70_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_70_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_70_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_70_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_70_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_70_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_70_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( cbx_1__1__75_ccff_tail ) , 
    .chany_top_out ( sb_1__1__64_chany_top_out ) , 
    .chanx_right_out ( sb_1__1__64_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__1__64_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__1__64_chanx_left_out ) , 
    .ccff_tail ( sb_1__1__64_ccff_tail ) ) ;
sb_1__1_ sb_6__11_ (
    .prog_clk ( { ctsbuf_net_2332215 } ) ,
    .chany_top_in ( cby_1__1__71_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_71_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_71_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_71_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_71_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_71_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_71_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_71_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_71_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__1__76_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_83_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_83_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_83_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_83_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_83_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_83_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_83_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_83_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_1__1__70_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_70_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_70_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_70_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_70_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_70_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_70_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_70_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_70_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__65_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_71_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_71_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_71_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_71_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_71_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_71_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_71_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_71_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( cbx_1__1__76_ccff_tail ) , 
    .chany_top_out ( sb_1__1__65_chany_top_out ) , 
    .chanx_right_out ( sb_1__1__65_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__1__65_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__1__65_chanx_left_out ) , 
    .ccff_tail ( sb_1__1__65_ccff_tail ) ) ;
sb_1__1_ sb_7__1_ (
    .prog_clk ( { ctsbuf_net_1832165 } ) ,
    .chany_top_in ( cby_1__1__73_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_73_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_73_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_73_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_73_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_73_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_73_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_73_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_73_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__1__77_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_85_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_85_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_85_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_85_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_85_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_85_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_85_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_85_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_1__1__72_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_72_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_72_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_72_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_72_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_72_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_72_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_72_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_72_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__66_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_73_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_73_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_73_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_73_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_73_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_73_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_73_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_73_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( cbx_1__1__77_ccff_tail ) , 
    .chany_top_out ( sb_1__1__66_chany_top_out ) , 
    .chanx_right_out ( sb_1__1__66_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__1__66_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__1__66_chanx_left_out ) , 
    .ccff_tail ( sb_1__1__66_ccff_tail ) ) ;
sb_1__1_ sb_7__2_ (
    .prog_clk ( { ctsbuf_net_2282210 } ) ,
    .chany_top_in ( cby_1__1__74_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_74_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_74_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_74_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_74_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_74_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_74_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_74_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_74_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__1__78_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_86_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_86_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_86_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_86_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_86_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_86_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_86_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_86_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_1__1__73_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_73_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_73_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_73_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_73_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_73_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_73_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_73_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_73_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__67_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_74_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_74_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_74_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_74_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_74_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_74_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_74_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_74_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( cbx_1__1__78_ccff_tail ) , 
    .chany_top_out ( sb_1__1__67_chany_top_out ) , 
    .chanx_right_out ( sb_1__1__67_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__1__67_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__1__67_chanx_left_out ) , 
    .ccff_tail ( sb_1__1__67_ccff_tail ) ) ;
sb_1__1_ sb_7__3_ (
    .prog_clk ( { ctsbuf_net_2742256 } ) ,
    .chany_top_in ( cby_1__1__75_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_75_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_75_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_75_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_75_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_75_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_75_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_75_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_75_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__1__79_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_87_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_87_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_87_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_87_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_87_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_87_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_87_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_87_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_1__1__74_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_74_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_74_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_74_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_74_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_74_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_74_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_74_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_74_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__68_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_75_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_75_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_75_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_75_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_75_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_75_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_75_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_75_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( cbx_1__1__79_ccff_tail ) , 
    .chany_top_out ( sb_1__1__68_chany_top_out ) , 
    .chanx_right_out ( sb_1__1__68_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__1__68_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__1__68_chanx_left_out ) , 
    .ccff_tail ( sb_1__1__68_ccff_tail ) ) ;
sb_1__1_ sb_7__4_ (
    .prog_clk ( { ctsbuf_net_3202302 } ) ,
    .chany_top_in ( cby_1__1__76_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_76_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_76_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_76_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_76_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_76_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_76_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_76_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_76_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__1__80_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_88_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_88_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_88_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_88_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_88_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_88_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_88_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_88_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_1__1__75_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_75_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_75_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_75_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_75_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_75_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_75_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_75_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_75_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__69_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_76_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_76_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_76_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_76_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_76_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_76_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_76_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_76_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( cbx_1__1__80_ccff_tail ) , 
    .chany_top_out ( sb_1__1__69_chany_top_out ) , 
    .chanx_right_out ( sb_1__1__69_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__1__69_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__1__69_chanx_left_out ) , 
    .ccff_tail ( sb_1__1__69_ccff_tail ) ) ;
sb_1__1_ sb_7__5_ (
    .prog_clk ( { ctsbuf_net_3652347 } ) ,
    .chany_top_in ( cby_1__1__77_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_77_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_77_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_77_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_77_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_77_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_77_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_77_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_77_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__1__81_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_89_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_89_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_89_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_89_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_89_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_89_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_89_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_89_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_1__1__76_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_76_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_76_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_76_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_76_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_76_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_76_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_76_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_76_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__70_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_77_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_77_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_77_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_77_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_77_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_77_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_77_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_77_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( cbx_1__1__81_ccff_tail ) , 
    .chany_top_out ( sb_1__1__70_chany_top_out ) , 
    .chanx_right_out ( sb_1__1__70_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__1__70_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__1__70_chanx_left_out ) , 
    .ccff_tail ( sb_1__1__70_ccff_tail ) ) ;
sb_1__1_ sb_7__6_ (
    .prog_clk ( { ctsbuf_net_4092391 } ) ,
    .chany_top_in ( cby_1__1__78_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_78_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_78_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_78_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_78_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_78_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_78_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_78_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_78_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__1__82_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_90_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_90_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_90_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_90_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_90_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_90_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_90_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_90_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_1__1__77_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_77_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_77_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_77_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_77_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_77_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_77_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_77_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_77_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__71_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_78_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_78_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_78_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_78_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_78_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_78_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_78_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_78_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( cbx_1__1__82_ccff_tail ) , 
    .chany_top_out ( sb_1__1__71_chany_top_out ) , 
    .chanx_right_out ( sb_1__1__71_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__1__71_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__1__71_chanx_left_out ) , 
    .ccff_tail ( sb_1__1__71_ccff_tail ) ) ;
sb_1__1_ sb_7__7_ (
    .prog_clk ( { ctsbuf_net_3722354 } ) ,
    .chany_top_in ( cby_1__1__79_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_79_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_79_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_79_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_79_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_79_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_79_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_79_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_79_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__1__83_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_91_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_91_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_91_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_91_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_91_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_91_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_91_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_91_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_1__1__78_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_78_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_78_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_78_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_78_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_78_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_78_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_78_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_78_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__72_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_79_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_79_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_79_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_79_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_79_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_79_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_79_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_79_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( cbx_1__1__83_ccff_tail ) , 
    .chany_top_out ( sb_1__1__72_chany_top_out ) , 
    .chanx_right_out ( sb_1__1__72_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__1__72_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__1__72_chanx_left_out ) , 
    .ccff_tail ( sb_1__1__72_ccff_tail ) ) ;
sb_1__1_ sb_7__8_ (
    .prog_clk ( { ctsbuf_net_3272309 } ) ,
    .chany_top_in ( cby_1__1__80_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_80_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_80_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_80_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_80_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_80_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_80_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_80_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_80_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__1__84_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_92_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_92_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_92_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_92_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_92_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_92_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_92_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_92_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_1__1__79_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_79_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_79_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_79_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_79_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_79_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_79_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_79_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_79_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__73_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_80_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_80_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_80_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_80_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_80_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_80_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_80_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_80_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( cbx_1__1__84_ccff_tail ) , 
    .chany_top_out ( sb_1__1__73_chany_top_out ) , 
    .chanx_right_out ( sb_1__1__73_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__1__73_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__1__73_chanx_left_out ) , 
    .ccff_tail ( sb_1__1__73_ccff_tail ) ) ;
sb_1__1_ sb_7__9_ (
    .prog_clk ( { ctsbuf_net_2812263 } ) ,
    .chany_top_in ( cby_1__1__81_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_81_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_81_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_81_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_81_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_81_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_81_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_81_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_81_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__1__85_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_93_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_93_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_93_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_93_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_93_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_93_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_93_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_93_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_1__1__80_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_80_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_80_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_80_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_80_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_80_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_80_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_80_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_80_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__74_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_81_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_81_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_81_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_81_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_81_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_81_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_81_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_81_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( cbx_1__1__85_ccff_tail ) , 
    .chany_top_out ( sb_1__1__74_chany_top_out ) , 
    .chanx_right_out ( sb_1__1__74_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__1__74_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__1__74_chanx_left_out ) , 
    .ccff_tail ( sb_1__1__74_ccff_tail ) ) ;
sb_1__1_ sb_7__10_ (
    .prog_clk ( { ctsbuf_net_2352217 } ) ,
    .chany_top_in ( cby_1__1__82_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_82_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_82_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_82_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_82_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_82_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_82_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_82_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_82_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__1__86_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_94_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_94_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_94_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_94_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_94_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_94_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_94_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_94_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_1__1__81_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_81_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_81_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_81_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_81_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_81_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_81_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_81_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_81_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__75_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_82_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_82_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_82_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_82_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_82_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_82_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_82_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_82_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( cbx_1__1__86_ccff_tail ) , 
    .chany_top_out ( sb_1__1__75_chany_top_out ) , 
    .chanx_right_out ( sb_1__1__75_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__1__75_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__1__75_chanx_left_out ) , 
    .ccff_tail ( sb_1__1__75_ccff_tail ) ) ;
sb_1__1_ sb_7__11_ (
    .prog_clk ( { ctsbuf_net_1882170 } ) ,
    .chany_top_in ( cby_1__1__83_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_83_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_83_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_83_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_83_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_83_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_83_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_83_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_83_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__1__87_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_95_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_95_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_95_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_95_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_95_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_95_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_95_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_95_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_1__1__82_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_82_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_82_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_82_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_82_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_82_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_82_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_82_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_82_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__76_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_83_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_83_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_83_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_83_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_83_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_83_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_83_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_83_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( cbx_1__1__87_ccff_tail ) , 
    .chany_top_out ( sb_1__1__76_chany_top_out ) , 
    .chanx_right_out ( sb_1__1__76_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__1__76_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__1__76_chanx_left_out ) , 
    .ccff_tail ( sb_1__1__76_ccff_tail ) ) ;
sb_1__1_ sb_8__1_ (
    .prog_clk ( { ctsbuf_net_1442126 } ) ,
    .chany_top_in ( cby_1__1__85_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_85_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_85_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_85_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_85_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_85_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_85_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_85_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_85_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__1__88_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_97_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_97_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_97_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_97_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_97_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_97_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_97_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_97_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_1__1__84_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_84_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_84_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_84_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_84_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_84_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_84_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_84_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_84_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__77_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_85_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_85_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_85_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_85_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_85_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_85_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_85_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_85_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( cbx_1__1__88_ccff_tail ) , 
    .chany_top_out ( sb_1__1__77_chany_top_out ) , 
    .chanx_right_out ( sb_1__1__77_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__1__77_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__1__77_chanx_left_out ) , 
    .ccff_tail ( sb_1__1__77_ccff_tail ) ) ;
sb_1__1_ sb_8__2_ (
    .prog_clk ( { ctsbuf_net_1842166 } ) ,
    .chany_top_in ( cby_1__1__86_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_86_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_86_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_86_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_86_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_86_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_86_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_86_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_86_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__1__89_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_98_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_98_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_98_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_98_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_98_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_98_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_98_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_98_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_1__1__85_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_85_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_85_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_85_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_85_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_85_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_85_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_85_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_85_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__78_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_86_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_86_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_86_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_86_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_86_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_86_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_86_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_86_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( cbx_1__1__89_ccff_tail ) , 
    .chany_top_out ( sb_1__1__78_chany_top_out ) , 
    .chanx_right_out ( sb_1__1__78_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__1__78_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__1__78_chanx_left_out ) , 
    .ccff_tail ( sb_1__1__78_ccff_tail ) ) ;
sb_1__1_ sb_8__3_ (
    .prog_clk ( { ctsbuf_net_2292211 } ) ,
    .chany_top_in ( cby_1__1__87_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_87_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_87_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_87_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_87_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_87_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_87_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_87_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_87_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__1__90_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_99_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_99_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_99_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_99_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_99_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_99_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_99_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_99_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_1__1__86_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_86_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_86_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_86_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_86_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_86_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_86_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_86_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_86_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__79_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_87_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_87_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_87_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_87_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_87_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_87_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_87_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_87_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( cbx_1__1__90_ccff_tail ) , 
    .chany_top_out ( sb_1__1__79_chany_top_out ) , 
    .chanx_right_out ( sb_1__1__79_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__1__79_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__1__79_chanx_left_out ) , 
    .ccff_tail ( sb_1__1__79_ccff_tail ) ) ;
sb_1__1_ sb_8__4_ (
    .prog_clk ( { ctsbuf_net_2752257 } ) ,
    .chany_top_in ( cby_1__1__88_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_88_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_88_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_88_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_88_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_88_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_88_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_88_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_88_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__1__91_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_100_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_100_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_100_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_100_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_100_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_100_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_100_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_100_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_1__1__87_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_87_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_87_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_87_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_87_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_87_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_87_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_87_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_87_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__80_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_88_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_88_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_88_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_88_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_88_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_88_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_88_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_88_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( cbx_1__1__91_ccff_tail ) , 
    .chany_top_out ( sb_1__1__80_chany_top_out ) , 
    .chanx_right_out ( sb_1__1__80_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__1__80_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__1__80_chanx_left_out ) , 
    .ccff_tail ( sb_1__1__80_ccff_tail ) ) ;
sb_1__1_ sb_8__5_ (
    .prog_clk ( { ctsbuf_net_3212303 } ) ,
    .chany_top_in ( cby_1__1__89_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_89_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_89_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_89_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_89_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_89_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_89_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_89_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_89_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__1__92_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_101_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_101_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_101_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_101_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_101_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_101_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_101_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_101_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_1__1__88_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_88_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_88_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_88_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_88_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_88_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_88_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_88_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_88_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__81_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_89_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_89_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_89_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_89_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_89_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_89_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_89_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_89_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( cbx_1__1__92_ccff_tail ) , 
    .chany_top_out ( sb_1__1__81_chany_top_out ) , 
    .chanx_right_out ( sb_1__1__81_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__1__81_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__1__81_chanx_left_out ) , 
    .ccff_tail ( sb_1__1__81_ccff_tail ) ) ;
sb_1__1_ sb_8__6_ (
    .prog_clk ( { ctsbuf_net_3662348 } ) ,
    .chany_top_in ( cby_1__1__90_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_90_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_90_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_90_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_90_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_90_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_90_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_90_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_90_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__1__93_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_102_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_102_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_102_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_102_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_102_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_102_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_102_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_102_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_1__1__89_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_89_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_89_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_89_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_89_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_89_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_89_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_89_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_89_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__82_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_90_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_90_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_90_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_90_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_90_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_90_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_90_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_90_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( cbx_1__1__93_ccff_tail ) , 
    .chany_top_out ( sb_1__1__82_chany_top_out ) , 
    .chanx_right_out ( sb_1__1__82_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__1__82_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__1__82_chanx_left_out ) , 
    .ccff_tail ( sb_1__1__82_ccff_tail ) ) ;
sb_1__1_ sb_8__7_ (
    .prog_clk ( { ctsbuf_net_3282310 } ) ,
    .chany_top_in ( cby_1__1__91_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_91_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_91_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_91_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_91_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_91_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_91_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_91_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_91_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__1__94_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_103_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_103_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_103_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_103_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_103_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_103_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_103_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_103_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_1__1__90_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_90_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_90_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_90_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_90_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_90_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_90_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_90_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_90_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__83_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_91_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_91_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_91_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_91_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_91_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_91_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_91_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_91_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( cbx_1__1__94_ccff_tail ) , 
    .chany_top_out ( sb_1__1__83_chany_top_out ) , 
    .chanx_right_out ( sb_1__1__83_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__1__83_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__1__83_chanx_left_out ) , 
    .ccff_tail ( sb_1__1__83_ccff_tail ) ) ;
sb_1__1_ sb_8__8_ (
    .prog_clk ( { ctsbuf_net_2822264 } ) ,
    .chany_top_in ( cby_1__1__92_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_92_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_92_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_92_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_92_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_92_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_92_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_92_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_92_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__1__95_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_104_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_104_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_104_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_104_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_104_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_104_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_104_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_104_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_1__1__91_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_91_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_91_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_91_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_91_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_91_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_91_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_91_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_91_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__84_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_92_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_92_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_92_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_92_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_92_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_92_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_92_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_92_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( cbx_1__1__95_ccff_tail ) , 
    .chany_top_out ( sb_1__1__84_chany_top_out ) , 
    .chanx_right_out ( sb_1__1__84_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__1__84_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__1__84_chanx_left_out ) , 
    .ccff_tail ( sb_1__1__84_ccff_tail ) ) ;
sb_1__1_ sb_8__9_ (
    .prog_clk ( { ctsbuf_net_2362218 } ) ,
    .chany_top_in ( cby_1__1__93_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_93_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_93_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_93_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_93_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_93_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_93_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_93_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_93_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__1__96_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_105_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_105_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_105_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_105_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_105_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_105_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_105_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_105_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_1__1__92_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_92_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_92_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_92_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_92_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_92_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_92_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_92_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_92_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__85_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_93_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_93_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_93_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_93_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_93_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_93_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_93_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_93_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( cbx_1__1__96_ccff_tail ) , 
    .chany_top_out ( sb_1__1__85_chany_top_out ) , 
    .chanx_right_out ( sb_1__1__85_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__1__85_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__1__85_chanx_left_out ) , 
    .ccff_tail ( sb_1__1__85_ccff_tail ) ) ;
sb_1__1_ sb_8__10_ (
    .prog_clk ( { ctsbuf_net_1902172 } ) ,
    .chany_top_in ( cby_1__1__94_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_94_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_94_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_94_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_94_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_94_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_94_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_94_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_94_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__1__97_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_106_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_106_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_106_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_106_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_106_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_106_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_106_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_106_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_1__1__93_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_93_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_93_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_93_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_93_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_93_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_93_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_93_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_93_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__86_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_94_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_94_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_94_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_94_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_94_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_94_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_94_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_94_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( cbx_1__1__97_ccff_tail ) , 
    .chany_top_out ( sb_1__1__86_chany_top_out ) , 
    .chanx_right_out ( sb_1__1__86_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__1__86_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__1__86_chanx_left_out ) , 
    .ccff_tail ( sb_1__1__86_ccff_tail ) ) ;
sb_1__1_ sb_8__11_ (
    .prog_clk ( { ctsbuf_net_1482130 } ) ,
    .chany_top_in ( cby_1__1__95_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_95_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_95_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_95_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_95_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_95_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_95_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_95_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_95_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__1__98_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_107_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_107_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_107_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_107_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_107_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_107_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_107_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_107_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_1__1__94_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_94_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_94_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_94_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_94_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_94_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_94_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_94_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_94_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__87_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_95_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_95_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_95_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_95_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_95_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_95_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_95_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_95_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( cbx_1__1__98_ccff_tail ) , 
    .chany_top_out ( sb_1__1__87_chany_top_out ) , 
    .chanx_right_out ( sb_1__1__87_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__1__87_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__1__87_chanx_left_out ) , 
    .ccff_tail ( sb_1__1__87_ccff_tail ) ) ;
sb_1__1_ sb_9__1_ (
    .prog_clk ( { ctsbuf_net_1122094 } ) ,
    .chany_top_in ( cby_1__1__97_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_97_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_97_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_97_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_97_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_97_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_97_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_97_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_97_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__1__99_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_109_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_109_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_109_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_109_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_109_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_109_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_109_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_109_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_1__1__96_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_96_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_96_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_96_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_96_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_96_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_96_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_96_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_96_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__88_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_97_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_97_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_97_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_97_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_97_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_97_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_97_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_97_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( cbx_1__1__99_ccff_tail ) , 
    .chany_top_out ( sb_1__1__88_chany_top_out ) , 
    .chanx_right_out ( sb_1__1__88_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__1__88_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__1__88_chanx_left_out ) , 
    .ccff_tail ( sb_1__1__88_ccff_tail ) ) ;
sb_1__1_ sb_9__2_ (
    .prog_clk ( { ctsbuf_net_1452127 } ) ,
    .chany_top_in ( cby_1__1__98_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_98_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_98_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_98_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_98_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_98_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_98_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_98_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_98_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__1__100_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_110_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_110_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_110_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_110_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_110_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_110_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_110_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_110_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_1__1__97_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_97_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_97_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_97_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_97_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_97_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_97_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_97_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_97_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__89_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_98_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_98_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_98_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_98_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_98_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_98_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_98_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_98_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( cbx_1__1__100_ccff_tail ) , 
    .chany_top_out ( sb_1__1__89_chany_top_out ) , 
    .chanx_right_out ( sb_1__1__89_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__1__89_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__1__89_chanx_left_out ) , 
    .ccff_tail ( sb_1__1__89_ccff_tail ) ) ;
sb_1__1_ sb_9__3_ (
    .prog_clk ( { ctsbuf_net_1852167 } ) ,
    .chany_top_in ( cby_1__1__99_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_99_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_99_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_99_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_99_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_99_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_99_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_99_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_99_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__1__101_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_111_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_111_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_111_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_111_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_111_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_111_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_111_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_111_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_1__1__98_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_98_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_98_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_98_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_98_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_98_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_98_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_98_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_98_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__90_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_99_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_99_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_99_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_99_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_99_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_99_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_99_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_99_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( cbx_1__1__101_ccff_tail ) , 
    .chany_top_out ( sb_1__1__90_chany_top_out ) , 
    .chanx_right_out ( sb_1__1__90_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__1__90_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__1__90_chanx_left_out ) , 
    .ccff_tail ( sb_1__1__90_ccff_tail ) ) ;
sb_1__1_ sb_9__4_ (
    .prog_clk ( { ctsbuf_net_2302212 } ) ,
    .chany_top_in ( cby_1__1__100_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_100_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_100_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_100_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_100_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_100_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_100_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_100_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_100_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__1__102_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_112_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_112_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_112_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_112_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_112_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_112_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_112_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_112_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_1__1__99_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_99_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_99_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_99_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_99_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_99_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_99_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_99_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_99_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__91_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_100_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_100_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_100_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_100_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_100_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_100_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_100_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_100_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( cbx_1__1__102_ccff_tail ) , 
    .chany_top_out ( sb_1__1__91_chany_top_out ) , 
    .chanx_right_out ( sb_1__1__91_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__1__91_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__1__91_chanx_left_out ) , 
    .ccff_tail ( sb_1__1__91_ccff_tail ) ) ;
sb_1__1_ sb_9__5_ (
    .prog_clk ( { ctsbuf_net_2762258 } ) ,
    .chany_top_in ( cby_1__1__101_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_101_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_101_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_101_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_101_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_101_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_101_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_101_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_101_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__1__103_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_113_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_113_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_113_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_113_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_113_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_113_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_113_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_113_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_1__1__100_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_100_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_100_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_100_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_100_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_100_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_100_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_100_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_100_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__92_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_101_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_101_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_101_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_101_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_101_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_101_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_101_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_101_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( cbx_1__1__103_ccff_tail ) , 
    .chany_top_out ( sb_1__1__92_chany_top_out ) , 
    .chanx_right_out ( sb_1__1__92_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__1__92_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__1__92_chanx_left_out ) , 
    .ccff_tail ( sb_1__1__92_ccff_tail ) ) ;
sb_1__1_ sb_9__6_ (
    .prog_clk ( { ctsbuf_net_3222304 } ) ,
    .chany_top_in ( cby_1__1__102_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_102_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_102_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_102_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_102_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_102_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_102_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_102_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_102_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__1__104_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_114_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_114_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_114_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_114_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_114_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_114_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_114_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_114_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_1__1__101_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_101_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_101_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_101_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_101_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_101_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_101_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_101_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_101_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__93_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_102_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_102_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_102_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_102_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_102_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_102_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_102_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_102_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( cbx_1__1__104_ccff_tail ) , 
    .chany_top_out ( sb_1__1__93_chany_top_out ) , 
    .chanx_right_out ( sb_1__1__93_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__1__93_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__1__93_chanx_left_out ) , 
    .ccff_tail ( sb_1__1__93_ccff_tail ) ) ;
sb_1__1_ sb_9__7_ (
    .prog_clk ( { ctsbuf_net_2832265 } ) ,
    .chany_top_in ( cby_1__1__103_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_103_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_103_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_103_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_103_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_103_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_103_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_103_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_103_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__1__105_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_115_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_115_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_115_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_115_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_115_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_115_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_115_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_115_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_1__1__102_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_102_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_102_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_102_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_102_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_102_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_102_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_102_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_102_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__94_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_103_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_103_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_103_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_103_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_103_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_103_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_103_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_103_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( cbx_1__1__105_ccff_tail ) , 
    .chany_top_out ( sb_1__1__94_chany_top_out ) , 
    .chanx_right_out ( sb_1__1__94_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__1__94_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__1__94_chanx_left_out ) , 
    .ccff_tail ( sb_1__1__94_ccff_tail ) ) ;
sb_1__1_ sb_9__8_ (
    .prog_clk ( { p_abuf11 } ) ,
    .chany_top_in ( cby_1__1__104_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_104_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_104_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_104_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_104_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_104_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_104_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_104_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_104_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__1__106_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_116_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_116_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_116_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_116_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_116_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_116_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_116_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_116_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_1__1__103_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_103_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_103_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_103_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_103_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_103_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_103_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_103_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_103_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__95_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_104_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_104_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_104_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_104_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_104_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_104_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_104_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_104_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( cbx_1__1__106_ccff_tail ) , 
    .chany_top_out ( sb_1__1__95_chany_top_out ) , 
    .chanx_right_out ( sb_1__1__95_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__1__95_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__1__95_chanx_left_out ) , 
    .ccff_tail ( sb_1__1__95_ccff_tail ) ) ;
sb_1__1_ sb_9__9_ (
    .prog_clk ( { ctsbuf_net_1912173 } ) ,
    .chany_top_in ( cby_1__1__105_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_105_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_105_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_105_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_105_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_105_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_105_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_105_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_105_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__1__107_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_117_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_117_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_117_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_117_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_117_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_117_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_117_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_117_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_1__1__104_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_104_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_104_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_104_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_104_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_104_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_104_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_104_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_104_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__96_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_105_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_105_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_105_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_105_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_105_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_105_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_105_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_105_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( cbx_1__1__107_ccff_tail ) , 
    .chany_top_out ( sb_1__1__96_chany_top_out ) , 
    .chanx_right_out ( sb_1__1__96_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__1__96_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__1__96_chanx_left_out ) , 
    .ccff_tail ( sb_1__1__96_ccff_tail ) ) ;
sb_1__1_ sb_9__10_ (
    .prog_clk ( { ctsbuf_net_1502132 } ) ,
    .chany_top_in ( cby_1__1__106_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_106_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_106_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_106_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_106_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_106_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_106_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_106_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_106_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__1__108_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_118_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_118_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_118_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_118_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_118_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_118_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_118_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_118_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_1__1__105_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_105_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_105_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_105_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_105_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_105_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_105_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_105_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_105_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__97_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_106_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_106_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_106_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_106_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_106_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_106_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_106_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_106_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( cbx_1__1__108_ccff_tail ) , 
    .chany_top_out ( sb_1__1__97_chany_top_out ) , 
    .chanx_right_out ( sb_1__1__97_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__1__97_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__1__97_chanx_left_out ) , 
    .ccff_tail ( sb_1__1__97_ccff_tail ) ) ;
sb_1__1_ sb_9__11_ (
    .prog_clk ( { ctsbuf_net_1152097 } ) ,
    .chany_top_in ( cby_1__1__107_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_107_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_107_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_107_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_107_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_107_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_107_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_107_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_107_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__1__109_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_119_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_119_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_119_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_119_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_119_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_119_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_119_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_119_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_1__1__106_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_106_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_106_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_106_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_106_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_106_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_106_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_106_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_106_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__98_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_107_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_107_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_107_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_107_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_107_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_107_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_107_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_107_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( cbx_1__1__109_ccff_tail ) , 
    .chany_top_out ( sb_1__1__98_chany_top_out ) , 
    .chanx_right_out ( sb_1__1__98_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__1__98_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__1__98_chanx_left_out ) , 
    .ccff_tail ( sb_1__1__98_ccff_tail ) ) ;
sb_1__1_ sb_10__1_ (
    .prog_clk ( { ctsbuf_net_842066 } ) ,
    .chany_top_in ( cby_1__1__109_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_109_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_109_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_109_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_109_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_109_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_109_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_109_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_109_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__1__110_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_121_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_121_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_121_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_121_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_121_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_121_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_121_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_121_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_1__1__108_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_108_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_108_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_108_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_108_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_108_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_108_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_108_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_108_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__99_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_109_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_109_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_109_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_109_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_109_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_109_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_109_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_109_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( cbx_1__1__110_ccff_tail ) , 
    .chany_top_out ( sb_1__1__99_chany_top_out ) , 
    .chanx_right_out ( sb_1__1__99_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__1__99_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__1__99_chanx_left_out ) , 
    .ccff_tail ( sb_1__1__99_ccff_tail ) ) ;
sb_1__1_ sb_10__2_ (
    .prog_clk ( { ctsbuf_net_1132095 } ) ,
    .chany_top_in ( cby_1__1__110_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_110_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_110_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_110_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_110_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_110_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_110_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_110_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_110_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__1__111_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_122_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_122_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_122_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_122_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_122_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_122_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_122_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_122_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_1__1__109_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_109_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_109_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_109_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_109_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_109_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_109_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_109_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_109_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__100_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_110_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_110_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_110_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_110_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_110_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_110_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_110_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_110_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( cbx_1__1__111_ccff_tail ) , 
    .chany_top_out ( sb_1__1__100_chany_top_out ) , 
    .chanx_right_out ( sb_1__1__100_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__1__100_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__1__100_chanx_left_out ) , 
    .ccff_tail ( sb_1__1__100_ccff_tail ) ) ;
sb_1__1_ sb_10__3_ (
    .prog_clk ( { ctsbuf_net_1462128 } ) ,
    .chany_top_in ( cby_1__1__111_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_111_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_111_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_111_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_111_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_111_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_111_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_111_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_111_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__1__112_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_123_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_123_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_123_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_123_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_123_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_123_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_123_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_123_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_1__1__110_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_110_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_110_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_110_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_110_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_110_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_110_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_110_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_110_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__101_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_111_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_111_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_111_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_111_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_111_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_111_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_111_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_111_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( cbx_1__1__112_ccff_tail ) , 
    .chany_top_out ( sb_1__1__101_chany_top_out ) , 
    .chanx_right_out ( sb_1__1__101_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__1__101_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__1__101_chanx_left_out ) , 
    .ccff_tail ( sb_1__1__101_ccff_tail ) ) ;
sb_1__1_ sb_10__4_ (
    .prog_clk ( { ctsbuf_net_1862168 } ) ,
    .chany_top_in ( cby_1__1__112_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_112_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_112_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_112_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_112_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_112_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_112_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_112_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_112_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__1__113_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_124_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_124_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_124_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_124_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_124_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_124_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_124_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_124_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_1__1__111_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_111_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_111_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_111_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_111_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_111_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_111_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_111_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_111_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__102_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_112_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_112_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_112_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_112_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_112_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_112_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_112_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_112_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( cbx_1__1__113_ccff_tail ) , 
    .chany_top_out ( sb_1__1__102_chany_top_out ) , 
    .chanx_right_out ( sb_1__1__102_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__1__102_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__1__102_chanx_left_out ) , 
    .ccff_tail ( sb_1__1__102_ccff_tail ) ) ;
sb_1__1_ sb_10__5_ (
    .prog_clk ( { ctsbuf_net_2312213 } ) ,
    .chany_top_in ( cby_1__1__113_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_113_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_113_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_113_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_113_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_113_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_113_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_113_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_113_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__1__114_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_125_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_125_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_125_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_125_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_125_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_125_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_125_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_125_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_1__1__112_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_112_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_112_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_112_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_112_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_112_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_112_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_112_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_112_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__103_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_113_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_113_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_113_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_113_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_113_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_113_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_113_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_113_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( cbx_1__1__114_ccff_tail ) , 
    .chany_top_out ( sb_1__1__103_chany_top_out ) , 
    .chanx_right_out ( sb_1__1__103_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__1__103_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__1__103_chanx_left_out ) , 
    .ccff_tail ( sb_1__1__103_ccff_tail ) ) ;
sb_1__1_ sb_10__6_ (
    .prog_clk ( { ctsbuf_net_2772259 } ) ,
    .chany_top_in ( cby_1__1__114_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_114_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_114_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_114_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_114_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_114_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_114_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_114_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_114_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__1__115_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_126_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_126_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_126_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_126_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_126_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_126_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_126_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_126_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_1__1__113_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_113_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_113_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_113_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_113_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_113_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_113_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_113_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_113_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__104_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_114_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_114_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_114_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_114_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_114_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_114_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_114_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_114_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( cbx_1__1__115_ccff_tail ) , 
    .chany_top_out ( sb_1__1__104_chany_top_out ) , 
    .chanx_right_out ( sb_1__1__104_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__1__104_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__1__104_chanx_left_out ) , 
    .ccff_tail ( sb_1__1__104_ccff_tail ) ) ;
sb_1__1_ sb_10__7_ (
    .prog_clk ( { ctsbuf_net_2382220 } ) ,
    .chany_top_in ( cby_1__1__115_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_115_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_115_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_115_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_115_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_115_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_115_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_115_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_115_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__1__116_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_127_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_127_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_127_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_127_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_127_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_127_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_127_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_127_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_1__1__114_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_114_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_114_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_114_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_114_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_114_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_114_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_114_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_114_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__105_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_115_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_115_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_115_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_115_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_115_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_115_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_115_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_115_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( cbx_1__1__116_ccff_tail ) , 
    .chany_top_out ( sb_1__1__105_chany_top_out ) , 
    .chanx_right_out ( sb_1__1__105_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__1__105_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__1__105_chanx_left_out ) , 
    .ccff_tail ( sb_1__1__105_ccff_tail ) ) ;
sb_1__1_ sb_10__8_ (
    .prog_clk ( { ctsbuf_net_1922174 } ) ,
    .chany_top_in ( cby_1__1__116_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_116_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_116_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_116_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_116_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_116_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_116_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_116_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_116_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__1__117_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_128_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_128_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_128_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_128_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_128_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_128_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_128_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_128_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_1__1__115_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_115_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_115_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_115_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_115_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_115_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_115_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_115_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_115_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__106_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_116_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_116_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_116_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_116_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_116_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_116_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_116_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_116_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( cbx_1__1__117_ccff_tail ) , 
    .chany_top_out ( sb_1__1__106_chany_top_out ) , 
    .chanx_right_out ( sb_1__1__106_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__1__106_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__1__106_chanx_left_out ) , 
    .ccff_tail ( sb_1__1__106_ccff_tail ) ) ;
sb_1__1_ sb_10__9_ (
    .prog_clk ( { ctsbuf_net_1512133 } ) ,
    .chany_top_in ( cby_1__1__117_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_117_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_117_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_117_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_117_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_117_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_117_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_117_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_117_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__1__118_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_129_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_129_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_129_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_129_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_129_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_129_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_129_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_129_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_1__1__116_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_116_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_116_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_116_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_116_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_116_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_116_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_116_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_116_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__107_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_117_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_117_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_117_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_117_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_117_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_117_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_117_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_117_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( cbx_1__1__118_ccff_tail ) , 
    .chany_top_out ( sb_1__1__107_chany_top_out ) , 
    .chanx_right_out ( sb_1__1__107_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__1__107_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__1__107_chanx_left_out ) , 
    .ccff_tail ( sb_1__1__107_ccff_tail ) ) ;
sb_1__1_ sb_10__10_ (
    .prog_clk ( { ctsbuf_net_1172099 } ) ,
    .chany_top_in ( cby_1__1__118_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_118_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_118_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_118_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_118_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_118_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_118_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_118_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_118_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__1__119_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_130_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_130_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_130_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_130_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_130_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_130_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_130_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_130_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_1__1__117_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_117_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_117_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_117_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_117_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_117_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_117_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_117_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_117_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__108_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_118_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_118_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_118_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_118_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_118_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_118_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_118_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_118_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( cbx_1__1__119_ccff_tail ) , 
    .chany_top_out ( sb_1__1__108_chany_top_out ) , 
    .chanx_right_out ( sb_1__1__108_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__1__108_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__1__108_chanx_left_out ) , 
    .ccff_tail ( sb_1__1__108_ccff_tail ) ) ;
sb_1__1_ sb_10__11_ (
    .prog_clk ( { ctsbuf_net_872069 } ) ,
    .chany_top_in ( cby_1__1__119_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_119_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_119_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_119_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_119_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_119_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_119_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_119_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_119_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__1__120_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_131_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_131_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_131_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_131_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_131_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_131_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_131_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_131_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_1__1__118_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_118_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_118_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_118_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_118_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_118_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_118_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_118_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_118_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__109_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_119_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_119_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_119_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_119_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_119_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_119_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_119_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_119_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( cbx_1__1__120_ccff_tail ) , 
    .chany_top_out ( sb_1__1__109_chany_top_out ) , 
    .chanx_right_out ( sb_1__1__109_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__1__109_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__1__109_chanx_left_out ) , 
    .ccff_tail ( sb_1__1__109_ccff_tail ) ) ;
sb_1__1_ sb_11__1_ (
    .prog_clk ( { p_abuf1 } ) ,
    .chany_top_in ( cby_1__1__121_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_121_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_121_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_121_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_121_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_121_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_121_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_121_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_121_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__1__121_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_133_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_133_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_133_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_133_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_133_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_133_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_133_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_133_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_1__1__120_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_120_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_120_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_120_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_120_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_120_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_120_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_120_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_120_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__110_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_121_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_121_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_121_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_121_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_121_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_121_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_121_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_121_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( cbx_1__1__121_ccff_tail ) , 
    .chany_top_out ( sb_1__1__110_chany_top_out ) , 
    .chanx_right_out ( sb_1__1__110_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__1__110_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__1__110_chanx_left_out ) , 
    .ccff_tail ( sb_1__1__110_ccff_tail ) ) ;
sb_1__1_ sb_11__2_ (
    .prog_clk ( { ctsbuf_net_852067 } ) ,
    .chany_top_in ( cby_1__1__122_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_122_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_122_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_122_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_122_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_122_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_122_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_122_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_122_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__1__122_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_134_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_134_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_134_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_134_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_134_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_134_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_134_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_134_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_1__1__121_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_121_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_121_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_121_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_121_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_121_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_121_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_121_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_121_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__111_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_122_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_122_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_122_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_122_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_122_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_122_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_122_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_122_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( cbx_1__1__122_ccff_tail ) , 
    .chany_top_out ( sb_1__1__111_chany_top_out ) , 
    .chanx_right_out ( sb_1__1__111_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__1__111_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__1__111_chanx_left_out ) , 
    .ccff_tail ( sb_1__1__111_ccff_tail ) ) ;
sb_1__1_ sb_11__3_ (
    .prog_clk ( { ctsbuf_net_1142096 } ) ,
    .chany_top_in ( cby_1__1__123_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_123_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_123_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_123_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_123_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_123_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_123_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_123_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_123_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__1__123_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_135_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_135_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_135_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_135_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_135_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_135_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_135_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_135_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_1__1__122_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_122_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_122_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_122_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_122_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_122_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_122_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_122_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_122_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__112_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_123_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_123_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_123_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_123_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_123_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_123_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_123_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_123_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( cbx_1__1__123_ccff_tail ) , 
    .chany_top_out ( sb_1__1__112_chany_top_out ) , 
    .chanx_right_out ( sb_1__1__112_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__1__112_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__1__112_chanx_left_out ) , 
    .ccff_tail ( sb_1__1__112_ccff_tail ) ) ;
sb_1__1_ sb_11__4_ (
    .prog_clk ( { ctsbuf_net_1472129 } ) ,
    .chany_top_in ( cby_1__1__124_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_124_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_124_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_124_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_124_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_124_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_124_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_124_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_124_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__1__124_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_136_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_136_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_136_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_136_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_136_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_136_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_136_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_136_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_1__1__123_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_123_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_123_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_123_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_123_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_123_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_123_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_123_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_123_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__113_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_124_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_124_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_124_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_124_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_124_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_124_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_124_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_124_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( cbx_1__1__124_ccff_tail ) , 
    .chany_top_out ( sb_1__1__113_chany_top_out ) , 
    .chanx_right_out ( sb_1__1__113_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__1__113_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__1__113_chanx_left_out ) , 
    .ccff_tail ( sb_1__1__113_ccff_tail ) ) ;
sb_1__1_ sb_11__5_ (
    .prog_clk ( { ctsbuf_net_1872169 } ) ,
    .chany_top_in ( cby_1__1__125_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_125_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_125_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_125_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_125_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_125_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_125_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_125_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_125_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__1__125_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_137_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_137_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_137_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_137_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_137_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_137_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_137_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_137_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_1__1__124_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_124_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_124_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_124_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_124_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_124_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_124_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_124_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_124_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__114_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_125_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_125_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_125_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_125_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_125_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_125_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_125_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_125_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( cbx_1__1__125_ccff_tail ) , 
    .chany_top_out ( sb_1__1__114_chany_top_out ) , 
    .chanx_right_out ( sb_1__1__114_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__1__114_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__1__114_chanx_left_out ) , 
    .ccff_tail ( sb_1__1__114_ccff_tail ) ) ;
sb_1__1_ sb_11__6_ (
    .prog_clk ( { ctsbuf_net_2322214 } ) ,
    .chany_top_in ( cby_1__1__126_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_126_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_126_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_126_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_126_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_126_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_126_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_126_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_126_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__1__126_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_138_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_138_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_138_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_138_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_138_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_138_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_138_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_138_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_1__1__125_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_125_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_125_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_125_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_125_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_125_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_125_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_125_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_125_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__115_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_126_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_126_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_126_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_126_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_126_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_126_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_126_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_126_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( cbx_1__1__126_ccff_tail ) , 
    .chany_top_out ( sb_1__1__115_chany_top_out ) , 
    .chanx_right_out ( sb_1__1__115_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__1__115_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__1__115_chanx_left_out ) , 
    .ccff_tail ( sb_1__1__115_ccff_tail ) ) ;
sb_1__1_ sb_11__7_ (
    .prog_clk ( { ctsbuf_net_1932175 } ) ,
    .chany_top_in ( cby_1__1__127_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_127_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_127_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_127_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_127_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_127_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_127_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_127_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_127_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__1__127_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_139_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_139_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_139_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_139_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_139_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_139_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_139_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_139_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_1__1__126_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_126_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_126_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_126_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_126_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_126_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_126_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_126_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_126_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__116_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_127_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_127_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_127_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_127_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_127_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_127_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_127_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_127_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( cbx_1__1__127_ccff_tail ) , 
    .chany_top_out ( sb_1__1__116_chany_top_out ) , 
    .chanx_right_out ( sb_1__1__116_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__1__116_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__1__116_chanx_left_out ) , 
    .ccff_tail ( sb_1__1__116_ccff_tail ) ) ;
sb_1__1_ sb_11__8_ (
    .prog_clk ( { ctsbuf_net_1522134 } ) ,
    .chany_top_in ( cby_1__1__128_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_128_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_128_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_128_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_128_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_128_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_128_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_128_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_128_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__1__128_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_140_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_140_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_140_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_140_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_140_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_140_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_140_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_140_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_1__1__127_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_127_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_127_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_127_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_127_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_127_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_127_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_127_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_127_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__117_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_128_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_128_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_128_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_128_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_128_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_128_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_128_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_128_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( cbx_1__1__128_ccff_tail ) , 
    .chany_top_out ( sb_1__1__117_chany_top_out ) , 
    .chanx_right_out ( sb_1__1__117_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__1__117_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__1__117_chanx_left_out ) , 
    .ccff_tail ( sb_1__1__117_ccff_tail ) ) ;
sb_1__1_ sb_11__9_ (
    .prog_clk ( { ctsbuf_net_1182100 } ) ,
    .chany_top_in ( cby_1__1__129_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_129_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_129_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_129_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_129_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_129_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_129_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_129_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_129_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__1__129_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_141_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_141_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_141_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_141_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_141_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_141_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_141_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_141_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_1__1__128_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_128_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_128_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_128_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_128_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_128_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_128_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_128_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_128_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__118_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_129_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_129_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_129_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_129_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_129_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_129_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_129_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_129_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( cbx_1__1__129_ccff_tail ) , 
    .chany_top_out ( sb_1__1__118_chany_top_out ) , 
    .chanx_right_out ( sb_1__1__118_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__1__118_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__1__118_chanx_left_out ) , 
    .ccff_tail ( sb_1__1__118_ccff_tail ) ) ;
sb_1__1_ sb_11__10_ (
    .prog_clk ( { ctsbuf_net_892071 } ) ,
    .chany_top_in ( cby_1__1__130_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_130_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_130_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_130_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_130_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_130_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_130_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_130_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_130_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__1__130_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_142_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_142_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_142_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_142_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_142_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_142_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_142_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_142_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_1__1__129_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_129_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_129_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_129_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_129_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_129_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_129_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_129_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_129_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__119_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_130_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_130_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_130_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_130_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_130_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_130_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_130_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_130_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( cbx_1__1__130_ccff_tail ) , 
    .chany_top_out ( sb_1__1__119_chany_top_out ) , 
    .chanx_right_out ( sb_1__1__119_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__1__119_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__1__119_chanx_left_out ) , 
    .ccff_tail ( sb_1__1__119_ccff_tail ) ) ;
sb_1__1_ sb_11__11_ (
    .prog_clk ( { ctsbuf_net_722054 } ) ,
    .chany_top_in ( cby_1__1__131_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_131_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_131_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_131_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_131_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_131_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_131_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_131_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_131_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__1__131_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_143_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_143_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_143_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_143_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_143_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_143_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_143_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_143_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_1__1__130_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_130_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_130_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_130_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_130_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_130_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_130_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_130_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_130_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__120_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_131_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_131_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_131_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_131_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_131_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_131_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_131_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_131_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( cbx_1__1__131_ccff_tail ) , 
    .chany_top_out ( sb_1__1__120_chany_top_out ) , 
    .chanx_right_out ( sb_1__1__120_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__1__120_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__1__120_chanx_left_out ) , 
    .ccff_tail ( sb_1__1__120_ccff_tail ) ) ;
sb_1__2_ sb_1__12_ (
    .prog_clk ( { ctsbuf_net_3882370 } ) ,
    .chanx_right_in ( cbx_1__12__1_chanx_left_out ) , 
    .right_top_grid_pin_1_ ( grid_io_top_1_bottom_width_0_height_0__pin_1_upper ) , 
    .chany_bottom_in ( cby_1__1__11_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_11_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_11_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_11_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_11_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_11_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_11_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_11_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_11_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__12__0_chanx_right_out ) , 
    .left_top_grid_pin_1_ ( grid_io_top_0_bottom_width_0_height_0__pin_1_lower ) , 
    .ccff_head ( grid_io_top_1_ccff_tail ) , 
    .chanx_right_out ( sb_1__12__0_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__12__0_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__12__0_chanx_left_out ) , 
    .ccff_tail ( sb_1__12__0_ccff_tail ) ) ;
sb_1__2_ sb_2__12_ (
    .prog_clk ( { ctsbuf_net_3292311 } ) ,
    .chanx_right_in ( cbx_1__12__2_chanx_left_out ) , 
    .right_top_grid_pin_1_ ( grid_io_top_2_bottom_width_0_height_0__pin_1_upper ) , 
    .chany_bottom_in ( cby_1__1__23_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_23_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_23_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_23_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_23_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_23_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_23_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_23_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_23_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__12__1_chanx_right_out ) , 
    .left_top_grid_pin_1_ ( grid_io_top_1_bottom_width_0_height_0__pin_1_lower ) , 
    .ccff_head ( grid_io_top_2_ccff_tail ) , 
    .chanx_right_out ( sb_1__12__1_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__12__1_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__12__1_chanx_left_out ) , 
    .ccff_tail ( sb_1__12__1_ccff_tail ) ) ;
sb_1__2_ sb_3__12_ (
    .prog_clk ( { ctsbuf_net_3002282 } ) ,
    .chanx_right_in ( cbx_1__12__3_chanx_left_out ) , 
    .right_top_grid_pin_1_ ( grid_io_top_3_bottom_width_0_height_0__pin_1_upper ) , 
    .chany_bottom_in ( cby_1__1__35_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_35_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_35_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_35_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_35_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_35_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_35_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_35_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_35_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__12__2_chanx_right_out ) , 
    .left_top_grid_pin_1_ ( grid_io_top_2_bottom_width_0_height_0__pin_1_lower ) , 
    .ccff_head ( grid_io_top_3_ccff_tail ) , 
    .chanx_right_out ( sb_1__12__2_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__12__2_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__12__2_chanx_left_out ) , 
    .ccff_tail ( sb_1__12__2_ccff_tail ) ) ;
sb_1__2_ sb_4__12_ (
    .prog_clk ( { p_abuf13 } ) ,
    .chanx_right_in ( cbx_1__12__4_chanx_left_out ) , 
    .right_top_grid_pin_1_ ( grid_io_top_4_bottom_width_0_height_0__pin_1_upper ) , 
    .chany_bottom_in ( cby_1__1__47_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_47_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_47_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_47_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_47_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_47_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_47_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_47_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_47_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__12__3_chanx_right_out ) , 
    .left_top_grid_pin_1_ ( grid_io_top_3_bottom_width_0_height_0__pin_1_lower ) , 
    .ccff_head ( grid_io_top_4_ccff_tail ) , 
    .chanx_right_out ( sb_1__12__3_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__12__3_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__12__3_chanx_left_out ) , 
    .ccff_tail ( sb_1__12__3_ccff_tail ) ) ;
sb_1__2_ sb_5__12_ (
    .prog_clk ( { ctsbuf_net_2102192 } ) ,
    .chanx_right_in ( cbx_1__12__5_chanx_left_out ) , 
    .right_top_grid_pin_1_ ( grid_io_top_5_bottom_width_0_height_0__pin_1_upper ) , 
    .chany_bottom_in ( cby_1__1__59_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_59_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_59_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_59_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_59_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_59_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_59_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_59_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_59_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__12__4_chanx_right_out ) , 
    .left_top_grid_pin_1_ ( grid_io_top_4_bottom_width_0_height_0__pin_1_lower ) , 
    .ccff_head ( grid_io_top_5_ccff_tail ) , 
    .chanx_right_out ( sb_1__12__4_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__12__4_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__12__4_chanx_left_out ) , 
    .ccff_tail ( sb_1__12__4_ccff_tail ) ) ;
sb_1__2_ sb_6__12_ (
    .prog_clk ( { ctsbuf_net_1532135 } ) ,
    .chanx_right_in ( cbx_1__12__6_chanx_left_out ) , 
    .right_top_grid_pin_1_ ( grid_io_top_6_bottom_width_0_height_0__pin_1_upper ) , 
    .chany_bottom_in ( cby_1__1__71_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_71_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_71_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_71_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_71_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_71_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_71_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_71_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_71_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__12__5_chanx_right_out ) , 
    .left_top_grid_pin_1_ ( grid_io_top_5_bottom_width_0_height_0__pin_1_lower ) , 
    .ccff_head ( grid_io_top_6_ccff_tail ) , 
    .chanx_right_out ( sb_1__12__5_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__12__5_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__12__5_chanx_left_out ) , 
    .ccff_tail ( sb_1__12__5_ccff_tail ) ) ;
sb_1__2_ sb_7__12_ (
    .prog_clk ( { ctsbuf_net_1312113 } ) ,
    .chanx_right_in ( cbx_1__12__7_chanx_left_out ) , 
    .right_top_grid_pin_1_ ( grid_io_top_7_bottom_width_0_height_0__pin_1_upper ) , 
    .chany_bottom_in ( cby_1__1__83_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_83_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_83_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_83_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_83_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_83_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_83_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_83_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_83_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__12__6_chanx_right_out ) , 
    .left_top_grid_pin_1_ ( grid_io_top_6_bottom_width_0_height_0__pin_1_lower ) , 
    .ccff_head ( grid_io_top_7_ccff_tail ) , 
    .chanx_right_out ( sb_1__12__6_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__12__6_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__12__6_chanx_left_out ) , 
    .ccff_tail ( sb_1__12__6_ccff_tail ) ) ;
sb_1__2_ sb_8__12_ (
    .prog_clk ( { p_abuf4 } ) ,
    .chanx_right_in ( cbx_1__12__8_chanx_left_out ) , 
    .right_top_grid_pin_1_ ( grid_io_top_8_bottom_width_0_height_0__pin_1_upper ) , 
    .chany_bottom_in ( cby_1__1__95_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_95_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_95_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_95_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_95_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_95_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_95_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_95_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_95_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__12__7_chanx_right_out ) , 
    .left_top_grid_pin_1_ ( grid_io_top_7_bottom_width_0_height_0__pin_1_lower ) , 
    .ccff_head ( grid_io_top_8_ccff_tail ) , 
    .chanx_right_out ( sb_1__12__7_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__12__7_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__12__7_chanx_left_out ) , 
    .ccff_tail ( sb_1__12__7_ccff_tail ) ) ;
sb_1__2_ sb_9__12_ (
    .prog_clk ( { ctsbuf_net_752057 } ) ,
    .chanx_right_in ( cbx_1__12__9_chanx_left_out ) , 
    .right_top_grid_pin_1_ ( grid_io_top_9_bottom_width_0_height_0__pin_1_upper ) , 
    .chany_bottom_in ( cby_1__1__107_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_107_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_107_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_107_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_107_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_107_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_107_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_107_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_107_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__12__8_chanx_right_out ) , 
    .left_top_grid_pin_1_ ( grid_io_top_8_bottom_width_0_height_0__pin_1_lower ) , 
    .ccff_head ( grid_io_top_9_ccff_tail ) , 
    .chanx_right_out ( sb_1__12__8_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__12__8_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__12__8_chanx_left_out ) , 
    .ccff_tail ( sb_1__12__8_ccff_tail ) ) ;
sb_1__2_ sb_10__12_ (
    .prog_clk ( { ctsbuf_net_532035 } ) ,
    .chanx_right_in ( cbx_1__12__10_chanx_left_out ) , 
    .right_top_grid_pin_1_ ( grid_io_top_10_bottom_width_0_height_0__pin_1_upper ) , 
    .chany_bottom_in ( cby_1__1__119_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_119_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_119_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_119_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_119_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_119_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_119_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_119_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_119_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__12__9_chanx_right_out ) , 
    .left_top_grid_pin_1_ ( grid_io_top_9_bottom_width_0_height_0__pin_1_lower ) , 
    .ccff_head ( grid_io_top_10_ccff_tail ) , 
    .chanx_right_out ( sb_1__12__9_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__12__9_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__12__9_chanx_left_out ) , 
    .ccff_tail ( sb_1__12__9_ccff_tail ) ) ;
sb_1__2_ sb_11__12_ (
    .prog_clk ( { ctsbuf_net_512033 } ) ,
    .chanx_right_in ( cbx_1__12__11_chanx_left_out ) , 
    .right_top_grid_pin_1_ ( grid_io_top_11_bottom_width_0_height_0__pin_1_upper ) , 
    .chany_bottom_in ( cby_1__1__131_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_131_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_131_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_131_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_131_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_131_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_131_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_131_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_131_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__12__10_chanx_right_out ) , 
    .left_top_grid_pin_1_ ( grid_io_top_10_bottom_width_0_height_0__pin_1_lower ) , 
    .ccff_head ( grid_io_top_11_ccff_tail ) , 
    .chanx_right_out ( sb_1__12__10_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__12__10_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__12__10_chanx_left_out ) , 
    .ccff_tail ( sb_1__12__10_ccff_tail ) ) ;
sb_2__0_ sb_12__0_ (
    .prog_clk ( { ctsbuf_net_452027 } ) ,
    .chany_top_in ( cby_1__1__132_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_132_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_132_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_132_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_132_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_132_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_132_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_132_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_132_right_width_0_height_0__pin_41_lower ) , 
    .top_right_grid_pin_1_ ( grid_io_right_0_left_width_0_height_0__pin_1_lower ) , 
    .chanx_left_in ( cbx_1__0__11_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_132_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_132_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_132_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_132_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_132_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_132_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_132_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_132_bottom_width_0_height_0__pin_49_lower ) , 
    .left_bottom_grid_pin_1_ ( grid_io_bottom_11_top_width_0_height_0__pin_1_lower ) , 
    .ccff_head ( grid_io_right_0_ccff_tail ) , 
    .chany_top_out ( sb_12__0__0_chany_top_out ) , 
    .chanx_left_out ( sb_12__0__0_chanx_left_out ) , 
    .ccff_tail ( sb_12__0__0_ccff_tail ) ) ;
sb_2__1_ sb_12__1_ (
    .prog_clk ( { ctsbuf_net_502032 } ) ,
    .chany_top_in ( cby_1__1__133_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_133_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_133_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_133_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_133_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_133_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_133_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_133_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_133_right_width_0_height_0__pin_41_lower ) , 
    .top_right_grid_pin_1_ ( grid_io_right_1_left_width_0_height_0__pin_1_lower ) , 
    .chany_bottom_in ( cby_1__1__132_chany_top_out ) , 
    .bottom_right_grid_pin_1_ ( grid_io_right_0_left_width_0_height_0__pin_1_upper ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_132_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_132_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_132_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_132_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_132_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_132_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_132_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_132_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__121_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_133_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_133_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_133_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_133_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_133_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_133_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_133_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_133_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( grid_io_right_1_ccff_tail ) , 
    .chany_top_out ( sb_12__1__0_chany_top_out ) , 
    .chany_bottom_out ( sb_12__1__0_chany_bottom_out ) , 
    .chanx_left_out ( sb_12__1__0_chanx_left_out ) , 
    .ccff_tail ( sb_12__1__0_ccff_tail ) ) ;
sb_2__1_ sb_12__2_ (
    .prog_clk ( { ctsbuf_net_652047 } ) ,
    .chany_top_in ( cby_1__1__134_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_134_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_134_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_134_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_134_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_134_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_134_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_134_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_134_right_width_0_height_0__pin_41_lower ) , 
    .top_right_grid_pin_1_ ( grid_io_right_2_left_width_0_height_0__pin_1_lower ) , 
    .chany_bottom_in ( cby_1__1__133_chany_top_out ) , 
    .bottom_right_grid_pin_1_ ( grid_io_right_1_left_width_0_height_0__pin_1_upper ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_133_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_133_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_133_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_133_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_133_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_133_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_133_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_133_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__122_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_134_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_134_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_134_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_134_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_134_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_134_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_134_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_134_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( grid_io_right_2_ccff_tail ) , 
    .chany_top_out ( sb_12__1__1_chany_top_out ) , 
    .chany_bottom_out ( sb_12__1__1_chany_bottom_out ) , 
    .chanx_left_out ( sb_12__1__1_chanx_left_out ) , 
    .ccff_tail ( sb_12__1__1_ccff_tail ) ) ;
sb_2__1_ sb_12__3_ (
    .prog_clk ( { ctsbuf_net_862068 } ) ,
    .chany_top_in ( cby_1__1__135_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_135_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_135_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_135_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_135_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_135_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_135_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_135_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_135_right_width_0_height_0__pin_41_lower ) , 
    .top_right_grid_pin_1_ ( grid_io_right_3_left_width_0_height_0__pin_1_lower ) , 
    .chany_bottom_in ( cby_1__1__134_chany_top_out ) , 
    .bottom_right_grid_pin_1_ ( grid_io_right_2_left_width_0_height_0__pin_1_upper ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_134_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_134_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_134_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_134_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_134_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_134_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_134_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_134_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__123_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_135_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_135_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_135_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_135_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_135_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_135_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_135_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_135_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( grid_io_right_3_ccff_tail ) , 
    .chany_top_out ( sb_12__1__2_chany_top_out ) , 
    .chany_bottom_out ( sb_12__1__2_chany_bottom_out ) , 
    .chanx_left_out ( sb_12__1__2_chanx_left_out ) , 
    .ccff_tail ( sb_12__1__2_ccff_tail ) ) ;
sb_2__1_ sb_12__4_ (
    .prog_clk ( { ctsbuf_net_1112093 } ) ,
    .chany_top_in ( cby_1__1__136_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_136_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_136_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_136_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_136_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_136_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_136_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_136_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_136_right_width_0_height_0__pin_41_lower ) , 
    .top_right_grid_pin_1_ ( grid_io_right_4_left_width_0_height_0__pin_1_lower ) , 
    .chany_bottom_in ( cby_1__1__135_chany_top_out ) , 
    .bottom_right_grid_pin_1_ ( grid_io_right_3_left_width_0_height_0__pin_1_upper ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_135_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_135_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_135_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_135_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_135_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_135_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_135_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_135_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__124_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_136_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_136_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_136_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_136_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_136_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_136_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_136_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_136_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( grid_io_right_4_ccff_tail ) , 
    .chany_top_out ( sb_12__1__3_chany_top_out ) , 
    .chany_bottom_out ( sb_12__1__3_chany_bottom_out ) , 
    .chanx_left_out ( sb_12__1__3_chanx_left_out ) , 
    .ccff_tail ( sb_12__1__3_ccff_tail ) ) ;
sb_2__1_ sb_12__5_ (
    .prog_clk ( { ctsbuf_net_1432125 } ) ,
    .chany_top_in ( cby_1__1__137_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_137_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_137_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_137_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_137_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_137_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_137_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_137_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_137_right_width_0_height_0__pin_41_lower ) , 
    .top_right_grid_pin_1_ ( grid_io_right_5_left_width_0_height_0__pin_1_lower ) , 
    .chany_bottom_in ( cby_1__1__136_chany_top_out ) , 
    .bottom_right_grid_pin_1_ ( grid_io_right_4_left_width_0_height_0__pin_1_upper ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_136_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_136_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_136_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_136_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_136_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_136_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_136_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_136_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__125_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_137_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_137_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_137_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_137_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_137_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_137_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_137_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_137_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( grid_io_right_5_ccff_tail ) , 
    .chany_top_out ( sb_12__1__4_chany_top_out ) , 
    .chany_bottom_out ( sb_12__1__4_chany_bottom_out ) , 
    .chanx_left_out ( sb_12__1__4_chanx_left_out ) , 
    .ccff_tail ( sb_12__1__4_ccff_tail ) ) ;
sb_2__1_ sb_12__6_ (
    .prog_clk ( { ctsbuf_net_1762158 } ) ,
    .chany_top_in ( cby_1__1__138_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_138_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_138_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_138_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_138_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_138_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_138_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_138_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_138_right_width_0_height_0__pin_41_lower ) , 
    .top_right_grid_pin_1_ ( grid_io_right_6_left_width_0_height_0__pin_1_lower ) , 
    .chany_bottom_in ( cby_1__1__137_chany_top_out ) , 
    .bottom_right_grid_pin_1_ ( grid_io_right_5_left_width_0_height_0__pin_1_upper ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_137_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_137_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_137_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_137_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_137_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_137_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_137_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_137_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__126_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_138_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_138_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_138_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_138_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_138_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_138_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_138_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_138_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( grid_io_right_6_ccff_tail ) , 
    .chany_top_out ( sb_12__1__5_chany_top_out ) , 
    .chany_bottom_out ( sb_12__1__5_chany_bottom_out ) , 
    .chanx_left_out ( sb_12__1__5_chanx_left_out ) , 
    .ccff_tail ( sb_12__1__5_ccff_tail ) ) ;
sb_2__1_ sb_12__7_ (
    .prog_clk ( { ctsbuf_net_1202102 } ) ,
    .chany_top_in ( cby_1__1__139_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_139_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_139_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_139_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_139_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_139_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_139_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_139_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_139_right_width_0_height_0__pin_41_lower ) , 
    .top_right_grid_pin_1_ ( grid_io_right_7_left_width_0_height_0__pin_1_lower ) , 
    .chany_bottom_in ( cby_1__1__138_chany_top_out ) , 
    .bottom_right_grid_pin_1_ ( grid_io_right_6_left_width_0_height_0__pin_1_upper ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_138_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_138_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_138_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_138_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_138_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_138_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_138_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_138_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__127_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_139_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_139_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_139_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_139_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_139_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_139_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_139_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_139_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( grid_io_right_7_ccff_tail ) , 
    .chany_top_out ( sb_12__1__6_chany_top_out ) , 
    .chany_bottom_out ( sb_12__1__6_chany_bottom_out ) , 
    .chanx_left_out ( sb_12__1__6_chanx_left_out ) , 
    .ccff_tail ( sb_12__1__6_ccff_tail ) ) ;
sb_2__1_ sb_12__8_ (
    .prog_clk ( { ctsbuf_net_1192101 } ) ,
    .chany_top_in ( cby_1__1__140_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_140_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_140_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_140_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_140_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_140_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_140_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_140_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_140_right_width_0_height_0__pin_41_lower ) , 
    .top_right_grid_pin_1_ ( grid_io_right_8_left_width_0_height_0__pin_1_lower ) , 
    .chany_bottom_in ( cby_1__1__139_chany_top_out ) , 
    .bottom_right_grid_pin_1_ ( grid_io_right_7_left_width_0_height_0__pin_1_upper ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_139_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_139_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_139_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_139_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_139_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_139_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_139_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_139_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__128_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_140_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_140_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_140_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_140_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_140_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_140_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_140_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_140_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( grid_io_right_8_ccff_tail ) , 
    .chany_top_out ( sb_12__1__7_chany_top_out ) , 
    .chany_bottom_out ( sb_12__1__7_chany_bottom_out ) , 
    .chanx_left_out ( sb_12__1__7_chanx_left_out ) , 
    .ccff_tail ( sb_12__1__7_ccff_tail ) ) ;
sb_2__1_ sb_12__9_ (
    .prog_clk ( { ctsbuf_net_902072 } ) ,
    .chany_top_in ( cby_1__1__141_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_141_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_141_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_141_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_141_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_141_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_141_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_141_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_141_right_width_0_height_0__pin_41_lower ) , 
    .top_right_grid_pin_1_ ( grid_io_right_9_left_width_0_height_0__pin_1_lower ) , 
    .chany_bottom_in ( cby_1__1__140_chany_top_out ) , 
    .bottom_right_grid_pin_1_ ( grid_io_right_8_left_width_0_height_0__pin_1_upper ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_140_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_140_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_140_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_140_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_140_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_140_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_140_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_140_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__129_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_141_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_141_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_141_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_141_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_141_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_141_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_141_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_141_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( grid_io_right_9_ccff_tail ) , 
    .chany_top_out ( sb_12__1__8_chany_top_out ) , 
    .chany_bottom_out ( sb_12__1__8_chany_bottom_out ) , 
    .chanx_left_out ( sb_12__1__8_chanx_left_out ) , 
    .ccff_tail ( sb_12__1__8_ccff_tail ) ) ;
sb_2__1_ sb_12__10_ (
    .prog_clk ( { ctsbuf_net_602042 } ) ,
    .chany_top_in ( cby_1__1__142_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_142_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_142_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_142_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_142_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_142_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_142_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_142_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_142_right_width_0_height_0__pin_41_lower ) , 
    .top_right_grid_pin_1_ ( grid_io_right_10_left_width_0_height_0__pin_1_lower ) , 
    .chany_bottom_in ( cby_1__1__141_chany_top_out ) , 
    .bottom_right_grid_pin_1_ ( grid_io_right_9_left_width_0_height_0__pin_1_upper ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_141_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_141_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_141_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_141_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_141_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_141_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_141_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_141_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__130_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_142_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_142_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_142_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_142_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_142_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_142_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_142_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_142_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( grid_io_right_10_ccff_tail ) , 
    .chany_top_out ( sb_12__1__9_chany_top_out ) , 
    .chany_bottom_out ( sb_12__1__9_chany_bottom_out ) , 
    .chanx_left_out ( sb_12__1__9_chanx_left_out ) , 
    .ccff_tail ( sb_12__1__9_ccff_tail ) ) ;
sb_2__1_ sb_12__11_ (
    .prog_clk ( { ctsbuf_net_472029 } ) ,
    .chany_top_in ( cby_1__1__143_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_143_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_143_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_143_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_143_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_143_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_143_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_143_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_143_right_width_0_height_0__pin_41_lower ) , 
    .top_right_grid_pin_1_ ( grid_io_right_11_left_width_0_height_0__pin_1_lower ) , 
    .chany_bottom_in ( cby_1__1__142_chany_top_out ) , 
    .bottom_right_grid_pin_1_ ( grid_io_right_10_left_width_0_height_0__pin_1_upper ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_142_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_142_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_142_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_142_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_142_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_142_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_142_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_142_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__131_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_143_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_143_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_143_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_143_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_143_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_143_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_143_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_143_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( grid_io_right_11_ccff_tail ) , 
    .chany_top_out ( sb_12__1__10_chany_top_out ) , 
    .chany_bottom_out ( sb_12__1__10_chany_bottom_out ) , 
    .chanx_left_out ( sb_12__1__10_chanx_left_out ) , 
    .ccff_tail ( sb_12__1__10_ccff_tail ) ) ;
sb_2__2_ sb_12__12_ (
    .prog_clk ( { ctsbuf_net_462028 } ) ,
    .chany_bottom_in ( cby_1__1__143_chany_top_out ) , 
    .bottom_right_grid_pin_1_ ( grid_io_right_11_left_width_0_height_0__pin_1_upper ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_143_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_143_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_143_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_143_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_143_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_143_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_143_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_143_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__12__11_chanx_right_out ) , 
    .left_top_grid_pin_1_ ( grid_io_top_11_bottom_width_0_height_0__pin_1_lower ) , 
    .ccff_head ( ccff_head ) , 
    .chany_bottom_out ( sb_12__12__0_chany_bottom_out ) , 
    .chanx_left_out ( sb_12__12__0_chanx_left_out ) , 
    .ccff_tail ( sb_12__12__0_ccff_tail ) ) ;
cbx_1__0_ cbx_1__0_ (
    .prog_clk ( { ctsbuf_net_4172399 } ) ,
    .chanx_left_in ( sb_0__0__0_chanx_right_out ) , 
    .chanx_right_in ( sb_1__0__0_chanx_left_out ) , 
    .ccff_head ( sb_1__0__0_ccff_tail ) , 
    .chanx_left_out ( cbx_1__0__0_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__0__0_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__0__0_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__0__0_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__0__0_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__0__0_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__0__0_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__0__0_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__0__0_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__0__0_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__0__0_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__0__0_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__0__0_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__0__0_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__0__0_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__0__0_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__0__0_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__0__0_top_grid_pin_31_ ) , 
    .bottom_grid_pin_0_ ( cbx_1__0__0_bottom_grid_pin_0_ ) , 
    .ccff_tail ( cbx_1__0__0_ccff_tail ) ) ;
cbx_1__0_ cbx_2__0_ (
    .prog_clk ( { ctsbuf_net_3732355 } ) ,
    .chanx_left_in ( sb_1__0__0_chanx_right_out ) , 
    .chanx_right_in ( sb_1__0__1_chanx_left_out ) , 
    .ccff_head ( sb_1__0__1_ccff_tail ) , 
    .chanx_left_out ( cbx_1__0__1_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__0__1_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__0__1_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__0__1_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__0__1_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__0__1_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__0__1_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__0__1_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__0__1_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__0__1_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__0__1_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__0__1_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__0__1_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__0__1_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__0__1_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__0__1_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__0__1_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__0__1_top_grid_pin_31_ ) , 
    .bottom_grid_pin_0_ ( cbx_1__0__1_bottom_grid_pin_0_ ) , 
    .ccff_tail ( cbx_1__0__1_ccff_tail ) ) ;
cbx_1__0_ cbx_3__0_ (
    .prog_clk ( { ctsbuf_net_3302312 } ) ,
    .chanx_left_in ( sb_1__0__1_chanx_right_out ) , 
    .chanx_right_in ( sb_1__0__2_chanx_left_out ) , 
    .ccff_head ( sb_1__0__2_ccff_tail ) , 
    .chanx_left_out ( cbx_1__0__2_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__0__2_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__0__2_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__0__2_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__0__2_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__0__2_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__0__2_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__0__2_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__0__2_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__0__2_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__0__2_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__0__2_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__0__2_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__0__2_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__0__2_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__0__2_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__0__2_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__0__2_top_grid_pin_31_ ) , 
    .bottom_grid_pin_0_ ( cbx_1__0__2_bottom_grid_pin_0_ ) , 
    .ccff_tail ( cbx_1__0__2_ccff_tail ) ) ;
cbx_1__0_ cbx_4__0_ (
    .prog_clk ( { ctsbuf_net_2842266 } ) ,
    .chanx_left_in ( sb_1__0__2_chanx_right_out ) , 
    .chanx_right_in ( sb_1__0__3_chanx_left_out ) , 
    .ccff_head ( sb_1__0__3_ccff_tail ) , 
    .chanx_left_out ( cbx_1__0__3_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__0__3_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__0__3_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__0__3_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__0__3_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__0__3_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__0__3_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__0__3_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__0__3_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__0__3_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__0__3_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__0__3_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__0__3_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__0__3_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__0__3_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__0__3_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__0__3_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__0__3_top_grid_pin_31_ ) , 
    .bottom_grid_pin_0_ ( cbx_1__0__3_bottom_grid_pin_0_ ) , 
    .ccff_tail ( cbx_1__0__3_ccff_tail ) ) ;
cbx_1__0_ cbx_5__0_ (
    .prog_clk ( { ctsbuf_net_2402222 } ) ,
    .chanx_left_in ( sb_1__0__3_chanx_right_out ) , 
    .chanx_right_in ( sb_1__0__4_chanx_left_out ) , 
    .ccff_head ( sb_1__0__4_ccff_tail ) , 
    .chanx_left_out ( cbx_1__0__4_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__0__4_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__0__4_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__0__4_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__0__4_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__0__4_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__0__4_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__0__4_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__0__4_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__0__4_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__0__4_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__0__4_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__0__4_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__0__4_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__0__4_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__0__4_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__0__4_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__0__4_top_grid_pin_31_ ) , 
    .bottom_grid_pin_0_ ( cbx_1__0__4_bottom_grid_pin_0_ ) , 
    .ccff_tail ( cbx_1__0__4_ccff_tail ) ) ;
cbx_1__0_ cbx_6__0_ (
    .prog_clk ( { ctsbuf_net_1942176 } ) ,
    .chanx_left_in ( sb_1__0__4_chanx_right_out ) , 
    .chanx_right_in ( sb_1__0__5_chanx_left_out ) , 
    .ccff_head ( sb_1__0__5_ccff_tail ) , 
    .chanx_left_out ( cbx_1__0__5_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__0__5_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__0__5_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__0__5_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__0__5_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__0__5_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__0__5_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__0__5_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__0__5_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__0__5_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__0__5_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__0__5_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__0__5_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__0__5_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__0__5_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__0__5_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__0__5_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__0__5_top_grid_pin_31_ ) , 
    .bottom_grid_pin_0_ ( cbx_1__0__5_bottom_grid_pin_0_ ) , 
    .ccff_tail ( cbx_1__0__5_ccff_tail ) ) ;
cbx_1__0_ cbx_7__0_ (
    .prog_clk ( { ctsbuf_net_1542136 } ) ,
    .chanx_left_in ( sb_1__0__5_chanx_right_out ) , 
    .chanx_right_in ( sb_1__0__6_chanx_left_out ) , 
    .ccff_head ( sb_1__0__6_ccff_tail ) , 
    .chanx_left_out ( cbx_1__0__6_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__0__6_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__0__6_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__0__6_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__0__6_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__0__6_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__0__6_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__0__6_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__0__6_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__0__6_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__0__6_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__0__6_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__0__6_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__0__6_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__0__6_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__0__6_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__0__6_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__0__6_top_grid_pin_31_ ) , 
    .bottom_grid_pin_0_ ( cbx_1__0__6_bottom_grid_pin_0_ ) , 
    .ccff_tail ( cbx_1__0__6_ccff_tail ) ) ;
cbx_1__0_ cbx_8__0_ (
    .prog_clk ( { ctsbuf_net_1212103 } ) ,
    .chanx_left_in ( sb_1__0__6_chanx_right_out ) , 
    .chanx_right_in ( sb_1__0__7_chanx_left_out ) , 
    .ccff_head ( sb_1__0__7_ccff_tail ) , 
    .chanx_left_out ( cbx_1__0__7_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__0__7_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__0__7_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__0__7_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__0__7_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__0__7_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__0__7_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__0__7_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__0__7_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__0__7_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__0__7_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__0__7_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__0__7_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__0__7_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__0__7_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__0__7_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__0__7_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__0__7_top_grid_pin_31_ ) , 
    .bottom_grid_pin_0_ ( cbx_1__0__7_bottom_grid_pin_0_ ) , 
    .ccff_tail ( cbx_1__0__7_ccff_tail ) ) ;
cbx_1__0_ cbx_9__0_ (
    .prog_clk ( { ctsbuf_net_932075 } ) ,
    .chanx_left_in ( sb_1__0__7_chanx_right_out ) , 
    .chanx_right_in ( sb_1__0__8_chanx_left_out ) , 
    .ccff_head ( sb_1__0__8_ccff_tail ) , 
    .chanx_left_out ( cbx_1__0__8_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__0__8_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__0__8_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__0__8_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__0__8_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__0__8_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__0__8_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__0__8_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__0__8_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__0__8_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__0__8_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__0__8_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__0__8_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__0__8_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__0__8_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__0__8_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__0__8_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__0__8_top_grid_pin_31_ ) , 
    .bottom_grid_pin_0_ ( cbx_1__0__8_bottom_grid_pin_0_ ) , 
    .ccff_tail ( cbx_1__0__8_ccff_tail ) ) ;
cbx_1__0_ cbx_10__0_ (
    .prog_clk ( { ctsbuf_net_692051 } ) ,
    .chanx_left_in ( sb_1__0__8_chanx_right_out ) , 
    .chanx_right_in ( sb_1__0__9_chanx_left_out ) , 
    .ccff_head ( sb_1__0__9_ccff_tail ) , 
    .chanx_left_out ( cbx_1__0__9_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__0__9_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__0__9_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__0__9_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__0__9_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__0__9_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__0__9_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__0__9_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__0__9_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__0__9_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__0__9_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__0__9_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__0__9_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__0__9_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__0__9_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__0__9_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__0__9_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__0__9_top_grid_pin_31_ ) , 
    .bottom_grid_pin_0_ ( cbx_1__0__9_bottom_grid_pin_0_ ) , 
    .ccff_tail ( cbx_1__0__9_ccff_tail ) ) ;
cbx_1__0_ cbx_11__0_ (
    .prog_clk ( { ctsbuf_net_542036 } ) ,
    .chanx_left_in ( sb_1__0__9_chanx_right_out ) , 
    .chanx_right_in ( sb_1__0__10_chanx_left_out ) , 
    .ccff_head ( sb_1__0__10_ccff_tail ) , 
    .chanx_left_out ( cbx_1__0__10_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__0__10_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__0__10_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__0__10_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__0__10_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__0__10_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__0__10_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__0__10_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__0__10_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__0__10_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__0__10_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__0__10_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__0__10_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__0__10_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__0__10_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__0__10_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__0__10_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__0__10_top_grid_pin_31_ ) , 
    .bottom_grid_pin_0_ ( cbx_1__0__10_bottom_grid_pin_0_ ) , 
    .ccff_tail ( cbx_1__0__10_ccff_tail ) ) ;
cbx_1__0_ cbx_12__0_ (
    .prog_clk ( { ctsbuf_net_482030 } ) ,
    .chanx_left_in ( sb_1__0__10_chanx_right_out ) , 
    .chanx_right_in ( sb_12__0__0_chanx_left_out ) , 
    .ccff_head ( sb_12__0__0_ccff_tail ) , 
    .chanx_left_out ( cbx_1__0__11_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__0__11_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__0__11_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__0__11_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__0__11_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__0__11_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__0__11_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__0__11_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__0__11_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__0__11_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__0__11_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__0__11_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__0__11_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__0__11_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__0__11_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__0__11_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__0__11_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__0__11_top_grid_pin_31_ ) , 
    .bottom_grid_pin_0_ ( cbx_1__0__11_bottom_grid_pin_0_ ) , 
    .ccff_tail ( cbx_1__0__11_ccff_tail ) ) ;
cbx_1__1_ cbx_1__1_ (
    .prog_clk ( { ctsbuf_net_4482430 } ) ,
    .chanx_left_in ( sb_0__1__0_chanx_right_out ) , 
    .chanx_right_in ( sb_1__1__0_chanx_left_out ) , 
    .ccff_head ( sb_1__1__0_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__0_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__0_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__0_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__0_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__0_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__0_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__0_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__0_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__0_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__0_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__0_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__0_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__0_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__0_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__0_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__0_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__0_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__0_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__0_ccff_tail ) ) ;
cbx_1__1_ cbx_1__2_ (
    .prog_clk ( { ctsbuf_net_4942476 } ) ,
    .chanx_left_in ( sb_0__1__1_chanx_right_out ) , 
    .chanx_right_in ( sb_1__1__1_chanx_left_out ) , 
    .ccff_head ( sb_1__1__1_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__1_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__1_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__1_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__1_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__1_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__1_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__1_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__1_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__1_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__1_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__1_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__1_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__1_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__1_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__1_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__1_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__1_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__1_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__1_ccff_tail ) ) ;
cbx_1__1_ cbx_1__3_ (
    .prog_clk ( { ctsbuf_net_5212503 } ) ,
    .chanx_left_in ( sb_0__1__2_chanx_right_out ) , 
    .chanx_right_in ( sb_1__1__2_chanx_left_out ) , 
    .ccff_head ( sb_1__1__2_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__2_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__2_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__2_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__2_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__2_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__2_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__2_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__2_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__2_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__2_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__2_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__2_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__2_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__2_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__2_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__2_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__2_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__2_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__2_ccff_tail ) ) ;
cbx_1__1_ cbx_1__4_ (
    .prog_clk ( { ctsbuf_net_5512533 } ) ,
    .chanx_left_in ( sb_0__1__3_chanx_right_out ) , 
    .chanx_right_in ( sb_1__1__3_chanx_left_out ) , 
    .ccff_head ( sb_1__1__3_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__3_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__3_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__3_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__3_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__3_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__3_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__3_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__3_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__3_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__3_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__3_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__3_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__3_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__3_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__3_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__3_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__3_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__3_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__3_ccff_tail ) ) ;
cbx_1__1_ cbx_1__5_ (
    .prog_clk ( { ctsbuf_net_5692551 } ) ,
    .chanx_left_in ( sb_0__1__4_chanx_right_out ) , 
    .chanx_right_in ( sb_1__1__4_chanx_left_out ) , 
    .ccff_head ( sb_1__1__4_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__4_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__4_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__4_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__4_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__4_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__4_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__4_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__4_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__4_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__4_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__4_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__4_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__4_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__4_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__4_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__4_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__4_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__4_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__4_ccff_tail ) ) ;
cbx_1__1_ cbx_1__6_ (
    .prog_clk ( { ctsbuf_net_5802562 } ) ,
    .chanx_left_in ( sb_0__1__5_chanx_right_out ) , 
    .chanx_right_in ( sb_1__1__5_chanx_left_out ) , 
    .ccff_head ( sb_1__1__5_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__5_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__5_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__5_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__5_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__5_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__5_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__5_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__5_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__5_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__5_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__5_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__5_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__5_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__5_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__5_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__5_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__5_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__5_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__5_ccff_tail ) ) ;
cbx_1__1_ cbx_1__7_ (
    .prog_clk ( { ctsbuf_net_5752557 } ) ,
    .chanx_left_in ( sb_0__1__6_chanx_right_out ) , 
    .chanx_right_in ( sb_1__1__6_chanx_left_out ) , 
    .ccff_head ( sb_1__1__6_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__6_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__6_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__6_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__6_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__6_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__6_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__6_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__6_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__6_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__6_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__6_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__6_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__6_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__6_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__6_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__6_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__6_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__6_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__6_ccff_tail ) ) ;
cbx_1__1_ cbx_1__8_ (
    .prog_clk ( { ctsbuf_net_5522534 } ) ,
    .chanx_left_in ( sb_0__1__7_chanx_right_out ) , 
    .chanx_right_in ( sb_1__1__7_chanx_left_out ) , 
    .ccff_head ( sb_1__1__7_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__7_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__7_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__7_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__7_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__7_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__7_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__7_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__7_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__7_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__7_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__7_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__7_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__7_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__7_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__7_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__7_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__7_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__7_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__7_ccff_tail ) ) ;
cbx_1__1_ cbx_1__9_ (
    .prog_clk ( { ctsbuf_net_5392521 } ) ,
    .chanx_left_in ( sb_0__1__8_chanx_right_out ) , 
    .chanx_right_in ( sb_1__1__8_chanx_left_out ) , 
    .ccff_head ( sb_1__1__8_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__8_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__8_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__8_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__8_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__8_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__8_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__8_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__8_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__8_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__8_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__8_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__8_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__8_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__8_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__8_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__8_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__8_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__8_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__8_ccff_tail ) ) ;
cbx_1__1_ cbx_1__10_ (
    .prog_clk ( { ctsbuf_net_4952477 } ) ,
    .chanx_left_in ( sb_0__1__9_chanx_right_out ) , 
    .chanx_right_in ( sb_1__1__9_chanx_left_out ) , 
    .ccff_head ( sb_1__1__9_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__9_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__9_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__9_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__9_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__9_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__9_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__9_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__9_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__9_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__9_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__9_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__9_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__9_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__9_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__9_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__9_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__9_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__9_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__9_ccff_tail ) ) ;
cbx_1__1_ cbx_1__11_ (
    .prog_clk ( { ctsbuf_net_4752457 } ) ,
    .chanx_left_in ( sb_0__1__10_chanx_right_out ) , 
    .chanx_right_in ( sb_1__1__10_chanx_left_out ) , 
    .ccff_head ( sb_1__1__10_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__10_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__10_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__10_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__10_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__10_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__10_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__10_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__10_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__10_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__10_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__10_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__10_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__10_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__10_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__10_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__10_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__10_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__10_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__10_ccff_tail ) ) ;
cbx_1__1_ cbx_2__1_ (
    .prog_clk ( { ctsbuf_net_4042386 } ) ,
    .chanx_left_in ( sb_1__1__0_chanx_right_out ) , 
    .chanx_right_in ( sb_1__1__11_chanx_left_out ) , 
    .ccff_head ( sb_1__1__11_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__11_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__11_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__11_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__11_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__11_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__11_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__11_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__11_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__11_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__11_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__11_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__11_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__11_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__11_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__11_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__11_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__11_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__11_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__11_ccff_tail ) ) ;
cbx_1__1_ cbx_2__2_ (
    .prog_clk ( { ctsbuf_net_4672449 } ) ,
    .chanx_left_in ( sb_1__1__1_chanx_right_out ) , 
    .chanx_right_in ( sb_1__1__12_chanx_left_out ) , 
    .ccff_head ( sb_1__1__12_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__12_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__12_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__12_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__12_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__12_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__12_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__12_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__12_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__12_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__12_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__12_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__12_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__12_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__12_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__12_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__12_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__12_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__12_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__12_ccff_tail ) ) ;
cbx_1__1_ cbx_2__3_ (
    .prog_clk ( { ctsbuf_net_4902472 } ) ,
    .chanx_left_in ( sb_1__1__2_chanx_right_out ) , 
    .chanx_right_in ( sb_1__1__13_chanx_left_out ) , 
    .ccff_head ( sb_1__1__13_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__13_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__13_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__13_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__13_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__13_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__13_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__13_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__13_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__13_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__13_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__13_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__13_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__13_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__13_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__13_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__13_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__13_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__13_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__13_ccff_tail ) ) ;
cbx_1__1_ cbx_2__4_ (
    .prog_clk ( { ctsbuf_net_5342516 } ) ,
    .chanx_left_in ( sb_1__1__3_chanx_right_out ) , 
    .chanx_right_in ( sb_1__1__14_chanx_left_out ) , 
    .ccff_head ( sb_1__1__14_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__14_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__14_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__14_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__14_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__14_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__14_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__14_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__14_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__14_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__14_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__14_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__14_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__14_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__14_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__14_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__14_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__14_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__14_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__14_ccff_tail ) ) ;
cbx_1__1_ cbx_2__5_ (
    .prog_clk ( { ctsbuf_net_5582540 } ) ,
    .chanx_left_in ( sb_1__1__4_chanx_right_out ) , 
    .chanx_right_in ( sb_1__1__15_chanx_left_out ) , 
    .ccff_head ( sb_1__1__15_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__15_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__15_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__15_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__15_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__15_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__15_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__15_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__15_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__15_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__15_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__15_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__15_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__15_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__15_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__15_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__15_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__15_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__15_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__15_ccff_tail ) ) ;
cbx_1__1_ cbx_2__6_ (
    .prog_clk ( { ctsbuf_net_5742556 } ) ,
    .chanx_left_in ( sb_1__1__5_chanx_right_out ) , 
    .chanx_right_in ( sb_1__1__16_chanx_left_out ) , 
    .ccff_head ( sb_1__1__16_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__16_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__16_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__16_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__16_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__16_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__16_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__16_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__16_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__16_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__16_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__16_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__16_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__16_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__16_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__16_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__16_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__16_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__16_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__16_ccff_tail ) ) ;
cbx_1__1_ cbx_2__7_ (
    .prog_clk ( { ctsbuf_net_5622544 } ) ,
    .chanx_left_in ( sb_1__1__6_chanx_right_out ) , 
    .chanx_right_in ( sb_1__1__17_chanx_left_out ) , 
    .ccff_head ( sb_1__1__17_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__17_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__17_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__17_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__17_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__17_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__17_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__17_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__17_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__17_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__17_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__17_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__17_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__17_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__17_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__17_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__17_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__17_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__17_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__17_ccff_tail ) ) ;
cbx_1__1_ cbx_2__8_ (
    .prog_clk ( { ctsbuf_net_5272509 } ) ,
    .chanx_left_in ( sb_1__1__7_chanx_right_out ) , 
    .chanx_right_in ( sb_1__1__18_chanx_left_out ) , 
    .ccff_head ( sb_1__1__18_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__18_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__18_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__18_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__18_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__18_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__18_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__18_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__18_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__18_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__18_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__18_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__18_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__18_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__18_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__18_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__18_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__18_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__18_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__18_ccff_tail ) ) ;
cbx_1__1_ cbx_2__9_ (
    .prog_clk ( { ctsbuf_net_5112493 } ) ,
    .chanx_left_in ( sb_1__1__8_chanx_right_out ) , 
    .chanx_right_in ( sb_1__1__19_chanx_left_out ) , 
    .ccff_head ( sb_1__1__19_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__19_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__19_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__19_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__19_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__19_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__19_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__19_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__19_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__19_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__19_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__19_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__19_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__19_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__19_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__19_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__19_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__19_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__19_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__19_ccff_tail ) ) ;
cbx_1__1_ cbx_2__10_ (
    .prog_clk ( { ctsbuf_net_4562438 } ) ,
    .chanx_left_in ( sb_1__1__9_chanx_right_out ) , 
    .chanx_right_in ( sb_1__1__20_chanx_left_out ) , 
    .ccff_head ( sb_1__1__20_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__20_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__20_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__20_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__20_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__20_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__20_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__20_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__20_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__20_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__20_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__20_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__20_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__20_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__20_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__20_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__20_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__20_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__20_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__20_ccff_tail ) ) ;
cbx_1__1_ cbx_2__11_ (
    .prog_clk ( { ctsbuf_net_4342416 } ) ,
    .chanx_left_in ( sb_1__1__10_chanx_right_out ) , 
    .chanx_right_in ( sb_1__1__21_chanx_left_out ) , 
    .ccff_head ( sb_1__1__21_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__21_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__21_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__21_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__21_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__21_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__21_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__21_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__21_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__21_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__21_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__21_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__21_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__21_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__21_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__21_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__21_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__21_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__21_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__21_ccff_tail ) ) ;
cbx_1__1_ cbx_3__1_ (
    .prog_clk ( { ctsbuf_net_3612343 } ) ,
    .chanx_left_in ( sb_1__1__11_chanx_right_out ) , 
    .chanx_right_in ( sb_1__1__22_chanx_left_out ) , 
    .ccff_head ( sb_1__1__22_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__22_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__22_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__22_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__22_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__22_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__22_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__22_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__22_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__22_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__22_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__22_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__22_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__22_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__22_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__22_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__22_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__22_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__22_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__22_ccff_tail ) ) ;
cbx_1__1_ cbx_3__2_ (
    .prog_clk ( { ctsbuf_net_4252407 } ) ,
    .chanx_left_in ( sb_1__1__12_chanx_right_out ) , 
    .chanx_right_in ( sb_1__1__23_chanx_left_out ) , 
    .ccff_head ( sb_1__1__23_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__23_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__23_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__23_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__23_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__23_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__23_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__23_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__23_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__23_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__23_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__23_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__23_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__23_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__23_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__23_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__23_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__23_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__23_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__23_ccff_tail ) ) ;
cbx_1__1_ cbx_3__3_ (
    .prog_clk ( { ctsbuf_net_4502432 } ) ,
    .chanx_left_in ( sb_1__1__13_chanx_right_out ) , 
    .chanx_right_in ( sb_1__1__24_chanx_left_out ) , 
    .ccff_head ( sb_1__1__24_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__24_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__24_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__24_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__24_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__24_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__24_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__24_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__24_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__24_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__24_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__24_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__24_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__24_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__24_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__24_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__24_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__24_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__24_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__24_ccff_tail ) ) ;
cbx_1__1_ cbx_3__4_ (
    .prog_clk ( { ctsbuf_net_5062488 } ) ,
    .chanx_left_in ( sb_1__1__14_chanx_right_out ) , 
    .chanx_right_in ( sb_1__1__25_chanx_left_out ) , 
    .ccff_head ( sb_1__1__25_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__25_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__25_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__25_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__25_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__25_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__25_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__25_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__25_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__25_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__25_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__25_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__25_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__25_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__25_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__25_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__25_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__25_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__25_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__25_ccff_tail ) ) ;
cbx_1__1_ cbx_3__5_ (
    .prog_clk ( { ctsbuf_net_5362518 } ) ,
    .chanx_left_in ( sb_1__1__15_chanx_right_out ) , 
    .chanx_right_in ( sb_1__1__26_chanx_left_out ) , 
    .ccff_head ( sb_1__1__26_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__26_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__26_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__26_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__26_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__26_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__26_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__26_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__26_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__26_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__26_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__26_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__26_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__26_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__26_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__26_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__26_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__26_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__26_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__26_ccff_tail ) ) ;
cbx_1__1_ cbx_3__6_ (
    .prog_clk ( { ctsbuf_net_5602542 } ) ,
    .chanx_left_in ( sb_1__1__16_chanx_right_out ) , 
    .chanx_right_in ( sb_1__1__27_chanx_left_out ) , 
    .ccff_head ( sb_1__1__27_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__27_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__27_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__27_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__27_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__27_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__27_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__27_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__27_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__27_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__27_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__27_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__27_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__27_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__27_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__27_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__27_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__27_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__27_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__27_ccff_tail ) ) ;
cbx_1__1_ cbx_3__7_ (
    .prog_clk ( { ctsbuf_net_5422524 } ) ,
    .chanx_left_in ( sb_1__1__17_chanx_right_out ) , 
    .chanx_right_in ( sb_1__1__28_chanx_left_out ) , 
    .ccff_head ( sb_1__1__28_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__28_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__28_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__28_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__28_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__28_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__28_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__28_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__28_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__28_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__28_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__28_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__28_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__28_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__28_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__28_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__28_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__28_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__28_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__28_ccff_tail ) ) ;
cbx_1__1_ cbx_3__8_ (
    .prog_clk ( { ctsbuf_net_4972479 } ) ,
    .chanx_left_in ( sb_1__1__18_chanx_right_out ) , 
    .chanx_right_in ( sb_1__1__29_chanx_left_out ) , 
    .ccff_head ( sb_1__1__29_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__29_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__29_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__29_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__29_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__29_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__29_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__29_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__29_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__29_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__29_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__29_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__29_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__29_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__29_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__29_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__29_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__29_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__29_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__29_ccff_tail ) ) ;
cbx_1__1_ cbx_3__9_ (
    .prog_clk ( { p_abuf20 } ) ,
    .chanx_left_in ( sb_1__1__19_chanx_right_out ) , 
    .chanx_right_in ( sb_1__1__30_chanx_left_out ) , 
    .ccff_head ( sb_1__1__30_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__30_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__30_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__30_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__30_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__30_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__30_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__30_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__30_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__30_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__30_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__30_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__30_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__30_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__30_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__30_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__30_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__30_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__30_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__30_ccff_tail ) ) ;
cbx_1__1_ cbx_3__10_ (
    .prog_clk ( { ctsbuf_net_4122394 } ) ,
    .chanx_left_in ( sb_1__1__20_chanx_right_out ) , 
    .chanx_right_in ( sb_1__1__31_chanx_left_out ) , 
    .ccff_head ( sb_1__1__31_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__31_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__31_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__31_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__31_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__31_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__31_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__31_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__31_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__31_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__31_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__31_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__31_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__31_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__31_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__31_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__31_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__31_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__31_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__31_ccff_tail ) ) ;
cbx_1__1_ cbx_3__11_ (
    .prog_clk ( { ctsbuf_net_3902372 } ) ,
    .chanx_left_in ( sb_1__1__21_chanx_right_out ) , 
    .chanx_right_in ( sb_1__1__32_chanx_left_out ) , 
    .ccff_head ( sb_1__1__32_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__32_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__32_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__32_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__32_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__32_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__32_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__32_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__32_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__32_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__32_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__32_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__32_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__32_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__32_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__32_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__32_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__32_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__32_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__32_ccff_tail ) ) ;
cbx_1__1_ cbx_4__1_ (
    .prog_clk ( { ctsbuf_net_3172299 } ) ,
    .chanx_left_in ( sb_1__1__22_chanx_right_out ) , 
    .chanx_right_in ( sb_1__1__33_chanx_left_out ) , 
    .ccff_head ( sb_1__1__33_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__33_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__33_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__33_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__33_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__33_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__33_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__33_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__33_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__33_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__33_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__33_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__33_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__33_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__33_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__33_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__33_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__33_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__33_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__33_ccff_tail ) ) ;
cbx_1__1_ cbx_4__2_ (
    .prog_clk ( { ctsbuf_net_3812363 } ) ,
    .chanx_left_in ( sb_1__1__23_chanx_right_out ) , 
    .chanx_right_in ( sb_1__1__34_chanx_left_out ) , 
    .ccff_head ( sb_1__1__34_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__34_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__34_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__34_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__34_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__34_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__34_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__34_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__34_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__34_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__34_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__34_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__34_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__34_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__34_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__34_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__34_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__34_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__34_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__34_ccff_tail ) ) ;
cbx_1__1_ cbx_4__3_ (
    .prog_clk ( { ctsbuf_net_4062388 } ) ,
    .chanx_left_in ( sb_1__1__24_chanx_right_out ) , 
    .chanx_right_in ( sb_1__1__35_chanx_left_out ) , 
    .ccff_head ( sb_1__1__35_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__35_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__35_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__35_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__35_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__35_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__35_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__35_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__35_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__35_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__35_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__35_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__35_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__35_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__35_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__35_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__35_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__35_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__35_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__35_ccff_tail ) ) ;
cbx_1__1_ cbx_4__4_ (
    .prog_clk ( { ctsbuf_net_4702452 } ) ,
    .chanx_left_in ( sb_1__1__25_chanx_right_out ) , 
    .chanx_right_in ( sb_1__1__36_chanx_left_out ) , 
    .ccff_head ( sb_1__1__36_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__36_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__36_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__36_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__36_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__36_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__36_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__36_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__36_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__36_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__36_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__36_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__36_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__36_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__36_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__36_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__36_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__36_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__36_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__36_ccff_tail ) ) ;
cbx_1__1_ cbx_4__5_ (
    .prog_clk ( { ctsbuf_net_4922474 } ) ,
    .chanx_left_in ( sb_1__1__26_chanx_right_out ) , 
    .chanx_right_in ( sb_1__1__37_chanx_left_out ) , 
    .ccff_head ( sb_1__1__37_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__37_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__37_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__37_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__37_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__37_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__37_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__37_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__37_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__37_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__37_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__37_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__37_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__37_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__37_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__37_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__37_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__37_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__37_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__37_ccff_tail ) ) ;
cbx_1__1_ cbx_4__6_ (
    .prog_clk ( { ctsbuf_net_5382520 } ) ,
    .chanx_left_in ( sb_1__1__27_chanx_right_out ) , 
    .chanx_right_in ( sb_1__1__38_chanx_left_out ) , 
    .ccff_head ( sb_1__1__38_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__38_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__38_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__38_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__38_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__38_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__38_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__38_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__38_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__38_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__38_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__38_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__38_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__38_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__38_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__38_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__38_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__38_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__38_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__38_ccff_tail ) ) ;
cbx_1__1_ cbx_4__7_ (
    .prog_clk ( { ctsbuf_net_5142496 } ) ,
    .chanx_left_in ( sb_1__1__28_chanx_right_out ) , 
    .chanx_right_in ( sb_1__1__39_chanx_left_out ) , 
    .ccff_head ( sb_1__1__39_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__39_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__39_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__39_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__39_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__39_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__39_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__39_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__39_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__39_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__39_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__39_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__39_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__39_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__39_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__39_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__39_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__39_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__39_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__39_ccff_tail ) ) ;
cbx_1__1_ cbx_4__8_ (
    .prog_clk ( { ctsbuf_net_4582440 } ) ,
    .chanx_left_in ( sb_1__1__29_chanx_right_out ) , 
    .chanx_right_in ( sb_1__1__40_chanx_left_out ) , 
    .ccff_head ( sb_1__1__40_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__40_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__40_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__40_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__40_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__40_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__40_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__40_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__40_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__40_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__40_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__40_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__40_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__40_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__40_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__40_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__40_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__40_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__40_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__40_ccff_tail ) ) ;
cbx_1__1_ cbx_4__9_ (
    .prog_clk ( { ctsbuf_net_4372419 } ) ,
    .chanx_left_in ( sb_1__1__30_chanx_right_out ) , 
    .chanx_right_in ( sb_1__1__41_chanx_left_out ) , 
    .ccff_head ( sb_1__1__41_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__41_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__41_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__41_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__41_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__41_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__41_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__41_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__41_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__41_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__41_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__41_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__41_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__41_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__41_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__41_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__41_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__41_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__41_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__41_ccff_tail ) ) ;
cbx_1__1_ cbx_4__10_ (
    .prog_clk ( { ctsbuf_net_3692351 } ) ,
    .chanx_left_in ( sb_1__1__31_chanx_right_out ) , 
    .chanx_right_in ( sb_1__1__42_chanx_left_out ) , 
    .ccff_head ( sb_1__1__42_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__42_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__42_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__42_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__42_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__42_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__42_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__42_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__42_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__42_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__42_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__42_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__42_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__42_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__42_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__42_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__42_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__42_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__42_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__42_ccff_tail ) ) ;
cbx_1__1_ cbx_4__11_ (
    .prog_clk ( { ctsbuf_net_3472329 } ) ,
    .chanx_left_in ( sb_1__1__32_chanx_right_out ) , 
    .chanx_right_in ( sb_1__1__43_chanx_left_out ) , 
    .ccff_head ( sb_1__1__43_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__43_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__43_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__43_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__43_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__43_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__43_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__43_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__43_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__43_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__43_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__43_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__43_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__43_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__43_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__43_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__43_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__43_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__43_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__43_ccff_tail ) ) ;
cbx_1__1_ cbx_5__1_ (
    .prog_clk ( { ctsbuf_net_2722254 } ) ,
    .chanx_left_in ( sb_1__1__33_chanx_right_out ) , 
    .chanx_right_in ( sb_1__1__44_chanx_left_out ) , 
    .ccff_head ( sb_1__1__44_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__44_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__44_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__44_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__44_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__44_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__44_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__44_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__44_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__44_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__44_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__44_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__44_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__44_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__44_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__44_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__44_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__44_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__44_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__44_ccff_tail ) ) ;
cbx_1__1_ cbx_5__2_ (
    .prog_clk ( { ctsbuf_net_3382320 } ) ,
    .chanx_left_in ( sb_1__1__34_chanx_right_out ) , 
    .chanx_right_in ( sb_1__1__45_chanx_left_out ) , 
    .ccff_head ( sb_1__1__45_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__45_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__45_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__45_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__45_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__45_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__45_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__45_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__45_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__45_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__45_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__45_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__45_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__45_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__45_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__45_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__45_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__45_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__45_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__45_ccff_tail ) ) ;
cbx_1__1_ cbx_5__3_ (
    .prog_clk ( { ctsbuf_net_3632345 } ) ,
    .chanx_left_in ( sb_1__1__35_chanx_right_out ) , 
    .chanx_right_in ( sb_1__1__46_chanx_left_out ) , 
    .ccff_head ( sb_1__1__46_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__46_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__46_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__46_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__46_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__46_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__46_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__46_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__46_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__46_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__46_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__46_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__46_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__46_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__46_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__46_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__46_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__46_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__46_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__46_ccff_tail ) ) ;
cbx_1__1_ cbx_5__4_ (
    .prog_clk ( { ctsbuf_net_4282410 } ) ,
    .chanx_left_in ( sb_1__1__36_chanx_right_out ) , 
    .chanx_right_in ( sb_1__1__47_chanx_left_out ) , 
    .ccff_head ( sb_1__1__47_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__47_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__47_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__47_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__47_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__47_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__47_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__47_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__47_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__47_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__47_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__47_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__47_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__47_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__47_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__47_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__47_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__47_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__47_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__47_ccff_tail ) ) ;
cbx_1__1_ cbx_5__5_ (
    .prog_clk ( { ctsbuf_net_4722454 } ) ,
    .chanx_left_in ( sb_1__1__37_chanx_right_out ) , 
    .chanx_right_in ( sb_1__1__48_chanx_left_out ) , 
    .ccff_head ( sb_1__1__48_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__48_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__48_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__48_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__48_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__48_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__48_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__48_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__48_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__48_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__48_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__48_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__48_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__48_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__48_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__48_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__48_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__48_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__48_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__48_ccff_tail ) ) ;
cbx_1__1_ cbx_5__6_ (
    .prog_clk ( { ctsbuf_net_5092491 } ) ,
    .chanx_left_in ( sb_1__1__38_chanx_right_out ) , 
    .chanx_right_in ( sb_1__1__49_chanx_left_out ) , 
    .ccff_head ( sb_1__1__49_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__49_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__49_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__49_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__49_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__49_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__49_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__49_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__49_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__49_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__49_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__49_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__49_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__49_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__49_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__49_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__49_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__49_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__49_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__49_ccff_tail ) ) ;
cbx_1__1_ cbx_5__7_ (
    .prog_clk ( { ctsbuf_net_4812463 } ) ,
    .chanx_left_in ( sb_1__1__39_chanx_right_out ) , 
    .chanx_right_in ( sb_1__1__50_chanx_left_out ) , 
    .ccff_head ( sb_1__1__50_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__50_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__50_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__50_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__50_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__50_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__50_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__50_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__50_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__50_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__50_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__50_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__50_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__50_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__50_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__50_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__50_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__50_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__50_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__50_ccff_tail ) ) ;
cbx_1__1_ cbx_5__8_ (
    .prog_clk ( { ctsbuf_net_4142396 } ) ,
    .chanx_left_in ( sb_1__1__40_chanx_right_out ) , 
    .chanx_right_in ( sb_1__1__51_chanx_left_out ) , 
    .ccff_head ( sb_1__1__51_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__51_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__51_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__51_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__51_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__51_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__51_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__51_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__51_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__51_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__51_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__51_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__51_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__51_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__51_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__51_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__51_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__51_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__51_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__51_ccff_tail ) ) ;
cbx_1__1_ cbx_5__9_ (
    .prog_clk ( { ctsbuf_net_3932375 } ) ,
    .chanx_left_in ( sb_1__1__41_chanx_right_out ) , 
    .chanx_right_in ( sb_1__1__52_chanx_left_out ) , 
    .ccff_head ( sb_1__1__52_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__52_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__52_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__52_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__52_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__52_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__52_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__52_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__52_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__52_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__52_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__52_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__52_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__52_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__52_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__52_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__52_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__52_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__52_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__52_ccff_tail ) ) ;
cbx_1__1_ cbx_5__10_ (
    .prog_clk ( { ctsbuf_net_3252307 } ) ,
    .chanx_left_in ( sb_1__1__42_chanx_right_out ) , 
    .chanx_right_in ( sb_1__1__53_chanx_left_out ) , 
    .ccff_head ( sb_1__1__53_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__53_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__53_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__53_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__53_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__53_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__53_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__53_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__53_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__53_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__53_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__53_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__53_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__53_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__53_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__53_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__53_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__53_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__53_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__53_ccff_tail ) ) ;
cbx_1__1_ cbx_5__11_ (
    .prog_clk ( { ctsbuf_net_3022284 } ) ,
    .chanx_left_in ( sb_1__1__43_chanx_right_out ) , 
    .chanx_right_in ( sb_1__1__54_chanx_left_out ) , 
    .ccff_head ( sb_1__1__54_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__54_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__54_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__54_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__54_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__54_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__54_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__54_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__54_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__54_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__54_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__54_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__54_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__54_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__54_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__54_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__54_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__54_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__54_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__54_ccff_tail ) ) ;
cbx_1__1_ cbx_6__1_ (
    .prog_clk ( { ctsbuf_net_2272209 } ) ,
    .chanx_left_in ( sb_1__1__44_chanx_right_out ) , 
    .chanx_right_in ( sb_1__1__55_chanx_left_out ) , 
    .ccff_head ( sb_1__1__55_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__55_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__55_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__55_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__55_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__55_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__55_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__55_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__55_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__55_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__55_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__55_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__55_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__55_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__55_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__55_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__55_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__55_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__55_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__55_ccff_tail ) ) ;
cbx_1__1_ cbx_6__2_ (
    .prog_clk ( { ctsbuf_net_2922274 } ) ,
    .chanx_left_in ( sb_1__1__45_chanx_right_out ) , 
    .chanx_right_in ( sb_1__1__56_chanx_left_out ) , 
    .ccff_head ( sb_1__1__56_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__56_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__56_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__56_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__56_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__56_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__56_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__56_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__56_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__56_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__56_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__56_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__56_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__56_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__56_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__56_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__56_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__56_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__56_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__56_ccff_tail ) ) ;
cbx_1__1_ cbx_6__3_ (
    .prog_clk ( { p_abuf14 } ) ,
    .chanx_left_in ( sb_1__1__46_chanx_right_out ) , 
    .chanx_right_in ( sb_1__1__57_chanx_left_out ) , 
    .ccff_head ( sb_1__1__57_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__57_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__57_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__57_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__57_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__57_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__57_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__57_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__57_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__57_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__57_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__57_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__57_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__57_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__57_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__57_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__57_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__57_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__57_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__57_ccff_tail ) ) ;
cbx_1__1_ cbx_6__4_ (
    .prog_clk ( { ctsbuf_net_3842366 } ) ,
    .chanx_left_in ( sb_1__1__47_chanx_right_out ) , 
    .chanx_right_in ( sb_1__1__58_chanx_left_out ) , 
    .ccff_head ( sb_1__1__58_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__58_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__58_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__58_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__58_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__58_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__58_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__58_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__58_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__58_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__58_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__58_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__58_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__58_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__58_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__58_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__58_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__58_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__58_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__58_ccff_tail ) ) ;
cbx_1__1_ cbx_6__5_ (
    .prog_clk ( { ctsbuf_net_4302412 } ) ,
    .chanx_left_in ( sb_1__1__48_chanx_right_out ) , 
    .chanx_right_in ( sb_1__1__59_chanx_left_out ) , 
    .ccff_head ( sb_1__1__59_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__59_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__59_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__59_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__59_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__59_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__59_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__59_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__59_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__59_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__59_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__59_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__59_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__59_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__59_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__59_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__59_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__59_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__59_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__59_ccff_tail ) ) ;
cbx_1__1_ cbx_6__6_ (
    .prog_clk ( { ctsbuf_net_4742456 } ) ,
    .chanx_left_in ( sb_1__1__49_chanx_right_out ) , 
    .chanx_right_in ( sb_1__1__60_chanx_left_out ) , 
    .ccff_head ( sb_1__1__60_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__60_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__60_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__60_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__60_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__60_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__60_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__60_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__60_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__60_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__60_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__60_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__60_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__60_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__60_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__60_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__60_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__60_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__60_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__60_ccff_tail ) ) ;
cbx_1__1_ cbx_6__7_ (
    .prog_clk ( { ctsbuf_net_4402422 } ) ,
    .chanx_left_in ( sb_1__1__50_chanx_right_out ) , 
    .chanx_right_in ( sb_1__1__61_chanx_left_out ) , 
    .ccff_head ( sb_1__1__61_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__61_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__61_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__61_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__61_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__61_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__61_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__61_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__61_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__61_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__61_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__61_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__61_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__61_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__61_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__61_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__61_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__61_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__61_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__61_ccff_tail ) ) ;
cbx_1__1_ cbx_6__8_ (
    .prog_clk ( { ctsbuf_net_3712353 } ) ,
    .chanx_left_in ( sb_1__1__51_chanx_right_out ) , 
    .chanx_right_in ( sb_1__1__62_chanx_left_out ) , 
    .ccff_head ( sb_1__1__62_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__62_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__62_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__62_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__62_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__62_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__62_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__62_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__62_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__62_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__62_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__62_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__62_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__62_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__62_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__62_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__62_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__62_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__62_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__62_ccff_tail ) ) ;
cbx_1__1_ cbx_6__9_ (
    .prog_clk ( { p_abuf17 } ) ,
    .chanx_left_in ( sb_1__1__52_chanx_right_out ) , 
    .chanx_right_in ( sb_1__1__63_chanx_left_out ) , 
    .ccff_head ( sb_1__1__63_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__63_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__63_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__63_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__63_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__63_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__63_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__63_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__63_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__63_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__63_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__63_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__63_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__63_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__63_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__63_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__63_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__63_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__63_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__63_ccff_tail ) ) ;
cbx_1__1_ cbx_6__10_ (
    .prog_clk ( { ctsbuf_net_2802262 } ) ,
    .chanx_left_in ( sb_1__1__53_chanx_right_out ) , 
    .chanx_right_in ( sb_1__1__64_chanx_left_out ) , 
    .ccff_head ( sb_1__1__64_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__64_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__64_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__64_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__64_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__64_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__64_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__64_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__64_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__64_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__64_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__64_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__64_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__64_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__64_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__64_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__64_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__64_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__64_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__64_ccff_tail ) ) ;
cbx_1__1_ cbx_6__11_ (
    .prog_clk ( { ctsbuf_net_2572239 } ) ,
    .chanx_left_in ( sb_1__1__54_chanx_right_out ) , 
    .chanx_right_in ( sb_1__1__65_chanx_left_out ) , 
    .ccff_head ( sb_1__1__65_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__65_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__65_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__65_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__65_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__65_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__65_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__65_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__65_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__65_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__65_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__65_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__65_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__65_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__65_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__65_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__65_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__65_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__65_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__65_ccff_tail ) ) ;
cbx_1__1_ cbx_7__1_ (
    .prog_clk ( { ctsbuf_net_1832165 } ) ,
    .chanx_left_in ( sb_1__1__55_chanx_right_out ) , 
    .chanx_right_in ( sb_1__1__66_chanx_left_out ) , 
    .ccff_head ( sb_1__1__66_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__66_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__66_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__66_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__66_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__66_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__66_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__66_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__66_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__66_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__66_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__66_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__66_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__66_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__66_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__66_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__66_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__66_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__66_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__66_ccff_tail ) ) ;
cbx_1__1_ cbx_7__2_ (
    .prog_clk ( { ctsbuf_net_2482230 } ) ,
    .chanx_left_in ( sb_1__1__56_chanx_right_out ) , 
    .chanx_right_in ( sb_1__1__67_chanx_left_out ) , 
    .ccff_head ( sb_1__1__67_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__67_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__67_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__67_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__67_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__67_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__67_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__67_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__67_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__67_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__67_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__67_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__67_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__67_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__67_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__67_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__67_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__67_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__67_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__67_ccff_tail ) ) ;
cbx_1__1_ cbx_7__3_ (
    .prog_clk ( { ctsbuf_net_2742256 } ) ,
    .chanx_left_in ( sb_1__1__57_chanx_right_out ) , 
    .chanx_right_in ( sb_1__1__68_chanx_left_out ) , 
    .ccff_head ( sb_1__1__68_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__68_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__68_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__68_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__68_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__68_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__68_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__68_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__68_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__68_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__68_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__68_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__68_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__68_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__68_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__68_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__68_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__68_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__68_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__68_ccff_tail ) ) ;
cbx_1__1_ cbx_7__4_ (
    .prog_clk ( { ctsbuf_net_3412323 } ) ,
    .chanx_left_in ( sb_1__1__58_chanx_right_out ) , 
    .chanx_right_in ( sb_1__1__69_chanx_left_out ) , 
    .ccff_head ( sb_1__1__69_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__69_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__69_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__69_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__69_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__69_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__69_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__69_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__69_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__69_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__69_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__69_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__69_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__69_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__69_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__69_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__69_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__69_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__69_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__69_ccff_tail ) ) ;
cbx_1__1_ cbx_7__5_ (
    .prog_clk ( { ctsbuf_net_3652347 } ) ,
    .chanx_left_in ( sb_1__1__59_chanx_right_out ) , 
    .chanx_right_in ( sb_1__1__70_chanx_left_out ) , 
    .ccff_head ( sb_1__1__70_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__70_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__70_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__70_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__70_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__70_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__70_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__70_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__70_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__70_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__70_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__70_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__70_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__70_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__70_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__70_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__70_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__70_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__70_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__70_ccff_tail ) ) ;
cbx_1__1_ cbx_7__6_ (
    .prog_clk ( { ctsbuf_net_4322414 } ) ,
    .chanx_left_in ( sb_1__1__60_chanx_right_out ) , 
    .chanx_right_in ( sb_1__1__71_chanx_left_out ) , 
    .ccff_head ( sb_1__1__71_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__71_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__71_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__71_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__71_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__71_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__71_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__71_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__71_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__71_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__71_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__71_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__71_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__71_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__71_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__71_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__71_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__71_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__71_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__71_ccff_tail ) ) ;
cbx_1__1_ cbx_7__7_ (
    .prog_clk ( { ctsbuf_net_3962378 } ) ,
    .chanx_left_in ( sb_1__1__61_chanx_right_out ) , 
    .chanx_right_in ( sb_1__1__72_chanx_left_out ) , 
    .ccff_head ( sb_1__1__72_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__72_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__72_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__72_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__72_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__72_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__72_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__72_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__72_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__72_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__72_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__72_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__72_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__72_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__72_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__72_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__72_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__72_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__72_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__72_ccff_tail ) ) ;
cbx_1__1_ cbx_7__8_ (
    .prog_clk ( { ctsbuf_net_3272309 } ) ,
    .chanx_left_in ( sb_1__1__62_chanx_right_out ) , 
    .chanx_right_in ( sb_1__1__73_chanx_left_out ) , 
    .ccff_head ( sb_1__1__73_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__73_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__73_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__73_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__73_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__73_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__73_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__73_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__73_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__73_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__73_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__73_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__73_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__73_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__73_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__73_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__73_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__73_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__73_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__73_ccff_tail ) ) ;
cbx_1__1_ cbx_7__9_ (
    .prog_clk ( { ctsbuf_net_3052287 } ) ,
    .chanx_left_in ( sb_1__1__63_chanx_right_out ) , 
    .chanx_right_in ( sb_1__1__74_chanx_left_out ) , 
    .ccff_head ( sb_1__1__74_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__74_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__74_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__74_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__74_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__74_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__74_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__74_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__74_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__74_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__74_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__74_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__74_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__74_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__74_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__74_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__74_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__74_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__74_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__74_ccff_tail ) ) ;
cbx_1__1_ cbx_7__10_ (
    .prog_clk ( { ctsbuf_net_2352217 } ) ,
    .chanx_left_in ( sb_1__1__64_chanx_right_out ) , 
    .chanx_right_in ( sb_1__1__75_chanx_left_out ) , 
    .ccff_head ( sb_1__1__75_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__75_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__75_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__75_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__75_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__75_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__75_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__75_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__75_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__75_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__75_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__75_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__75_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__75_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__75_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__75_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__75_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__75_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__75_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__75_ccff_tail ) ) ;
cbx_1__1_ cbx_7__11_ (
    .prog_clk ( { ctsbuf_net_2122194 } ) ,
    .chanx_left_in ( sb_1__1__65_chanx_right_out ) , 
    .chanx_right_in ( sb_1__1__76_chanx_left_out ) , 
    .ccff_head ( sb_1__1__76_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__76_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__76_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__76_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__76_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__76_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__76_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__76_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__76_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__76_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__76_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__76_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__76_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__76_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__76_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__76_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__76_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__76_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__76_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__76_ccff_tail ) ) ;
cbx_1__1_ cbx_8__1_ (
    .prog_clk ( { ctsbuf_net_1442126 } ) ,
    .chanx_left_in ( sb_1__1__66_chanx_right_out ) , 
    .chanx_right_in ( sb_1__1__77_chanx_left_out ) , 
    .ccff_head ( sb_1__1__77_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__77_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__77_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__77_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__77_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__77_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__77_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__77_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__77_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__77_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__77_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__77_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__77_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__77_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__77_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__77_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__77_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__77_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__77_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__77_ccff_tail ) ) ;
cbx_1__1_ cbx_8__2_ (
    .prog_clk ( { ctsbuf_net_2022184 } ) ,
    .chanx_left_in ( sb_1__1__67_chanx_right_out ) , 
    .chanx_right_in ( sb_1__1__78_chanx_left_out ) , 
    .ccff_head ( sb_1__1__78_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__78_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__78_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__78_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__78_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__78_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__78_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__78_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__78_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__78_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__78_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__78_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__78_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__78_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__78_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__78_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__78_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__78_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__78_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__78_ccff_tail ) ) ;
cbx_1__1_ cbx_8__3_ (
    .prog_clk ( { ctsbuf_net_2292211 } ) ,
    .chanx_left_in ( sb_1__1__68_chanx_right_out ) , 
    .chanx_right_in ( sb_1__1__79_chanx_left_out ) , 
    .ccff_head ( sb_1__1__79_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__79_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__79_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__79_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__79_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__79_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__79_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__79_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__79_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__79_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__79_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__79_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__79_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__79_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__79_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__79_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__79_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__79_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__79_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__79_ccff_tail ) ) ;
cbx_1__1_ cbx_8__4_ (
    .prog_clk ( { ctsbuf_net_2952277 } ) ,
    .chanx_left_in ( sb_1__1__69_chanx_right_out ) , 
    .chanx_right_in ( sb_1__1__80_chanx_left_out ) , 
    .ccff_head ( sb_1__1__80_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__80_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__80_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__80_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__80_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__80_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__80_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__80_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__80_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__80_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__80_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__80_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__80_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__80_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__80_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__80_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__80_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__80_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__80_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__80_ccff_tail ) ) ;
cbx_1__1_ cbx_8__5_ (
    .prog_clk ( { ctsbuf_net_3432325 } ) ,
    .chanx_left_in ( sb_1__1__70_chanx_right_out ) , 
    .chanx_right_in ( sb_1__1__81_chanx_left_out ) , 
    .ccff_head ( sb_1__1__81_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__81_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__81_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__81_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__81_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__81_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__81_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__81_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__81_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__81_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__81_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__81_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__81_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__81_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__81_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__81_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__81_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__81_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__81_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__81_ccff_tail ) ) ;
cbx_1__1_ cbx_8__6_ (
    .prog_clk ( { ctsbuf_net_3872369 } ) ,
    .chanx_left_in ( sb_1__1__71_chanx_right_out ) , 
    .chanx_right_in ( sb_1__1__82_chanx_left_out ) , 
    .ccff_head ( sb_1__1__82_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__82_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__82_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__82_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__82_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__82_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__82_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__82_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__82_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__82_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__82_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__82_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__82_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__82_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__82_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__82_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__82_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__82_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__82_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__82_ccff_tail ) ) ;
cbx_1__1_ cbx_8__7_ (
    .prog_clk ( { ctsbuf_net_3532335 } ) ,
    .chanx_left_in ( sb_1__1__72_chanx_right_out ) , 
    .chanx_right_in ( sb_1__1__83_chanx_left_out ) , 
    .ccff_head ( sb_1__1__83_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__83_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__83_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__83_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__83_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__83_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__83_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__83_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__83_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__83_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__83_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__83_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__83_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__83_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__83_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__83_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__83_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__83_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__83_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__83_ccff_tail ) ) ;
cbx_1__1_ cbx_8__8_ (
    .prog_clk ( { ctsbuf_net_3072289 } ) ,
    .chanx_left_in ( sb_1__1__73_chanx_right_out ) , 
    .chanx_right_in ( sb_1__1__84_chanx_left_out ) , 
    .ccff_head ( sb_1__1__84_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__84_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__84_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__84_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__84_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__84_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__84_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__84_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__84_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__84_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__84_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__84_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__84_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__84_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__84_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__84_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__84_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__84_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__84_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__84_ccff_tail ) ) ;
cbx_1__1_ cbx_8__9_ (
    .prog_clk ( { ctsbuf_net_2602242 } ) ,
    .chanx_left_in ( sb_1__1__74_chanx_right_out ) , 
    .chanx_right_in ( sb_1__1__85_chanx_left_out ) , 
    .ccff_head ( sb_1__1__85_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__85_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__85_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__85_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__85_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__85_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__85_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__85_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__85_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__85_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__85_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__85_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__85_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__85_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__85_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__85_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__85_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__85_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__85_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__85_ccff_tail ) ) ;
cbx_1__1_ cbx_8__10_ (
    .prog_clk ( { ctsbuf_net_2142196 } ) ,
    .chanx_left_in ( sb_1__1__75_chanx_right_out ) , 
    .chanx_right_in ( sb_1__1__86_chanx_left_out ) , 
    .ccff_head ( sb_1__1__86_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__86_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__86_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__86_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__86_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__86_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__86_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__86_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__86_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__86_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__86_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__86_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__86_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__86_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__86_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__86_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__86_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__86_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__86_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__86_ccff_tail ) ) ;
cbx_1__1_ cbx_8__11_ (
    .prog_clk ( { ctsbuf_net_1682150 } ) ,
    .chanx_left_in ( sb_1__1__76_chanx_right_out ) , 
    .chanx_right_in ( sb_1__1__87_chanx_left_out ) , 
    .ccff_head ( sb_1__1__87_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__87_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__87_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__87_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__87_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__87_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__87_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__87_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__87_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__87_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__87_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__87_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__87_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__87_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__87_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__87_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__87_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__87_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__87_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__87_ccff_tail ) ) ;
cbx_1__1_ cbx_9__1_ (
    .prog_clk ( { ctsbuf_net_1122094 } ) ,
    .chanx_left_in ( sb_1__1__77_chanx_right_out ) , 
    .chanx_right_in ( sb_1__1__88_chanx_left_out ) , 
    .ccff_head ( sb_1__1__88_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__88_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__88_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__88_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__88_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__88_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__88_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__88_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__88_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__88_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__88_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__88_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__88_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__88_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__88_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__88_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__88_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__88_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__88_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__88_ccff_tail ) ) ;
cbx_1__1_ cbx_9__2_ (
    .prog_clk ( { ctsbuf_net_1612143 } ) ,
    .chanx_left_in ( sb_1__1__78_chanx_right_out ) , 
    .chanx_right_in ( sb_1__1__89_chanx_left_out ) , 
    .ccff_head ( sb_1__1__89_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__89_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__89_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__89_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__89_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__89_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__89_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__89_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__89_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__89_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__89_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__89_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__89_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__89_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__89_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__89_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__89_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__89_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__89_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__89_ccff_tail ) ) ;
cbx_1__1_ cbx_9__3_ (
    .prog_clk ( { ctsbuf_net_1852167 } ) ,
    .chanx_left_in ( sb_1__1__79_chanx_right_out ) , 
    .chanx_right_in ( sb_1__1__90_chanx_left_out ) , 
    .ccff_head ( sb_1__1__90_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__90_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__90_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__90_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__90_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__90_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__90_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__90_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__90_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__90_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__90_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__90_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__90_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__90_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__90_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__90_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__90_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__90_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__90_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__90_ccff_tail ) ) ;
cbx_1__1_ cbx_9__4_ (
    .prog_clk ( { ctsbuf_net_2512233 } ) ,
    .chanx_left_in ( sb_1__1__80_chanx_right_out ) , 
    .chanx_right_in ( sb_1__1__91_chanx_left_out ) , 
    .ccff_head ( sb_1__1__91_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__91_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__91_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__91_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__91_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__91_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__91_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__91_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__91_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__91_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__91_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__91_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__91_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__91_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__91_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__91_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__91_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__91_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__91_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__91_ccff_tail ) ) ;
cbx_1__1_ cbx_9__5_ (
    .prog_clk ( { ctsbuf_net_2972279 } ) ,
    .chanx_left_in ( sb_1__1__81_chanx_right_out ) , 
    .chanx_right_in ( sb_1__1__92_chanx_left_out ) , 
    .ccff_head ( sb_1__1__92_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__92_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__92_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__92_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__92_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__92_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__92_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__92_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__92_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__92_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__92_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__92_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__92_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__92_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__92_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__92_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__92_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__92_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__92_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__92_ccff_tail ) ) ;
cbx_1__1_ cbx_9__6_ (
    .prog_clk ( { ctsbuf_net_3452327 } ) ,
    .chanx_left_in ( sb_1__1__82_chanx_right_out ) , 
    .chanx_right_in ( sb_1__1__93_chanx_left_out ) , 
    .ccff_head ( sb_1__1__93_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__93_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__93_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__93_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__93_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__93_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__93_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__93_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__93_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__93_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__93_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__93_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__93_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__93_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__93_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__93_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__93_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__93_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__93_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__93_ccff_tail ) ) ;
cbx_1__1_ cbx_9__7_ (
    .prog_clk ( { ctsbuf_net_3092291 } ) ,
    .chanx_left_in ( sb_1__1__83_chanx_right_out ) , 
    .chanx_right_in ( sb_1__1__94_chanx_left_out ) , 
    .ccff_head ( sb_1__1__94_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__94_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__94_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__94_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__94_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__94_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__94_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__94_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__94_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__94_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__94_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__94_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__94_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__94_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__94_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__94_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__94_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__94_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__94_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__94_ccff_tail ) ) ;
cbx_1__1_ cbx_9__8_ (
    .prog_clk ( { ctsbuf_net_2622244 } ) ,
    .chanx_left_in ( sb_1__1__84_chanx_right_out ) , 
    .chanx_right_in ( sb_1__1__95_chanx_left_out ) , 
    .ccff_head ( sb_1__1__95_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__95_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__95_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__95_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__95_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__95_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__95_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__95_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__95_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__95_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__95_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__95_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__95_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__95_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__95_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__95_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__95_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__95_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__95_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__95_ccff_tail ) ) ;
cbx_1__1_ cbx_9__9_ (
    .prog_clk ( { ctsbuf_net_2162198 } ) ,
    .chanx_left_in ( sb_1__1__85_chanx_right_out ) , 
    .chanx_right_in ( sb_1__1__96_chanx_left_out ) , 
    .ccff_head ( sb_1__1__96_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__96_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__96_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__96_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__96_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__96_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__96_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__96_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__96_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__96_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__96_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__96_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__96_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__96_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__96_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__96_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__96_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__96_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__96_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__96_ccff_tail ) ) ;
cbx_1__1_ cbx_9__10_ (
    .prog_clk ( { ctsbuf_net_1702152 } ) ,
    .chanx_left_in ( sb_1__1__86_chanx_right_out ) , 
    .chanx_right_in ( sb_1__1__97_chanx_left_out ) , 
    .ccff_head ( sb_1__1__97_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__97_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__97_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__97_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__97_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__97_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__97_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__97_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__97_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__97_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__97_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__97_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__97_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__97_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__97_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__97_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__97_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__97_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__97_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__97_ccff_tail ) ) ;
cbx_1__1_ cbx_9__11_ (
    .prog_clk ( { ctsbuf_net_1332115 } ) ,
    .chanx_left_in ( sb_1__1__87_chanx_right_out ) , 
    .chanx_right_in ( sb_1__1__98_chanx_left_out ) , 
    .ccff_head ( sb_1__1__98_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__98_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__98_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__98_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__98_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__98_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__98_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__98_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__98_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__98_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__98_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__98_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__98_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__98_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__98_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__98_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__98_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__98_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__98_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__98_ccff_tail ) ) ;
cbx_1__1_ cbx_10__1_ (
    .prog_clk ( { ctsbuf_net_982080 } ) ,
    .chanx_left_in ( sb_1__1__88_chanx_right_out ) , 
    .chanx_right_in ( sb_1__1__99_chanx_left_out ) , 
    .ccff_head ( sb_1__1__99_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__99_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__99_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__99_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__99_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__99_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__99_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__99_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__99_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__99_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__99_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__99_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__99_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__99_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__99_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__99_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__99_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__99_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__99_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__99_ccff_tail ) ) ;
cbx_1__1_ cbx_10__2_ (
    .prog_clk ( { ctsbuf_net_1272109 } ) ,
    .chanx_left_in ( sb_1__1__89_chanx_right_out ) , 
    .chanx_right_in ( sb_1__1__100_chanx_left_out ) , 
    .ccff_head ( sb_1__1__100_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__100_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__100_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__100_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__100_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__100_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__100_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__100_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__100_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__100_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__100_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__100_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__100_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__100_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__100_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__100_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__100_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__100_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__100_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__100_ccff_tail ) ) ;
cbx_1__1_ cbx_10__3_ (
    .prog_clk ( { ctsbuf_net_1462128 } ) ,
    .chanx_left_in ( sb_1__1__90_chanx_right_out ) , 
    .chanx_right_in ( sb_1__1__101_chanx_left_out ) , 
    .ccff_head ( sb_1__1__101_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__101_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__101_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__101_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__101_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__101_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__101_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__101_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__101_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__101_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__101_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__101_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__101_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__101_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__101_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__101_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__101_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__101_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__101_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__101_ccff_tail ) ) ;
cbx_1__1_ cbx_10__4_ (
    .prog_clk ( { ctsbuf_net_2052187 } ) ,
    .chanx_left_in ( sb_1__1__91_chanx_right_out ) , 
    .chanx_right_in ( sb_1__1__102_chanx_left_out ) , 
    .ccff_head ( sb_1__1__102_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__102_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__102_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__102_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__102_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__102_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__102_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__102_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__102_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__102_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__102_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__102_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__102_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__102_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__102_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__102_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__102_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__102_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__102_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__102_ccff_tail ) ) ;
cbx_1__1_ cbx_10__5_ (
    .prog_clk ( { ctsbuf_net_2532235 } ) ,
    .chanx_left_in ( sb_1__1__92_chanx_right_out ) , 
    .chanx_right_in ( sb_1__1__103_chanx_left_out ) , 
    .ccff_head ( sb_1__1__103_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__103_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__103_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__103_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__103_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__103_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__103_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__103_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__103_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__103_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__103_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__103_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__103_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__103_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__103_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__103_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__103_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__103_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__103_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__103_ccff_tail ) ) ;
cbx_1__1_ cbx_10__6_ (
    .prog_clk ( { ctsbuf_net_2992281 } ) ,
    .chanx_left_in ( sb_1__1__93_chanx_right_out ) , 
    .chanx_right_in ( sb_1__1__104_chanx_left_out ) , 
    .ccff_head ( sb_1__1__104_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__104_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__104_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__104_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__104_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__104_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__104_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__104_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__104_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__104_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__104_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__104_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__104_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__104_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__104_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__104_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__104_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__104_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__104_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__104_ccff_tail ) ) ;
cbx_1__1_ cbx_10__7_ (
    .prog_clk ( { ctsbuf_net_2642246 } ) ,
    .chanx_left_in ( sb_1__1__94_chanx_right_out ) , 
    .chanx_right_in ( sb_1__1__105_chanx_left_out ) , 
    .ccff_head ( sb_1__1__105_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__105_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__105_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__105_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__105_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__105_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__105_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__105_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__105_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__105_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__105_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__105_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__105_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__105_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__105_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__105_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__105_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__105_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__105_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__105_ccff_tail ) ) ;
cbx_1__1_ cbx_10__8_ (
    .prog_clk ( { ctsbuf_net_1922174 } ) ,
    .chanx_left_in ( sb_1__1__95_chanx_right_out ) , 
    .chanx_right_in ( sb_1__1__106_chanx_left_out ) , 
    .ccff_head ( sb_1__1__106_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__106_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__106_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__106_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__106_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__106_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__106_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__106_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__106_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__106_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__106_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__106_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__106_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__106_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__106_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__106_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__106_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__106_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__106_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__106_ccff_tail ) ) ;
cbx_1__1_ cbx_10__9_ (
    .prog_clk ( { p_abuf7 } ) ,
    .chanx_left_in ( sb_1__1__96_chanx_right_out ) , 
    .chanx_right_in ( sb_1__1__107_chanx_left_out ) , 
    .ccff_head ( sb_1__1__107_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__107_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__107_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__107_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__107_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__107_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__107_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__107_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__107_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__107_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__107_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__107_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__107_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__107_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__107_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__107_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__107_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__107_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__107_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__107_ccff_tail ) ) ;
cbx_1__1_ cbx_10__10_ (
    .prog_clk ( { ctsbuf_net_1172099 } ) ,
    .chanx_left_in ( sb_1__1__97_chanx_right_out ) , 
    .chanx_right_in ( sb_1__1__108_chanx_left_out ) , 
    .ccff_head ( sb_1__1__108_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__108_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__108_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__108_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__108_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__108_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__108_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__108_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__108_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__108_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__108_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__108_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__108_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__108_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__108_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__108_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__108_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__108_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__108_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__108_ccff_tail ) ) ;
cbx_1__1_ cbx_10__11_ (
    .prog_clk ( { ctsbuf_net_1032085 } ) ,
    .chanx_left_in ( sb_1__1__98_chanx_right_out ) , 
    .chanx_right_in ( sb_1__1__109_chanx_left_out ) , 
    .ccff_head ( sb_1__1__109_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__109_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__109_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__109_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__109_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__109_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__109_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__109_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__109_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__109_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__109_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__109_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__109_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__109_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__109_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__109_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__109_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__109_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__109_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__109_ccff_tail ) ) ;
cbx_1__1_ cbx_11__1_ (
    .prog_clk ( { ctsbuf_net_732055 } ) ,
    .chanx_left_in ( sb_1__1__99_chanx_right_out ) , 
    .chanx_right_in ( sb_1__1__110_chanx_left_out ) , 
    .ccff_head ( sb_1__1__110_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__110_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__110_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__110_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__110_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__110_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__110_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__110_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__110_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__110_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__110_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__110_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__110_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__110_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__110_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__110_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__110_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__110_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__110_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__110_ccff_tail ) ) ;
cbx_1__1_ cbx_11__2_ (
    .prog_clk ( { ctsbuf_net_1002082 } ) ,
    .chanx_left_in ( sb_1__1__100_chanx_right_out ) , 
    .chanx_right_in ( sb_1__1__111_chanx_left_out ) , 
    .ccff_head ( sb_1__1__111_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__111_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__111_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__111_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__111_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__111_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__111_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__111_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__111_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__111_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__111_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__111_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__111_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__111_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__111_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__111_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__111_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__111_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__111_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__111_ccff_tail ) ) ;
cbx_1__1_ cbx_11__3_ (
    .prog_clk ( { ctsbuf_net_1142096 } ) ,
    .chanx_left_in ( sb_1__1__101_chanx_right_out ) , 
    .chanx_right_in ( sb_1__1__112_chanx_left_out ) , 
    .ccff_head ( sb_1__1__112_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__112_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__112_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__112_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__112_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__112_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__112_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__112_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__112_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__112_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__112_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__112_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__112_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__112_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__112_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__112_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__112_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__112_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__112_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__112_ccff_tail ) ) ;
cbx_1__1_ cbx_11__4_ (
    .prog_clk ( { ctsbuf_net_1642146 } ) ,
    .chanx_left_in ( sb_1__1__102_chanx_right_out ) , 
    .chanx_right_in ( sb_1__1__113_chanx_left_out ) , 
    .ccff_head ( sb_1__1__113_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__113_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__113_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__113_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__113_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__113_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__113_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__113_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__113_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__113_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__113_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__113_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__113_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__113_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__113_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__113_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__113_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__113_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__113_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__113_ccff_tail ) ) ;
cbx_1__1_ cbx_11__5_ (
    .prog_clk ( { ctsbuf_net_2072189 } ) ,
    .chanx_left_in ( sb_1__1__103_chanx_right_out ) , 
    .chanx_right_in ( sb_1__1__114_chanx_left_out ) , 
    .ccff_head ( sb_1__1__114_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__114_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__114_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__114_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__114_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__114_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__114_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__114_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__114_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__114_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__114_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__114_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__114_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__114_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__114_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__114_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__114_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__114_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__114_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__114_ccff_tail ) ) ;
cbx_1__1_ cbx_11__6_ (
    .prog_clk ( { ctsbuf_net_2552237 } ) ,
    .chanx_left_in ( sb_1__1__104_chanx_right_out ) , 
    .chanx_right_in ( sb_1__1__115_chanx_left_out ) , 
    .ccff_head ( sb_1__1__115_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__115_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__115_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__115_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__115_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__115_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__115_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__115_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__115_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__115_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__115_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__115_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__115_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__115_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__115_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__115_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__115_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__115_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__115_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__115_ccff_tail ) ) ;
cbx_1__1_ cbx_11__7_ (
    .prog_clk ( { ctsbuf_net_2192201 } ) ,
    .chanx_left_in ( sb_1__1__105_chanx_right_out ) , 
    .chanx_right_in ( sb_1__1__116_chanx_left_out ) , 
    .ccff_head ( sb_1__1__116_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__116_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__116_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__116_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__116_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__116_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__116_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__116_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__116_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__116_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__116_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__116_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__116_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__116_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__116_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__116_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__116_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__116_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__116_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__116_ccff_tail ) ) ;
cbx_1__1_ cbx_11__8_ (
    .prog_clk ( { ctsbuf_net_1522134 } ) ,
    .chanx_left_in ( sb_1__1__106_chanx_right_out ) , 
    .chanx_right_in ( sb_1__1__117_chanx_left_out ) , 
    .ccff_head ( sb_1__1__117_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__117_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__117_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__117_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__117_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__117_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__117_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__117_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__117_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__117_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__117_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__117_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__117_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__117_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__117_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__117_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__117_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__117_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__117_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__117_ccff_tail ) ) ;
cbx_1__1_ cbx_11__9_ (
    .prog_clk ( { ctsbuf_net_1362118 } ) ,
    .chanx_left_in ( sb_1__1__107_chanx_right_out ) , 
    .chanx_right_in ( sb_1__1__118_chanx_left_out ) , 
    .ccff_head ( sb_1__1__118_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__118_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__118_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__118_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__118_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__118_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__118_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__118_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__118_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__118_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__118_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__118_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__118_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__118_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__118_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__118_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__118_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__118_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__118_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__118_ccff_tail ) ) ;
cbx_1__1_ cbx_11__10_ (
    .prog_clk ( { ctsbuf_net_1052087 } ) ,
    .chanx_left_in ( sb_1__1__108_chanx_right_out ) , 
    .chanx_right_in ( sb_1__1__119_chanx_left_out ) , 
    .ccff_head ( sb_1__1__119_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__119_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__119_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__119_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__119_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__119_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__119_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__119_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__119_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__119_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__119_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__119_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__119_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__119_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__119_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__119_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__119_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__119_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__119_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__119_ccff_tail ) ) ;
cbx_1__1_ cbx_11__11_ (
    .prog_clk ( { ctsbuf_net_772059 } ) ,
    .chanx_left_in ( sb_1__1__109_chanx_right_out ) , 
    .chanx_right_in ( sb_1__1__120_chanx_left_out ) , 
    .ccff_head ( sb_1__1__120_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__120_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__120_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__120_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__120_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__120_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__120_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__120_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__120_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__120_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__120_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__120_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__120_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__120_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__120_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__120_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__120_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__120_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__120_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__120_ccff_tail ) ) ;
cbx_1__1_ cbx_12__1_ (
    .prog_clk ( { ctsbuf_net_572039 } ) ,
    .chanx_left_in ( sb_1__1__110_chanx_right_out ) , 
    .chanx_right_in ( sb_12__1__0_chanx_left_out ) , 
    .ccff_head ( sb_12__1__0_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__121_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__121_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__121_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__121_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__121_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__121_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__121_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__121_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__121_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__121_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__121_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__121_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__121_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__121_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__121_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__121_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__121_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__121_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__121_ccff_tail ) ) ;
cbx_1__1_ cbx_12__2_ (
    .prog_clk ( { ctsbuf_net_652047 } ) ,
    .chanx_left_in ( sb_1__1__111_chanx_right_out ) , 
    .chanx_right_in ( sb_12__1__1_chanx_left_out ) , 
    .ccff_head ( sb_12__1__1_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__122_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__122_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__122_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__122_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__122_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__122_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__122_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__122_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__122_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__122_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__122_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__122_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__122_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__122_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__122_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__122_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__122_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__122_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__122_ccff_tail ) ) ;
cbx_1__1_ cbx_12__3_ (
    .prog_clk ( { ctsbuf_net_862068 } ) ,
    .chanx_left_in ( sb_1__1__112_chanx_right_out ) , 
    .chanx_right_in ( sb_12__1__2_chanx_left_out ) , 
    .ccff_head ( sb_12__1__2_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__123_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__123_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__123_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__123_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__123_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__123_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__123_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__123_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__123_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__123_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__123_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__123_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__123_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__123_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__123_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__123_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__123_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__123_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__123_ccff_tail ) ) ;
cbx_1__1_ cbx_12__4_ (
    .prog_clk ( { ctsbuf_net_1302112 } ) ,
    .chanx_left_in ( sb_1__1__113_chanx_right_out ) , 
    .chanx_right_in ( sb_12__1__3_chanx_left_out ) , 
    .ccff_head ( sb_12__1__3_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__124_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__124_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__124_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__124_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__124_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__124_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__124_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__124_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__124_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__124_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__124_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__124_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__124_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__124_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__124_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__124_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__124_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__124_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__124_ccff_tail ) ) ;
cbx_1__1_ cbx_12__5_ (
    .prog_clk ( { ctsbuf_net_1662148 } ) ,
    .chanx_left_in ( sb_1__1__114_chanx_right_out ) , 
    .chanx_right_in ( sb_12__1__4_chanx_left_out ) , 
    .ccff_head ( sb_12__1__4_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__125_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__125_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__125_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__125_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__125_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__125_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__125_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__125_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__125_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__125_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__125_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__125_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__125_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__125_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__125_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__125_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__125_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__125_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__125_ccff_tail ) ) ;
cbx_1__1_ cbx_12__6_ (
    .prog_clk ( { ctsbuf_net_2092191 } ) ,
    .chanx_left_in ( sb_1__1__115_chanx_right_out ) , 
    .chanx_right_in ( sb_12__1__5_chanx_left_out ) , 
    .ccff_head ( sb_12__1__5_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__126_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__126_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__126_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__126_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__126_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__126_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__126_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__126_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__126_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__126_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__126_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__126_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__126_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__126_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__126_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__126_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__126_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__126_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__126_ccff_tail ) ) ;
cbx_1__1_ cbx_12__7_ (
    .prog_clk ( { ctsbuf_net_1752157 } ) ,
    .chanx_left_in ( sb_1__1__116_chanx_right_out ) , 
    .chanx_right_in ( sb_12__1__6_chanx_left_out ) , 
    .ccff_head ( sb_12__1__6_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__127_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__127_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__127_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__127_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__127_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__127_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__127_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__127_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__127_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__127_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__127_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__127_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__127_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__127_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__127_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__127_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__127_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__127_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__127_ccff_tail ) ) ;
cbx_1__1_ cbx_12__8_ (
    .prog_clk ( { ctsbuf_net_1192101 } ) ,
    .chanx_left_in ( sb_1__1__117_chanx_right_out ) , 
    .chanx_right_in ( sb_12__1__7_chanx_left_out ) , 
    .ccff_head ( sb_12__1__7_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__128_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__128_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__128_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__128_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__128_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__128_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__128_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__128_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__128_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__128_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__128_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__128_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__128_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__128_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__128_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__128_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__128_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__128_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__128_ccff_tail ) ) ;
cbx_1__1_ cbx_12__9_ (
    .prog_clk ( { ctsbuf_net_902072 } ) ,
    .chanx_left_in ( sb_1__1__118_chanx_right_out ) , 
    .chanx_right_in ( sb_12__1__8_chanx_left_out ) , 
    .ccff_head ( sb_12__1__8_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__129_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__129_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__129_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__129_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__129_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__129_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__129_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__129_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__129_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__129_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__129_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__129_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__129_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__129_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__129_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__129_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__129_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__129_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__129_ccff_tail ) ) ;
cbx_1__1_ cbx_12__10_ (
    .prog_clk ( { ctsbuf_net_792061 } ) ,
    .chanx_left_in ( sb_1__1__119_chanx_right_out ) , 
    .chanx_right_in ( sb_12__1__9_chanx_left_out ) , 
    .ccff_head ( sb_12__1__9_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__130_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__130_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__130_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__130_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__130_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__130_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__130_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__130_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__130_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__130_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__130_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__130_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__130_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__130_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__130_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__130_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__130_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__130_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__130_ccff_tail ) ) ;
cbx_1__1_ cbx_12__11_ (
    .prog_clk ( { ctsbuf_net_592041 } ) ,
    .chanx_left_in ( sb_1__1__120_chanx_right_out ) , 
    .chanx_right_in ( sb_12__1__10_chanx_left_out ) , 
    .ccff_head ( sb_12__1__10_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__131_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__131_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__131_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__131_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__131_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__131_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__131_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__131_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__131_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__131_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__131_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__131_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__131_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__131_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__131_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__131_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__131_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__131_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__131_ccff_tail ) ) ;
cbx_1__2_ cbx_1__12_ (
    .prog_clk ( { ctsbuf_net_4162398 } ) ,
    .chanx_left_in ( sb_0__12__0_chanx_right_out ) , 
    .chanx_right_in ( sb_1__12__0_chanx_left_out ) , 
    .ccff_head ( sb_1__12__0_ccff_tail ) , 
    .chanx_left_out ( cbx_1__12__0_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__12__0_chanx_right_out ) , 
    .top_grid_pin_0_ ( cbx_1__12__0_top_grid_pin_0_ ) , 
    .ccff_tail ( cbx_1__12__0_ccff_tail ) ) ;
cbx_1__2_ cbx_2__12_ (
    .prog_clk ( { ctsbuf_net_3292311 } ) ,
    .chanx_left_in ( sb_1__12__0_chanx_right_out ) , 
    .chanx_right_in ( sb_1__12__1_chanx_left_out ) , 
    .ccff_head ( sb_1__12__1_ccff_tail ) , 
    .chanx_left_out ( cbx_1__12__1_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__12__1_chanx_right_out ) , 
    .top_grid_pin_0_ ( cbx_1__12__1_top_grid_pin_0_ ) , 
    .ccff_tail ( cbx_1__12__1_ccff_tail ) ) ;
cbx_1__2_ cbx_3__12_ (
    .prog_clk ( { ctsbuf_net_3292311 } ) ,
    .chanx_left_in ( sb_1__12__1_chanx_right_out ) , 
    .chanx_right_in ( sb_1__12__2_chanx_left_out ) , 
    .ccff_head ( sb_1__12__2_ccff_tail ) , 
    .chanx_left_out ( cbx_1__12__2_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__12__2_chanx_right_out ) , 
    .top_grid_pin_0_ ( cbx_1__12__2_top_grid_pin_0_ ) , 
    .ccff_tail ( cbx_1__12__2_ccff_tail ) ) ;
cbx_1__2_ cbx_4__12_ (
    .prog_clk ( { ctsbuf_net_3002282 } ) ,
    .chanx_left_in ( sb_1__12__2_chanx_right_out ) , 
    .chanx_right_in ( sb_1__12__3_chanx_left_out ) , 
    .ccff_head ( sb_1__12__3_ccff_tail ) , 
    .chanx_left_out ( cbx_1__12__3_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__12__3_chanx_right_out ) , 
    .top_grid_pin_0_ ( cbx_1__12__3_top_grid_pin_0_ ) , 
    .ccff_tail ( cbx_1__12__3_ccff_tail ) ) ;
cbx_1__2_ cbx_5__12_ (
    .prog_clk ( { p_abuf12 } ) ,
    .chanx_left_in ( sb_1__12__3_chanx_right_out ) , 
    .chanx_right_in ( sb_1__12__4_chanx_left_out ) , 
    .ccff_head ( sb_1__12__4_ccff_tail ) , 
    .chanx_left_out ( cbx_1__12__4_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__12__4_chanx_right_out ) , 
    .top_grid_pin_0_ ( cbx_1__12__4_top_grid_pin_0_ ) , 
    .ccff_tail ( cbx_1__12__4_ccff_tail ) ) ;
cbx_1__2_ cbx_6__12_ (
    .prog_clk ( { ctsbuf_net_2102192 } ) ,
    .chanx_left_in ( sb_1__12__4_chanx_right_out ) , 
    .chanx_right_in ( sb_1__12__5_chanx_left_out ) , 
    .ccff_head ( sb_1__12__5_ccff_tail ) , 
    .chanx_left_out ( cbx_1__12__5_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__12__5_chanx_right_out ) , 
    .top_grid_pin_0_ ( cbx_1__12__5_top_grid_pin_0_ ) , 
    .ccff_tail ( cbx_1__12__5_ccff_tail ) ) ;
cbx_1__2_ cbx_7__12_ (
    .prog_clk ( { ctsbuf_net_1532135 } ) ,
    .chanx_left_in ( sb_1__12__5_chanx_right_out ) , 
    .chanx_right_in ( sb_1__12__6_chanx_left_out ) , 
    .ccff_head ( sb_1__12__6_ccff_tail ) , 
    .chanx_left_out ( cbx_1__12__6_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__12__6_chanx_right_out ) , 
    .top_grid_pin_0_ ( cbx_1__12__6_top_grid_pin_0_ ) , 
    .ccff_tail ( cbx_1__12__6_ccff_tail ) ) ;
cbx_1__2_ cbx_8__12_ (
    .prog_clk ( { ctsbuf_net_1312113 } ) ,
    .chanx_left_in ( sb_1__12__6_chanx_right_out ) , 
    .chanx_right_in ( sb_1__12__7_chanx_left_out ) , 
    .ccff_head ( sb_1__12__7_ccff_tail ) , 
    .chanx_left_out ( cbx_1__12__7_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__12__7_chanx_right_out ) , 
    .top_grid_pin_0_ ( cbx_1__12__7_top_grid_pin_0_ ) , 
    .ccff_tail ( cbx_1__12__7_ccff_tail ) ) ;
cbx_1__2_ cbx_9__12_ (
    .prog_clk ( { p_abuf4 } ) ,
    .chanx_left_in ( sb_1__12__7_chanx_right_out ) , 
    .chanx_right_in ( sb_1__12__8_chanx_left_out ) , 
    .ccff_head ( sb_1__12__8_ccff_tail ) , 
    .chanx_left_out ( cbx_1__12__8_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__12__8_chanx_right_out ) , 
    .top_grid_pin_0_ ( cbx_1__12__8_top_grid_pin_0_ ) , 
    .ccff_tail ( cbx_1__12__8_ccff_tail ) ) ;
cbx_1__2_ cbx_10__12_ (
    .prog_clk ( { ctsbuf_net_752057 } ) ,
    .chanx_left_in ( sb_1__12__8_chanx_right_out ) , 
    .chanx_right_in ( sb_1__12__9_chanx_left_out ) , 
    .ccff_head ( sb_1__12__9_ccff_tail ) , 
    .chanx_left_out ( cbx_1__12__9_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__12__9_chanx_right_out ) , 
    .top_grid_pin_0_ ( cbx_1__12__9_top_grid_pin_0_ ) , 
    .ccff_tail ( cbx_1__12__9_ccff_tail ) ) ;
cbx_1__2_ cbx_11__12_ (
    .prog_clk ( { ctsbuf_net_512033 } ) ,
    .chanx_left_in ( sb_1__12__9_chanx_right_out ) , 
    .chanx_right_in ( sb_1__12__10_chanx_left_out ) , 
    .ccff_head ( sb_1__12__10_ccff_tail ) , 
    .chanx_left_out ( cbx_1__12__10_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__12__10_chanx_right_out ) , 
    .top_grid_pin_0_ ( cbx_1__12__10_top_grid_pin_0_ ) , 
    .ccff_tail ( cbx_1__12__10_ccff_tail ) ) ;
cbx_1__2_ cbx_12__12_ (
    .prog_clk ( { ctsbuf_net_462028 } ) ,
    .chanx_left_in ( sb_1__12__10_chanx_right_out ) , 
    .chanx_right_in ( sb_12__12__0_chanx_left_out ) , 
    .ccff_head ( sb_12__12__0_ccff_tail ) , 
    .chanx_left_out ( cbx_1__12__11_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__12__11_chanx_right_out ) , 
    .top_grid_pin_0_ ( cbx_1__12__11_top_grid_pin_0_ ) , 
    .ccff_tail ( cbx_1__12__11_ccff_tail ) ) ;
cby_0__1_ cby_0__1_ (
    .prog_clk ( { ctsbuf_net_4422424 } ) ,
    .chany_bottom_in ( sb_0__0__0_chany_top_out ) , 
    .chany_top_in ( sb_0__1__0_chany_bottom_out ) , 
    .ccff_head ( sb_0__1__0_ccff_tail ) , 
    .chany_bottom_out ( cby_0__1__0_chany_bottom_out ) , 
    .chany_top_out ( cby_0__1__0_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_0__1__0_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_0__1__0_left_grid_pin_0_ ) , 
    .ccff_tail ( cby_0__1__0_ccff_tail ) ) ;
cby_0__1_ cby_0__2_ (
    .prog_clk ( { ctsbuf_net_4942476 } ) ,
    .chany_bottom_in ( sb_0__1__0_chany_top_out ) , 
    .chany_top_in ( sb_0__1__1_chany_bottom_out ) , 
    .ccff_head ( sb_0__1__1_ccff_tail ) , 
    .chany_bottom_out ( cby_0__1__1_chany_bottom_out ) , 
    .chany_top_out ( cby_0__1__1_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_0__1__1_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_0__1__1_left_grid_pin_0_ ) , 
    .ccff_tail ( cby_0__1__1_ccff_tail ) ) ;
cby_0__1_ cby_0__3_ (
    .prog_clk ( { ctsbuf_net_5172499 } ) ,
    .chany_bottom_in ( sb_0__1__1_chany_top_out ) , 
    .chany_top_in ( sb_0__1__2_chany_bottom_out ) , 
    .ccff_head ( sb_0__1__2_ccff_tail ) , 
    .chany_bottom_out ( cby_0__1__2_chany_bottom_out ) , 
    .chany_top_out ( cby_0__1__2_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_0__1__2_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_0__1__2_left_grid_pin_0_ ) , 
    .ccff_tail ( cby_0__1__2_ccff_tail ) ) ;
cby_0__1_ cby_0__4_ (
    .prog_clk ( { ctsbuf_net_5512533 } ) ,
    .chany_bottom_in ( sb_0__1__2_chany_top_out ) , 
    .chany_top_in ( sb_0__1__3_chany_bottom_out ) , 
    .ccff_head ( sb_0__1__3_ccff_tail ) , 
    .chany_bottom_out ( cby_0__1__3_chany_bottom_out ) , 
    .chany_top_out ( cby_0__1__3_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_0__1__3_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_0__1__3_left_grid_pin_0_ ) , 
    .ccff_tail ( cby_0__1__3_ccff_tail ) ) ;
cby_0__1_ cby_0__5_ (
    .prog_clk ( { ctsbuf_net_5692551 } ) ,
    .chany_bottom_in ( sb_0__1__3_chany_top_out ) , 
    .chany_top_in ( sb_0__1__4_chany_bottom_out ) , 
    .ccff_head ( sb_0__1__4_ccff_tail ) , 
    .chany_bottom_out ( cby_0__1__4_chany_bottom_out ) , 
    .chany_top_out ( cby_0__1__4_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_0__1__4_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_0__1__4_left_grid_pin_0_ ) , 
    .ccff_tail ( cby_0__1__4_ccff_tail ) ) ;
cby_0__1_ cby_0__6_ (
    .prog_clk ( { ctsbuf_net_5782560 } ) ,
    .chany_bottom_in ( sb_0__1__4_chany_top_out ) , 
    .chany_top_in ( sb_0__1__5_chany_bottom_out ) , 
    .ccff_head ( sb_0__1__5_ccff_tail ) , 
    .chany_bottom_out ( cby_0__1__5_chany_bottom_out ) , 
    .chany_top_out ( cby_0__1__5_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_0__1__5_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_0__1__5_left_grid_pin_0_ ) , 
    .ccff_tail ( cby_0__1__5_ccff_tail ) ) ;
cby_0__1_ cby_0__7_ (
    .prog_clk ( { ctsbuf_net_5752557 } ) ,
    .chany_bottom_in ( sb_0__1__5_chany_top_out ) , 
    .chany_top_in ( sb_0__1__6_chany_bottom_out ) , 
    .ccff_head ( sb_0__1__6_ccff_tail ) , 
    .chany_bottom_out ( cby_0__1__6_chany_bottom_out ) , 
    .chany_top_out ( cby_0__1__6_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_0__1__6_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_0__1__6_left_grid_pin_0_ ) , 
    .ccff_tail ( cby_0__1__6_ccff_tail ) ) ;
cby_0__1_ cby_0__8_ (
    .prog_clk ( { ctsbuf_net_5642546 } ) ,
    .chany_bottom_in ( sb_0__1__6_chany_top_out ) , 
    .chany_top_in ( sb_0__1__7_chany_bottom_out ) , 
    .ccff_head ( sb_0__1__7_ccff_tail ) , 
    .chany_bottom_out ( cby_0__1__7_chany_bottom_out ) , 
    .chany_top_out ( cby_0__1__7_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_0__1__7_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_0__1__7_left_grid_pin_0_ ) , 
    .ccff_tail ( cby_0__1__7_ccff_tail ) ) ;
cby_0__1_ cby_0__9_ (
    .prog_clk ( { ctsbuf_net_5392521 } ) ,
    .chany_bottom_in ( sb_0__1__7_chany_top_out ) , 
    .chany_top_in ( sb_0__1__8_chany_bottom_out ) , 
    .ccff_head ( sb_0__1__8_ccff_tail ) , 
    .chany_bottom_out ( cby_0__1__8_chany_bottom_out ) , 
    .chany_top_out ( cby_0__1__8_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_0__1__8_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_0__1__8_left_grid_pin_0_ ) , 
    .ccff_tail ( cby_0__1__8_ccff_tail ) ) ;
cby_0__1_ cby_0__10_ (
    .prog_clk ( { ctsbuf_net_5162498 } ) ,
    .chany_bottom_in ( sb_0__1__8_chany_top_out ) , 
    .chany_top_in ( sb_0__1__9_chany_bottom_out ) , 
    .ccff_head ( sb_0__1__9_ccff_tail ) , 
    .chany_bottom_out ( cby_0__1__9_chany_bottom_out ) , 
    .chany_top_out ( cby_0__1__9_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_0__1__9_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_0__1__9_left_grid_pin_0_ ) , 
    .ccff_tail ( cby_0__1__9_ccff_tail ) ) ;
cby_0__1_ cby_0__11_ (
    .prog_clk ( { ctsbuf_net_4752457 } ) ,
    .chany_bottom_in ( sb_0__1__9_chany_top_out ) , 
    .chany_top_in ( sb_0__1__10_chany_bottom_out ) , 
    .ccff_head ( sb_0__1__10_ccff_tail ) , 
    .chany_bottom_out ( cby_0__1__10_chany_bottom_out ) , 
    .chany_top_out ( cby_0__1__10_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_0__1__10_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_0__1__10_left_grid_pin_0_ ) , 
    .ccff_tail ( cby_0__1__10_ccff_tail ) ) ;
cby_0__1_ cby_0__12_ (
    .prog_clk ( { ctsbuf_net_4162398 } ) ,
    .chany_bottom_in ( sb_0__1__10_chany_top_out ) , 
    .chany_top_in ( sb_0__12__0_chany_bottom_out ) , 
    .ccff_head ( sb_0__12__0_ccff_tail ) , 
    .chany_bottom_out ( cby_0__1__11_chany_bottom_out ) , 
    .chany_top_out ( cby_0__1__11_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_0__1__11_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_0__1__11_left_grid_pin_0_ ) , 
    .ccff_tail ( cby_0__1__11_ccff_tail ) ) ;
cby_1__1_ cby_1__1_ (
    .prog_clk ( { ctsbuf_net_4112393 } ) ,
    .chany_bottom_in ( sb_1__0__0_chany_top_out ) , 
    .chany_top_in ( sb_1__1__0_chany_bottom_out ) , 
    .ccff_head ( grid_clb_0_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__0_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__0_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__0_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__0_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__0_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__0_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__0_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__0_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__0_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__0_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__0_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__0_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__0_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__0_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__0_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__0_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__0_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__0_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__0_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__0_ccff_tail ) ) ;
cby_1__1_ cby_1__2_ (
    .prog_clk ( { ctsbuf_net_4602442 } ) ,
    .chany_bottom_in ( sb_1__1__0_chany_top_out ) , 
    .chany_top_in ( sb_1__1__1_chany_bottom_out ) , 
    .ccff_head ( grid_clb_1_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__1_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__1_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__1_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__1_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__1_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__1_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__1_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__1_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__1_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__1_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__1_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__1_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__1_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__1_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__1_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__1_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__1_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__1_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__1_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__1_ccff_tail ) ) ;
cby_1__1_ cby_1__3_ (
    .prog_clk ( { ctsbuf_net_4992481 } ) ,
    .chany_bottom_in ( sb_1__1__1_chany_top_out ) , 
    .chany_top_in ( sb_1__1__2_chany_bottom_out ) , 
    .ccff_head ( grid_clb_2_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__2_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__2_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__2_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__2_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__2_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__2_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__2_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__2_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__2_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__2_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__2_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__2_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__2_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__2_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__2_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__2_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__2_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__2_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__2_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__2_ccff_tail ) ) ;
cby_1__1_ cby_1__4_ (
    .prog_clk ( { ctsbuf_net_5292511 } ) ,
    .chany_bottom_in ( sb_1__1__2_chany_top_out ) , 
    .chany_top_in ( sb_1__1__3_chany_bottom_out ) , 
    .ccff_head ( grid_clb_3_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__3_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__3_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__3_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__3_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__3_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__3_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__3_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__3_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__3_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__3_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__3_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__3_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__3_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__3_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__3_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__3_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__3_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__3_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__3_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__3_ccff_tail ) ) ;
cby_1__1_ cby_1__5_ (
    .prog_clk ( { ctsbuf_net_5542536 } ) ,
    .chany_bottom_in ( sb_1__1__3_chany_top_out ) , 
    .chany_top_in ( sb_1__1__4_chany_bottom_out ) , 
    .ccff_head ( grid_clb_4_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__4_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__4_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__4_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__4_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__4_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__4_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__4_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__4_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__4_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__4_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__4_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__4_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__4_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__4_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__4_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__4_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__4_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__4_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__4_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__4_ccff_tail ) ) ;
cby_1__1_ cby_1__6_ (
    .prog_clk ( { ctsbuf_net_5712553 } ) ,
    .chany_bottom_in ( sb_1__1__4_chany_top_out ) , 
    .chany_top_in ( sb_1__1__5_chany_bottom_out ) , 
    .ccff_head ( grid_clb_5_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__5_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__5_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__5_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__5_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__5_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__5_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__5_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__5_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__5_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__5_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__5_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__5_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__5_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__5_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__5_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__5_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__5_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__5_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__5_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__5_ccff_tail ) ) ;
cby_1__1_ cby_1__7_ (
    .prog_clk ( { ctsbuf_net_5762558 } ) ,
    .chany_bottom_in ( sb_1__1__5_chany_top_out ) , 
    .chany_top_in ( sb_1__1__6_chany_bottom_out ) , 
    .ccff_head ( grid_clb_6_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__6_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__6_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__6_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__6_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__6_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__6_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__6_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__6_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__6_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__6_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__6_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__6_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__6_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__6_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__6_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__6_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__6_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__6_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__6_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__6_ccff_tail ) ) ;
cby_1__1_ cby_1__8_ (
    .prog_clk ( { ctsbuf_net_5612543 } ) ,
    .chany_bottom_in ( sb_1__1__6_chany_top_out ) , 
    .chany_top_in ( sb_1__1__7_chany_bottom_out ) , 
    .ccff_head ( grid_clb_7_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__7_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__7_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__7_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__7_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__7_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__7_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__7_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__7_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__7_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__7_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__7_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__7_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__7_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__7_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__7_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__7_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__7_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__7_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__7_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__7_ccff_tail ) ) ;
cby_1__1_ cby_1__9_ (
    .prog_clk ( { ctsbuf_net_5402522 } ) ,
    .chany_bottom_in ( sb_1__1__7_chany_top_out ) , 
    .chany_top_in ( sb_1__1__8_chany_bottom_out ) , 
    .ccff_head ( grid_clb_8_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__8_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__8_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__8_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__8_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__8_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__8_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__8_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__8_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__8_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__8_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__8_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__8_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__8_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__8_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__8_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__8_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__8_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__8_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__8_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__8_ccff_tail ) ) ;
cby_1__1_ cby_1__10_ (
    .prog_clk ( { ctsbuf_net_5102492 } ) ,
    .chany_bottom_in ( sb_1__1__8_chany_top_out ) , 
    .chany_top_in ( sb_1__1__9_chany_bottom_out ) , 
    .ccff_head ( grid_clb_9_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__9_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__9_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__9_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__9_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__9_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__9_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__9_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__9_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__9_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__9_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__9_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__9_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__9_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__9_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__9_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__9_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__9_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__9_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__9_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__9_ccff_tail ) ) ;
cby_1__1_ cby_1__11_ (
    .prog_clk ( { ctsbuf_net_4762458 } ) ,
    .chany_bottom_in ( sb_1__1__9_chany_top_out ) , 
    .chany_top_in ( sb_1__1__10_chany_bottom_out ) , 
    .ccff_head ( grid_clb_10_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__10_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__10_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__10_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__10_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__10_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__10_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__10_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__10_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__10_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__10_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__10_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__10_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__10_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__10_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__10_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__10_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__10_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__10_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__10_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__10_ccff_tail ) ) ;
cby_1__1_ cby_1__12_ (
    .prog_clk ( { ctsbuf_net_4332415 } ) ,
    .chany_bottom_in ( sb_1__1__10_chany_top_out ) , 
    .chany_top_in ( sb_1__12__0_chany_bottom_out ) , 
    .ccff_head ( grid_clb_11_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__11_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__11_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__11_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__11_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__11_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__11_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__11_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__11_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__11_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__11_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__11_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__11_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__11_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__11_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__11_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__11_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__11_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__11_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__11_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__11_ccff_tail ) ) ;
cby_1__1_ cby_2__1_ (
    .prog_clk ( { ctsbuf_net_3682350 } ) ,
    .chany_bottom_in ( sb_1__0__1_chany_top_out ) , 
    .chany_top_in ( sb_1__1__11_chany_bottom_out ) , 
    .ccff_head ( grid_clb_12_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__12_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__12_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__12_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__12_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__12_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__12_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__12_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__12_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__12_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__12_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__12_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__12_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__12_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__12_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__12_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__12_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__12_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__12_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__12_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__12_ccff_tail ) ) ;
cby_1__1_ cby_2__2_ (
    .prog_clk ( { ctsbuf_net_4182400 } ) ,
    .chany_bottom_in ( sb_1__1__11_chany_top_out ) , 
    .chany_top_in ( sb_1__1__12_chany_bottom_out ) , 
    .ccff_head ( grid_clb_13_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__13_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__13_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__13_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__13_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__13_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__13_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__13_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__13_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__13_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__13_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__13_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__13_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__13_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__13_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__13_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__13_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__13_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__13_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__13_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__13_ccff_tail ) ) ;
cby_1__1_ cby_2__3_ (
    .prog_clk ( { ctsbuf_net_4612443 } ) ,
    .chany_bottom_in ( sb_1__1__12_chany_top_out ) , 
    .chany_top_in ( sb_1__1__13_chany_bottom_out ) , 
    .ccff_head ( grid_clb_14_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__14_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__14_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__14_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__14_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__14_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__14_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__14_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__14_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__14_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__14_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__14_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__14_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__14_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__14_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__14_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__14_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__14_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__14_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__14_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__14_ccff_tail ) ) ;
cby_1__1_ cby_2__4_ (
    .prog_clk ( { ctsbuf_net_5002482 } ) ,
    .chany_bottom_in ( sb_1__1__13_chany_top_out ) , 
    .chany_top_in ( sb_1__1__14_chany_bottom_out ) , 
    .ccff_head ( grid_clb_15_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__15_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__15_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__15_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__15_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__15_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__15_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__15_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__15_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__15_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__15_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__15_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__15_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__15_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__15_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__15_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__15_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__15_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__15_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__15_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__15_ccff_tail ) ) ;
cby_1__1_ cby_2__5_ (
    .prog_clk ( { ctsbuf_net_5302512 } ) ,
    .chany_bottom_in ( sb_1__1__14_chany_top_out ) , 
    .chany_top_in ( sb_1__1__15_chany_bottom_out ) , 
    .ccff_head ( grid_clb_16_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__16_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__16_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__16_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__16_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__16_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__16_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__16_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__16_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__16_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__16_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__16_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__16_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__16_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__16_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__16_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__16_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__16_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__16_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__16_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__16_ccff_tail ) ) ;
cby_1__1_ cby_2__6_ (
    .prog_clk ( { ctsbuf_net_5552537 } ) ,
    .chany_bottom_in ( sb_1__1__15_chany_top_out ) , 
    .chany_top_in ( sb_1__1__16_chany_bottom_out ) , 
    .ccff_head ( grid_clb_17_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__17_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__17_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__17_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__17_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__17_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__17_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__17_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__17_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__17_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__17_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__17_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__17_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__17_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__17_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__17_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__17_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__17_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__17_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__17_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__17_ccff_tail ) ) ;
cby_1__1_ cby_2__7_ (
    .prog_clk ( { ctsbuf_net_5632545 } ) ,
    .chany_bottom_in ( sb_1__1__16_chany_top_out ) , 
    .chany_top_in ( sb_1__1__17_chany_bottom_out ) , 
    .ccff_head ( grid_clb_18_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__18_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__18_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__18_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__18_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__18_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__18_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__18_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__18_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__18_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__18_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__18_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__18_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__18_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__18_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__18_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__18_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__18_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__18_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__18_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__18_ccff_tail ) ) ;
cby_1__1_ cby_2__8_ (
    .prog_clk ( { ctsbuf_net_5412523 } ) ,
    .chany_bottom_in ( sb_1__1__17_chany_top_out ) , 
    .chany_top_in ( sb_1__1__18_chany_bottom_out ) , 
    .ccff_head ( grid_clb_19_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__19_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__19_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__19_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__19_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__19_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__19_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__19_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__19_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__19_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__19_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__19_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__19_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__19_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__19_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__19_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__19_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__19_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__19_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__19_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__19_ccff_tail ) ) ;
cby_1__1_ cby_2__9_ (
    .prog_clk ( { ctsbuf_net_5122494 } ) ,
    .chany_bottom_in ( sb_1__1__18_chany_top_out ) , 
    .chany_top_in ( sb_1__1__19_chany_bottom_out ) , 
    .ccff_head ( grid_clb_20_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__20_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__20_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__20_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__20_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__20_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__20_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__20_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__20_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__20_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__20_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__20_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__20_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__20_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__20_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__20_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__20_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__20_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__20_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__20_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__20_ccff_tail ) ) ;
cby_1__1_ cby_2__10_ (
    .prog_clk ( { ctsbuf_net_4772459 } ) ,
    .chany_bottom_in ( sb_1__1__19_chany_top_out ) , 
    .chany_top_in ( sb_1__1__20_chany_bottom_out ) , 
    .ccff_head ( grid_clb_21_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__21_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__21_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__21_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__21_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__21_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__21_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__21_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__21_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__21_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__21_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__21_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__21_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__21_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__21_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__21_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__21_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__21_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__21_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__21_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__21_ccff_tail ) ) ;
cby_1__1_ cby_2__11_ (
    .prog_clk ( { ctsbuf_net_4352417 } ) ,
    .chany_bottom_in ( sb_1__1__20_chany_top_out ) , 
    .chany_top_in ( sb_1__1__21_chany_bottom_out ) , 
    .ccff_head ( grid_clb_22_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__22_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__22_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__22_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__22_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__22_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__22_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__22_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__22_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__22_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__22_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__22_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__22_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__22_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__22_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__22_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__22_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__22_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__22_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__22_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__22_ccff_tail ) ) ;
cby_1__1_ cby_2__12_ (
    .prog_clk ( { ctsbuf_net_3892371 } ) ,
    .chany_bottom_in ( sb_1__1__21_chany_top_out ) , 
    .chany_top_in ( sb_1__12__1_chany_bottom_out ) , 
    .ccff_head ( grid_clb_23_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__23_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__23_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__23_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__23_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__23_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__23_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__23_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__23_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__23_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__23_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__23_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__23_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__23_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__23_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__23_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__23_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__23_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__23_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__23_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__23_ccff_tail ) ) ;
cby_1__1_ cby_3__1_ (
    .prog_clk ( { ctsbuf_net_3242306 } ) ,
    .chany_bottom_in ( sb_1__0__2_chany_top_out ) , 
    .chany_top_in ( sb_1__1__22_chany_bottom_out ) , 
    .ccff_head ( grid_clb_24_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__24_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__24_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__24_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__24_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__24_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__24_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__24_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__24_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__24_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__24_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__24_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__24_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__24_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__24_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__24_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__24_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__24_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__24_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__24_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__24_ccff_tail ) ) ;
cby_1__1_ cby_3__2_ (
    .prog_clk ( { ctsbuf_net_3742356 } ) ,
    .chany_bottom_in ( sb_1__1__22_chany_top_out ) , 
    .chany_top_in ( sb_1__1__23_chany_bottom_out ) , 
    .ccff_head ( grid_clb_25_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__25_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__25_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__25_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__25_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__25_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__25_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__25_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__25_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__25_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__25_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__25_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__25_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__25_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__25_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__25_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__25_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__25_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__25_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__25_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__25_ccff_tail ) ) ;
cby_1__1_ cby_3__3_ (
    .prog_clk ( { ctsbuf_net_4192401 } ) ,
    .chany_bottom_in ( sb_1__1__23_chany_top_out ) , 
    .chany_top_in ( sb_1__1__24_chany_bottom_out ) , 
    .ccff_head ( grid_clb_26_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__26_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__26_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__26_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__26_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__26_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__26_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__26_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__26_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__26_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__26_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__26_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__26_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__26_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__26_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__26_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__26_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__26_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__26_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__26_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__26_ccff_tail ) ) ;
cby_1__1_ cby_3__4_ (
    .prog_clk ( { ctsbuf_net_4622444 } ) ,
    .chany_bottom_in ( sb_1__1__24_chany_top_out ) , 
    .chany_top_in ( sb_1__1__25_chany_bottom_out ) , 
    .ccff_head ( grid_clb_27_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__27_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__27_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__27_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__27_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__27_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__27_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__27_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__27_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__27_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__27_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__27_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__27_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__27_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__27_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__27_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__27_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__27_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__27_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__27_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__27_ccff_tail ) ) ;
cby_1__1_ cby_3__5_ (
    .prog_clk ( { ctsbuf_net_5012483 } ) ,
    .chany_bottom_in ( sb_1__1__25_chany_top_out ) , 
    .chany_top_in ( sb_1__1__26_chany_bottom_out ) , 
    .ccff_head ( grid_clb_28_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__28_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__28_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__28_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__28_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__28_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__28_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__28_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__28_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__28_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__28_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__28_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__28_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__28_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__28_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__28_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__28_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__28_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__28_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__28_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__28_ccff_tail ) ) ;
cby_1__1_ cby_3__6_ (
    .prog_clk ( { ctsbuf_net_5312513 } ) ,
    .chany_bottom_in ( sb_1__1__26_chany_top_out ) , 
    .chany_top_in ( sb_1__1__27_chany_bottom_out ) , 
    .ccff_head ( grid_clb_29_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__29_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__29_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__29_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__29_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__29_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__29_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__29_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__29_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__29_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__29_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__29_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__29_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__29_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__29_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__29_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__29_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__29_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__29_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__29_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__29_ccff_tail ) ) ;
cby_1__1_ cby_3__7_ (
    .prog_clk ( { ctsbuf_net_5432525 } ) ,
    .chany_bottom_in ( sb_1__1__27_chany_top_out ) , 
    .chany_top_in ( sb_1__1__28_chany_bottom_out ) , 
    .ccff_head ( grid_clb_30_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__30_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__30_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__30_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__30_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__30_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__30_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__30_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__30_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__30_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__30_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__30_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__30_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__30_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__30_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__30_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__30_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__30_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__30_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__30_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__30_ccff_tail ) ) ;
cby_1__1_ cby_3__8_ (
    .prog_clk ( { ctsbuf_net_5132495 } ) ,
    .chany_bottom_in ( sb_1__1__28_chany_top_out ) , 
    .chany_top_in ( sb_1__1__29_chany_bottom_out ) , 
    .ccff_head ( grid_clb_31_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__31_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__31_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__31_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__31_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__31_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__31_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__31_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__31_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__31_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__31_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__31_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__31_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__31_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__31_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__31_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__31_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__31_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__31_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__31_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__31_ccff_tail ) ) ;
cby_1__1_ cby_3__9_ (
    .prog_clk ( { ctsbuf_net_4792461 } ) ,
    .chany_bottom_in ( sb_1__1__29_chany_top_out ) , 
    .chany_top_in ( sb_1__1__30_chany_bottom_out ) , 
    .ccff_head ( grid_clb_32_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__32_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__32_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__32_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__32_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__32_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__32_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__32_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__32_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__32_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__32_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__32_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__32_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__32_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__32_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__32_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__32_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__32_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__32_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__32_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__32_ccff_tail ) ) ;
cby_1__1_ cby_3__10_ (
    .prog_clk ( { ctsbuf_net_4362418 } ) ,
    .chany_bottom_in ( sb_1__1__30_chany_top_out ) , 
    .chany_top_in ( sb_1__1__31_chany_bottom_out ) , 
    .ccff_head ( grid_clb_33_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__33_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__33_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__33_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__33_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__33_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__33_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__33_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__33_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__33_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__33_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__33_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__33_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__33_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__33_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__33_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__33_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__33_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__33_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__33_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__33_ccff_tail ) ) ;
cby_1__1_ cby_3__11_ (
    .prog_clk ( { ctsbuf_net_3912373 } ) ,
    .chany_bottom_in ( sb_1__1__31_chany_top_out ) , 
    .chany_top_in ( sb_1__1__32_chany_bottom_out ) , 
    .ccff_head ( grid_clb_34_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__34_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__34_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__34_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__34_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__34_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__34_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__34_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__34_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__34_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__34_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__34_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__34_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__34_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__34_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__34_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__34_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__34_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__34_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__34_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__34_ccff_tail ) ) ;
cby_1__1_ cby_3__12_ (
    .prog_clk ( { ctsbuf_net_3462328 } ) ,
    .chany_bottom_in ( sb_1__1__32_chany_top_out ) , 
    .chany_top_in ( sb_1__12__2_chany_bottom_out ) , 
    .ccff_head ( grid_clb_35_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__35_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__35_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__35_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__35_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__35_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__35_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__35_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__35_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__35_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__35_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__35_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__35_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__35_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__35_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__35_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__35_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__35_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__35_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__35_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__35_ccff_tail ) ) ;
cby_1__1_ cby_4__1_ (
    .prog_clk ( { ctsbuf_net_2792261 } ) ,
    .chany_bottom_in ( sb_1__0__3_chany_top_out ) , 
    .chany_top_in ( sb_1__1__33_chany_bottom_out ) , 
    .ccff_head ( grid_clb_36_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__36_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__36_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__36_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__36_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__36_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__36_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__36_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__36_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__36_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__36_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__36_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__36_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__36_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__36_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__36_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__36_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__36_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__36_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__36_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__36_ccff_tail ) ) ;
cby_1__1_ cby_4__2_ (
    .prog_clk ( { ctsbuf_net_3312313 } ) ,
    .chany_bottom_in ( sb_1__1__33_chany_top_out ) , 
    .chany_top_in ( sb_1__1__34_chany_bottom_out ) , 
    .ccff_head ( grid_clb_37_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__37_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__37_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__37_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__37_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__37_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__37_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__37_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__37_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__37_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__37_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__37_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__37_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__37_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__37_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__37_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__37_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__37_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__37_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__37_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__37_ccff_tail ) ) ;
cby_1__1_ cby_4__3_ (
    .prog_clk ( { ctsbuf_net_3752357 } ) ,
    .chany_bottom_in ( sb_1__1__34_chany_top_out ) , 
    .chany_top_in ( sb_1__1__35_chany_bottom_out ) , 
    .ccff_head ( grid_clb_38_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__38_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__38_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__38_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__38_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__38_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__38_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__38_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__38_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__38_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__38_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__38_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__38_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__38_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__38_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__38_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__38_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__38_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__38_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__38_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__38_ccff_tail ) ) ;
cby_1__1_ cby_4__4_ (
    .prog_clk ( { ctsbuf_net_4202402 } ) ,
    .chany_bottom_in ( sb_1__1__35_chany_top_out ) , 
    .chany_top_in ( sb_1__1__36_chany_bottom_out ) , 
    .ccff_head ( grid_clb_39_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__39_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__39_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__39_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__39_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__39_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__39_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__39_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__39_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__39_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__39_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__39_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__39_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__39_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__39_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__39_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__39_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__39_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__39_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__39_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__39_ccff_tail ) ) ;
cby_1__1_ cby_4__5_ (
    .prog_clk ( { ctsbuf_net_4632445 } ) ,
    .chany_bottom_in ( sb_1__1__36_chany_top_out ) , 
    .chany_top_in ( sb_1__1__37_chany_bottom_out ) , 
    .ccff_head ( grid_clb_40_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__40_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__40_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__40_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__40_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__40_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__40_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__40_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__40_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__40_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__40_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__40_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__40_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__40_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__40_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__40_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__40_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__40_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__40_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__40_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__40_ccff_tail ) ) ;
cby_1__1_ cby_4__6_ (
    .prog_clk ( { ctsbuf_net_5022484 } ) ,
    .chany_bottom_in ( sb_1__1__37_chany_top_out ) , 
    .chany_top_in ( sb_1__1__38_chany_bottom_out ) , 
    .ccff_head ( grid_clb_41_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__41_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__41_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__41_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__41_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__41_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__41_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__41_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__41_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__41_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__41_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__41_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__41_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__41_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__41_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__41_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__41_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__41_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__41_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__41_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__41_ccff_tail ) ) ;
cby_1__1_ cby_4__7_ (
    .prog_clk ( { ctsbuf_net_5152497 } ) ,
    .chany_bottom_in ( sb_1__1__38_chany_top_out ) , 
    .chany_top_in ( sb_1__1__39_chany_bottom_out ) , 
    .ccff_head ( grid_clb_42_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__42_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__42_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__42_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__42_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__42_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__42_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__42_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__42_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__42_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__42_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__42_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__42_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__42_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__42_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__42_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__42_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__42_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__42_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__42_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__42_ccff_tail ) ) ;
cby_1__1_ cby_4__8_ (
    .prog_clk ( { ctsbuf_net_4802462 } ) ,
    .chany_bottom_in ( sb_1__1__39_chany_top_out ) , 
    .chany_top_in ( sb_1__1__40_chany_bottom_out ) , 
    .ccff_head ( grid_clb_43_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__43_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__43_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__43_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__43_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__43_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__43_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__43_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__43_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__43_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__43_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__43_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__43_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__43_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__43_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__43_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__43_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__43_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__43_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__43_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__43_ccff_tail ) ) ;
cby_1__1_ cby_4__9_ (
    .prog_clk ( { ctsbuf_net_4382420 } ) ,
    .chany_bottom_in ( sb_1__1__40_chany_top_out ) , 
    .chany_top_in ( sb_1__1__41_chany_bottom_out ) , 
    .ccff_head ( grid_clb_44_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__44_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__44_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__44_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__44_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__44_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__44_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__44_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__44_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__44_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__44_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__44_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__44_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__44_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__44_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__44_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__44_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__44_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__44_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__44_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__44_ccff_tail ) ) ;
cby_1__1_ cby_4__10_ (
    .prog_clk ( { ctsbuf_net_3922374 } ) ,
    .chany_bottom_in ( sb_1__1__41_chany_top_out ) , 
    .chany_top_in ( sb_1__1__42_chany_bottom_out ) , 
    .ccff_head ( grid_clb_45_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__45_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__45_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__45_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__45_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__45_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__45_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__45_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__45_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__45_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__45_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__45_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__45_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__45_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__45_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__45_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__45_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__45_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__45_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__45_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__45_ccff_tail ) ) ;
cby_1__1_ cby_4__11_ (
    .prog_clk ( { ctsbuf_net_3482330 } ) ,
    .chany_bottom_in ( sb_1__1__42_chany_top_out ) , 
    .chany_top_in ( sb_1__1__43_chany_bottom_out ) , 
    .ccff_head ( grid_clb_46_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__46_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__46_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__46_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__46_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__46_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__46_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__46_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__46_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__46_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__46_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__46_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__46_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__46_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__46_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__46_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__46_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__46_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__46_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__46_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__46_ccff_tail ) ) ;
cby_1__1_ cby_4__12_ (
    .prog_clk ( { ctsbuf_net_3012283 } ) ,
    .chany_bottom_in ( sb_1__1__43_chany_top_out ) , 
    .chany_top_in ( sb_1__12__3_chany_bottom_out ) , 
    .ccff_head ( grid_clb_47_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__47_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__47_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__47_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__47_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__47_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__47_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__47_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__47_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__47_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__47_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__47_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__47_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__47_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__47_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__47_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__47_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__47_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__47_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__47_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__47_ccff_tail ) ) ;
cby_1__1_ cby_5__1_ (
    .prog_clk ( { ctsbuf_net_2342216 } ) ,
    .chany_bottom_in ( sb_1__0__4_chany_top_out ) , 
    .chany_top_in ( sb_1__1__44_chany_bottom_out ) , 
    .ccff_head ( grid_clb_48_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__48_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__48_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__48_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__48_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__48_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__48_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__48_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__48_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__48_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__48_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__48_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__48_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__48_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__48_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__48_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__48_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__48_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__48_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__48_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__48_ccff_tail ) ) ;
cby_1__1_ cby_5__2_ (
    .prog_clk ( { ctsbuf_net_2852267 } ) ,
    .chany_bottom_in ( sb_1__1__44_chany_top_out ) , 
    .chany_top_in ( sb_1__1__45_chany_bottom_out ) , 
    .ccff_head ( grid_clb_49_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__49_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__49_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__49_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__49_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__49_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__49_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__49_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__49_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__49_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__49_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__49_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__49_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__49_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__49_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__49_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__49_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__49_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__49_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__49_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__49_ccff_tail ) ) ;
cby_1__1_ cby_5__3_ (
    .prog_clk ( { ctsbuf_net_3322314 } ) ,
    .chany_bottom_in ( sb_1__1__45_chany_top_out ) , 
    .chany_top_in ( sb_1__1__46_chany_bottom_out ) , 
    .ccff_head ( grid_clb_50_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__50_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__50_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__50_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__50_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__50_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__50_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__50_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__50_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__50_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__50_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__50_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__50_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__50_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__50_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__50_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__50_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__50_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__50_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__50_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__50_ccff_tail ) ) ;
cby_1__1_ cby_5__4_ (
    .prog_clk ( { ctsbuf_net_3762358 } ) ,
    .chany_bottom_in ( sb_1__1__46_chany_top_out ) , 
    .chany_top_in ( sb_1__1__47_chany_bottom_out ) , 
    .ccff_head ( grid_clb_51_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__51_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__51_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__51_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__51_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__51_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__51_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__51_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__51_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__51_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__51_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__51_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__51_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__51_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__51_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__51_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__51_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__51_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__51_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__51_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__51_ccff_tail ) ) ;
cby_1__1_ cby_5__5_ (
    .prog_clk ( { ctsbuf_net_4212403 } ) ,
    .chany_bottom_in ( sb_1__1__47_chany_top_out ) , 
    .chany_top_in ( sb_1__1__48_chany_bottom_out ) , 
    .ccff_head ( grid_clb_52_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__52_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__52_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__52_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__52_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__52_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__52_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__52_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__52_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__52_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__52_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__52_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__52_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__52_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__52_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__52_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__52_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__52_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__52_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__52_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__52_ccff_tail ) ) ;
cby_1__1_ cby_5__6_ (
    .prog_clk ( { ctsbuf_net_4642446 } ) ,
    .chany_bottom_in ( sb_1__1__48_chany_top_out ) , 
    .chany_top_in ( sb_1__1__49_chany_bottom_out ) , 
    .ccff_head ( grid_clb_53_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__53_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__53_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__53_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__53_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__53_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__53_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__53_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__53_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__53_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__53_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__53_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__53_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__53_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__53_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__53_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__53_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__53_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__53_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__53_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__53_ccff_tail ) ) ;
cby_1__1_ cby_5__7_ (
    .prog_clk ( { ctsbuf_net_4822464 } ) ,
    .chany_bottom_in ( sb_1__1__49_chany_top_out ) , 
    .chany_top_in ( sb_1__1__50_chany_bottom_out ) , 
    .ccff_head ( grid_clb_54_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__54_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__54_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__54_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__54_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__54_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__54_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__54_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__54_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__54_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__54_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__54_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__54_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__54_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__54_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__54_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__54_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__54_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__54_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__54_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__54_ccff_tail ) ) ;
cby_1__1_ cby_5__8_ (
    .prog_clk ( { ctsbuf_net_4392421 } ) ,
    .chany_bottom_in ( sb_1__1__50_chany_top_out ) , 
    .chany_top_in ( sb_1__1__51_chany_bottom_out ) , 
    .ccff_head ( grid_clb_55_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__55_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__55_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__55_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__55_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__55_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__55_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__55_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__55_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__55_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__55_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__55_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__55_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__55_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__55_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__55_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__55_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__55_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__55_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__55_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__55_ccff_tail ) ) ;
cby_1__1_ cby_5__9_ (
    .prog_clk ( { ctsbuf_net_3942376 } ) ,
    .chany_bottom_in ( sb_1__1__51_chany_top_out ) , 
    .chany_top_in ( sb_1__1__52_chany_bottom_out ) , 
    .ccff_head ( grid_clb_56_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__56_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__56_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__56_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__56_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__56_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__56_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__56_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__56_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__56_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__56_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__56_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__56_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__56_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__56_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__56_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__56_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__56_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__56_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__56_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__56_ccff_tail ) ) ;
cby_1__1_ cby_5__10_ (
    .prog_clk ( { ctsbuf_net_3492331 } ) ,
    .chany_bottom_in ( sb_1__1__52_chany_top_out ) , 
    .chany_top_in ( sb_1__1__53_chany_bottom_out ) , 
    .ccff_head ( grid_clb_57_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__57_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__57_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__57_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__57_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__57_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__57_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__57_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__57_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__57_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__57_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__57_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__57_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__57_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__57_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__57_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__57_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__57_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__57_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__57_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__57_ccff_tail ) ) ;
cby_1__1_ cby_5__11_ (
    .prog_clk ( { ctsbuf_net_3032285 } ) ,
    .chany_bottom_in ( sb_1__1__53_chany_top_out ) , 
    .chany_top_in ( sb_1__1__54_chany_bottom_out ) , 
    .ccff_head ( grid_clb_58_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__58_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__58_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__58_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__58_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__58_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__58_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__58_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__58_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__58_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__58_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__58_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__58_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__58_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__58_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__58_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__58_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__58_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__58_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__58_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__58_ccff_tail ) ) ;
cby_1__1_ cby_5__12_ (
    .prog_clk ( { ctsbuf_net_2562238 } ) ,
    .chany_bottom_in ( sb_1__1__54_chany_top_out ) , 
    .chany_top_in ( sb_1__12__4_chany_bottom_out ) , 
    .ccff_head ( grid_clb_59_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__59_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__59_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__59_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__59_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__59_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__59_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__59_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__59_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__59_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__59_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__59_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__59_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__59_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__59_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__59_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__59_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__59_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__59_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__59_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__59_ccff_tail ) ) ;
cby_1__1_ cby_6__1_ (
    .prog_clk ( { ctsbuf_net_1892171 } ) ,
    .chany_bottom_in ( sb_1__0__5_chany_top_out ) , 
    .chany_top_in ( sb_1__1__55_chany_bottom_out ) , 
    .ccff_head ( grid_clb_60_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__60_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__60_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__60_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__60_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__60_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__60_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__60_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__60_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__60_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__60_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__60_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__60_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__60_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__60_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__60_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__60_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__60_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__60_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__60_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__60_ccff_tail ) ) ;
cby_1__1_ cby_6__2_ (
    .prog_clk ( { ctsbuf_net_2412223 } ) ,
    .chany_bottom_in ( sb_1__1__55_chany_top_out ) , 
    .chany_top_in ( sb_1__1__56_chany_bottom_out ) , 
    .ccff_head ( grid_clb_61_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__61_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__61_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__61_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__61_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__61_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__61_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__61_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__61_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__61_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__61_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__61_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__61_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__61_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__61_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__61_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__61_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__61_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__61_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__61_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__61_ccff_tail ) ) ;
cby_1__1_ cby_6__3_ (
    .prog_clk ( { ctsbuf_net_2862268 } ) ,
    .chany_bottom_in ( sb_1__1__56_chany_top_out ) , 
    .chany_top_in ( sb_1__1__57_chany_bottom_out ) , 
    .ccff_head ( grid_clb_62_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__62_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__62_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__62_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__62_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__62_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__62_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__62_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__62_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__62_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__62_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__62_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__62_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__62_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__62_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__62_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__62_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__62_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__62_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__62_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__62_ccff_tail ) ) ;
cby_1__1_ cby_6__4_ (
    .prog_clk ( { ctsbuf_net_3332315 } ) ,
    .chany_bottom_in ( sb_1__1__57_chany_top_out ) , 
    .chany_top_in ( sb_1__1__58_chany_bottom_out ) , 
    .ccff_head ( grid_clb_63_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__63_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__63_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__63_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__63_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__63_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__63_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__63_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__63_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__63_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__63_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__63_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__63_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__63_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__63_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__63_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__63_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__63_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__63_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__63_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__63_ccff_tail ) ) ;
cby_1__1_ cby_6__5_ (
    .prog_clk ( { ctsbuf_net_3772359 } ) ,
    .chany_bottom_in ( sb_1__1__58_chany_top_out ) , 
    .chany_top_in ( sb_1__1__59_chany_bottom_out ) , 
    .ccff_head ( grid_clb_64_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__64_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__64_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__64_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__64_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__64_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__64_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__64_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__64_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__64_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__64_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__64_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__64_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__64_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__64_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__64_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__64_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__64_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__64_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__64_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__64_ccff_tail ) ) ;
cby_1__1_ cby_6__6_ (
    .prog_clk ( { ctsbuf_net_4222404 } ) ,
    .chany_bottom_in ( sb_1__1__59_chany_top_out ) , 
    .chany_top_in ( sb_1__1__60_chany_bottom_out ) , 
    .ccff_head ( grid_clb_65_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__65_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__65_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__65_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__65_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__65_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__65_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__65_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__65_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__65_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__65_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__65_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__65_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__65_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__65_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__65_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__65_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__65_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__65_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__65_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__65_ccff_tail ) ) ;
cby_1__1_ cby_6__7_ (
    .prog_clk ( { p_abuf21 } ) ,
    .chany_bottom_in ( sb_1__1__60_chany_top_out ) , 
    .chany_top_in ( sb_1__1__61_chany_bottom_out ) , 
    .ccff_head ( grid_clb_66_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__66_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__66_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__66_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__66_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__66_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__66_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__66_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__66_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__66_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__66_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__66_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__66_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__66_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__66_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__66_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__66_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__66_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__66_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__66_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__66_ccff_tail ) ) ;
cby_1__1_ cby_6__8_ (
    .prog_clk ( { ctsbuf_net_3952377 } ) ,
    .chany_bottom_in ( sb_1__1__61_chany_top_out ) , 
    .chany_top_in ( sb_1__1__62_chany_bottom_out ) , 
    .ccff_head ( grid_clb_67_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__67_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__67_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__67_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__67_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__67_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__67_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__67_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__67_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__67_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__67_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__67_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__67_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__67_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__67_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__67_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__67_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__67_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__67_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__67_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__67_ccff_tail ) ) ;
cby_1__1_ cby_6__9_ (
    .prog_clk ( { ctsbuf_net_3512333 } ) ,
    .chany_bottom_in ( sb_1__1__62_chany_top_out ) , 
    .chany_top_in ( sb_1__1__63_chany_bottom_out ) , 
    .ccff_head ( grid_clb_68_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__68_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__68_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__68_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__68_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__68_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__68_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__68_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__68_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__68_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__68_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__68_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__68_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__68_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__68_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__68_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__68_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__68_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__68_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__68_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__68_ccff_tail ) ) ;
cby_1__1_ cby_6__10_ (
    .prog_clk ( { ctsbuf_net_3042286 } ) ,
    .chany_bottom_in ( sb_1__1__63_chany_top_out ) , 
    .chany_top_in ( sb_1__1__64_chany_bottom_out ) , 
    .ccff_head ( grid_clb_69_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__69_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__69_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__69_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__69_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__69_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__69_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__69_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__69_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__69_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__69_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__69_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__69_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__69_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__69_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__69_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__69_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__69_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__69_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__69_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__69_ccff_tail ) ) ;
cby_1__1_ cby_6__11_ (
    .prog_clk ( { p_abuf9 } ) ,
    .chany_bottom_in ( sb_1__1__64_chany_top_out ) , 
    .chany_top_in ( sb_1__1__65_chany_bottom_out ) , 
    .ccff_head ( grid_clb_70_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__70_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__70_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__70_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__70_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__70_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__70_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__70_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__70_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__70_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__70_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__70_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__70_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__70_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__70_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__70_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__70_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__70_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__70_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__70_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__70_ccff_tail ) ) ;
cby_1__1_ cby_6__12_ (
    .prog_clk ( { ctsbuf_net_2112193 } ) ,
    .chany_bottom_in ( sb_1__1__65_chany_top_out ) , 
    .chany_top_in ( sb_1__12__5_chany_bottom_out ) , 
    .ccff_head ( grid_clb_71_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__71_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__71_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__71_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__71_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__71_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__71_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__71_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__71_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__71_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__71_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__71_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__71_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__71_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__71_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__71_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__71_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__71_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__71_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__71_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__71_ccff_tail ) ) ;
cby_1__1_ cby_7__1_ (
    .prog_clk ( { ctsbuf_net_1492131 } ) ,
    .chany_bottom_in ( sb_1__0__6_chany_top_out ) , 
    .chany_top_in ( sb_1__1__66_chany_bottom_out ) , 
    .ccff_head ( grid_clb_72_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__72_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__72_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__72_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__72_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__72_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__72_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__72_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__72_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__72_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__72_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__72_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__72_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__72_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__72_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__72_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__72_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__72_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__72_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__72_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__72_ccff_tail ) ) ;
cby_1__1_ cby_7__2_ (
    .prog_clk ( { ctsbuf_net_1952177 } ) ,
    .chany_bottom_in ( sb_1__1__66_chany_top_out ) , 
    .chany_top_in ( sb_1__1__67_chany_bottom_out ) , 
    .ccff_head ( grid_clb_73_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__73_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__73_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__73_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__73_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__73_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__73_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__73_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__73_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__73_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__73_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__73_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__73_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__73_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__73_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__73_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__73_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__73_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__73_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__73_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__73_ccff_tail ) ) ;
cby_1__1_ cby_7__3_ (
    .prog_clk ( { ctsbuf_net_2422224 } ) ,
    .chany_bottom_in ( sb_1__1__67_chany_top_out ) , 
    .chany_top_in ( sb_1__1__68_chany_bottom_out ) , 
    .ccff_head ( grid_clb_74_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__74_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__74_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__74_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__74_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__74_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__74_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__74_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__74_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__74_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__74_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__74_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__74_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__74_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__74_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__74_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__74_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__74_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__74_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__74_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__74_ccff_tail ) ) ;
cby_1__1_ cby_7__4_ (
    .prog_clk ( { ctsbuf_net_2872269 } ) ,
    .chany_bottom_in ( sb_1__1__68_chany_top_out ) , 
    .chany_top_in ( sb_1__1__69_chany_bottom_out ) , 
    .ccff_head ( grid_clb_75_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__75_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__75_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__75_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__75_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__75_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__75_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__75_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__75_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__75_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__75_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__75_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__75_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__75_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__75_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__75_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__75_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__75_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__75_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__75_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__75_ccff_tail ) ) ;
cby_1__1_ cby_7__5_ (
    .prog_clk ( { ctsbuf_net_3342316 } ) ,
    .chany_bottom_in ( sb_1__1__69_chany_top_out ) , 
    .chany_top_in ( sb_1__1__70_chany_bottom_out ) , 
    .ccff_head ( grid_clb_76_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__76_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__76_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__76_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__76_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__76_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__76_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__76_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__76_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__76_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__76_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__76_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__76_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__76_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__76_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__76_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__76_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__76_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__76_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__76_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__76_ccff_tail ) ) ;
cby_1__1_ cby_7__6_ (
    .prog_clk ( { ctsbuf_net_3782360 } ) ,
    .chany_bottom_in ( sb_1__1__70_chany_top_out ) , 
    .chany_top_in ( sb_1__1__71_chany_bottom_out ) , 
    .ccff_head ( grid_clb_77_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__77_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__77_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__77_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__77_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__77_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__77_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__77_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__77_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__77_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__77_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__77_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__77_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__77_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__77_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__77_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__77_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__77_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__77_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__77_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__77_ccff_tail ) ) ;
cby_1__1_ cby_7__7_ (
    .prog_clk ( { ctsbuf_net_3972379 } ) ,
    .chany_bottom_in ( sb_1__1__71_chany_top_out ) , 
    .chany_top_in ( sb_1__1__72_chany_bottom_out ) , 
    .ccff_head ( grid_clb_78_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__78_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__78_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__78_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__78_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__78_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__78_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__78_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__78_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__78_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__78_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__78_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__78_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__78_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__78_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__78_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__78_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__78_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__78_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__78_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__78_ccff_tail ) ) ;
cby_1__1_ cby_7__8_ (
    .prog_clk ( { ctsbuf_net_3522334 } ) ,
    .chany_bottom_in ( sb_1__1__72_chany_top_out ) , 
    .chany_top_in ( sb_1__1__73_chany_bottom_out ) , 
    .ccff_head ( grid_clb_79_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__79_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__79_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__79_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__79_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__79_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__79_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__79_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__79_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__79_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__79_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__79_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__79_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__79_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__79_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__79_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__79_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__79_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__79_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__79_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__79_ccff_tail ) ) ;
cby_1__1_ cby_7__9_ (
    .prog_clk ( { ctsbuf_net_3062288 } ) ,
    .chany_bottom_in ( sb_1__1__73_chany_top_out ) , 
    .chany_top_in ( sb_1__1__74_chany_bottom_out ) , 
    .ccff_head ( grid_clb_80_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__80_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__80_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__80_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__80_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__80_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__80_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__80_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__80_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__80_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__80_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__80_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__80_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__80_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__80_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__80_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__80_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__80_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__80_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__80_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__80_ccff_tail ) ) ;
cby_1__1_ cby_7__10_ (
    .prog_clk ( { ctsbuf_net_2592241 } ) ,
    .chany_bottom_in ( sb_1__1__74_chany_top_out ) , 
    .chany_top_in ( sb_1__1__75_chany_bottom_out ) , 
    .ccff_head ( grid_clb_81_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__81_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__81_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__81_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__81_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__81_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__81_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__81_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__81_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__81_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__81_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__81_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__81_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__81_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__81_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__81_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__81_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__81_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__81_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__81_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__81_ccff_tail ) ) ;
cby_1__1_ cby_7__11_ (
    .prog_clk ( { p_abuf5 } ) ,
    .chany_bottom_in ( sb_1__1__75_chany_top_out ) , 
    .chany_top_in ( sb_1__1__76_chany_bottom_out ) , 
    .ccff_head ( grid_clb_82_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__82_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__82_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__82_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__82_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__82_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__82_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__82_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__82_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__82_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__82_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__82_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__82_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__82_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__82_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__82_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__82_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__82_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__82_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__82_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__82_ccff_tail ) ) ;
cby_1__1_ cby_7__12_ (
    .prog_clk ( { ctsbuf_net_1672149 } ) ,
    .chany_bottom_in ( sb_1__1__76_chany_top_out ) , 
    .chany_top_in ( sb_1__12__6_chany_bottom_out ) , 
    .ccff_head ( grid_clb_83_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__83_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__83_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__83_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__83_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__83_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__83_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__83_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__83_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__83_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__83_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__83_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__83_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__83_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__83_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__83_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__83_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__83_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__83_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__83_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__83_ccff_tail ) ) ;
cby_1__1_ cby_8__1_ (
    .prog_clk ( { ctsbuf_net_1162098 } ) ,
    .chany_bottom_in ( sb_1__0__7_chany_top_out ) , 
    .chany_top_in ( sb_1__1__77_chany_bottom_out ) , 
    .ccff_head ( grid_clb_84_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__84_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__84_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__84_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__84_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__84_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__84_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__84_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__84_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__84_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__84_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__84_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__84_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__84_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__84_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__84_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__84_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__84_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__84_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__84_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__84_ccff_tail ) ) ;
cby_1__1_ cby_8__2_ (
    .prog_clk ( { p_abuf8 } ) ,
    .chany_bottom_in ( sb_1__1__77_chany_top_out ) , 
    .chany_top_in ( sb_1__1__78_chany_bottom_out ) , 
    .ccff_head ( grid_clb_85_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__85_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__85_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__85_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__85_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__85_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__85_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__85_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__85_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__85_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__85_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__85_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__85_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__85_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__85_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__85_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__85_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__85_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__85_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__85_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__85_ccff_tail ) ) ;
cby_1__1_ cby_8__3_ (
    .prog_clk ( { ctsbuf_net_1962178 } ) ,
    .chany_bottom_in ( sb_1__1__78_chany_top_out ) , 
    .chany_top_in ( sb_1__1__79_chany_bottom_out ) , 
    .ccff_head ( grid_clb_86_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__86_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__86_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__86_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__86_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__86_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__86_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__86_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__86_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__86_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__86_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__86_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__86_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__86_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__86_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__86_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__86_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__86_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__86_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__86_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__86_ccff_tail ) ) ;
cby_1__1_ cby_8__4_ (
    .prog_clk ( { ctsbuf_net_2432225 } ) ,
    .chany_bottom_in ( sb_1__1__79_chany_top_out ) , 
    .chany_top_in ( sb_1__1__80_chany_bottom_out ) , 
    .ccff_head ( grid_clb_87_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__87_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__87_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__87_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__87_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__87_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__87_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__87_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__87_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__87_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__87_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__87_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__87_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__87_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__87_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__87_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__87_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__87_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__87_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__87_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__87_ccff_tail ) ) ;
cby_1__1_ cby_8__5_ (
    .prog_clk ( { ctsbuf_net_2882270 } ) ,
    .chany_bottom_in ( sb_1__1__80_chany_top_out ) , 
    .chany_top_in ( sb_1__1__81_chany_bottom_out ) , 
    .ccff_head ( grid_clb_88_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__88_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__88_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__88_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__88_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__88_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__88_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__88_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__88_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__88_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__88_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__88_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__88_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__88_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__88_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__88_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__88_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__88_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__88_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__88_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__88_ccff_tail ) ) ;
cby_1__1_ cby_8__6_ (
    .prog_clk ( { ctsbuf_net_3352317 } ) ,
    .chany_bottom_in ( sb_1__1__81_chany_top_out ) , 
    .chany_top_in ( sb_1__1__82_chany_bottom_out ) , 
    .ccff_head ( grid_clb_89_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__89_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__89_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__89_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__89_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__89_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__89_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__89_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__89_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__89_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__89_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__89_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__89_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__89_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__89_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__89_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__89_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__89_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__89_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__89_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__89_ccff_tail ) ) ;
cby_1__1_ cby_8__7_ (
    .prog_clk ( { ctsbuf_net_3542336 } ) ,
    .chany_bottom_in ( sb_1__1__82_chany_top_out ) , 
    .chany_top_in ( sb_1__1__83_chany_bottom_out ) , 
    .ccff_head ( grid_clb_90_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__90_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__90_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__90_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__90_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__90_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__90_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__90_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__90_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__90_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__90_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__90_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__90_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__90_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__90_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__90_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__90_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__90_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__90_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__90_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__90_ccff_tail ) ) ;
cby_1__1_ cby_8__8_ (
    .prog_clk ( { ctsbuf_net_3082290 } ) ,
    .chany_bottom_in ( sb_1__1__83_chany_top_out ) , 
    .chany_top_in ( sb_1__1__84_chany_bottom_out ) , 
    .ccff_head ( grid_clb_91_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__91_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__91_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__91_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__91_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__91_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__91_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__91_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__91_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__91_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__91_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__91_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__91_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__91_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__91_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__91_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__91_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__91_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__91_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__91_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__91_ccff_tail ) ) ;
cby_1__1_ cby_8__9_ (
    .prog_clk ( { ctsbuf_net_2612243 } ) ,
    .chany_bottom_in ( sb_1__1__84_chany_top_out ) , 
    .chany_top_in ( sb_1__1__85_chany_bottom_out ) , 
    .ccff_head ( grid_clb_92_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__92_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__92_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__92_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__92_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__92_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__92_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__92_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__92_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__92_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__92_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__92_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__92_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__92_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__92_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__92_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__92_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__92_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__92_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__92_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__92_ccff_tail ) ) ;
cby_1__1_ cby_8__10_ (
    .prog_clk ( { ctsbuf_net_2152197 } ) ,
    .chany_bottom_in ( sb_1__1__85_chany_top_out ) , 
    .chany_top_in ( sb_1__1__86_chany_bottom_out ) , 
    .ccff_head ( grid_clb_93_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__93_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__93_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__93_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__93_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__93_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__93_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__93_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__93_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__93_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__93_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__93_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__93_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__93_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__93_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__93_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__93_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__93_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__93_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__93_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__93_ccff_tail ) ) ;
cby_1__1_ cby_8__11_ (
    .prog_clk ( { ctsbuf_net_1692151 } ) ,
    .chany_bottom_in ( sb_1__1__86_chany_top_out ) , 
    .chany_top_in ( sb_1__1__87_chany_bottom_out ) , 
    .ccff_head ( grid_clb_94_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__94_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__94_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__94_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__94_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__94_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__94_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__94_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__94_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__94_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__94_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__94_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__94_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__94_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__94_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__94_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__94_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__94_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__94_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__94_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__94_ccff_tail ) ) ;
cby_1__1_ cby_8__12_ (
    .prog_clk ( { ctsbuf_net_1322114 } ) ,
    .chany_bottom_in ( sb_1__1__87_chany_top_out ) , 
    .chany_top_in ( sb_1__12__7_chany_bottom_out ) , 
    .ccff_head ( grid_clb_95_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__95_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__95_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__95_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__95_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__95_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__95_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__95_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__95_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__95_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__95_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__95_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__95_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__95_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__95_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__95_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__95_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__95_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__95_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__95_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__95_ccff_tail ) ) ;
cby_1__1_ cby_9__1_ (
    .prog_clk ( { ctsbuf_net_942076 } ) ,
    .chany_bottom_in ( sb_1__0__8_chany_top_out ) , 
    .chany_top_in ( sb_1__1__88_chany_bottom_out ) , 
    .ccff_head ( grid_clb_96_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__96_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__96_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__96_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__96_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__96_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__96_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__96_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__96_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__96_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__96_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__96_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__96_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__96_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__96_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__96_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__96_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__96_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__96_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__96_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__96_ccff_tail ) ) ;
cby_1__1_ cby_9__2_ (
    .prog_clk ( { ctsbuf_net_1222104 } ) ,
    .chany_bottom_in ( sb_1__1__88_chany_top_out ) , 
    .chany_top_in ( sb_1__1__89_chany_bottom_out ) , 
    .ccff_head ( grid_clb_97_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__97_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__97_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__97_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__97_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__97_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__97_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__97_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__97_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__97_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__97_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__97_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__97_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__97_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__97_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__97_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__97_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__97_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__97_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__97_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__97_ccff_tail ) ) ;
cby_1__1_ cby_9__3_ (
    .prog_clk ( { ctsbuf_net_1562138 } ) ,
    .chany_bottom_in ( sb_1__1__89_chany_top_out ) , 
    .chany_top_in ( sb_1__1__90_chany_bottom_out ) , 
    .ccff_head ( grid_clb_98_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__98_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__98_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__98_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__98_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__98_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__98_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__98_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__98_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__98_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__98_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__98_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__98_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__98_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__98_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__98_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__98_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__98_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__98_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__98_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__98_ccff_tail ) ) ;
cby_1__1_ cby_9__4_ (
    .prog_clk ( { ctsbuf_net_1972179 } ) ,
    .chany_bottom_in ( sb_1__1__90_chany_top_out ) , 
    .chany_top_in ( sb_1__1__91_chany_bottom_out ) , 
    .ccff_head ( grid_clb_99_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__99_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__99_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__99_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__99_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__99_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__99_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__99_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__99_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__99_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__99_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__99_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__99_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__99_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__99_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__99_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__99_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__99_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__99_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__99_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__99_ccff_tail ) ) ;
cby_1__1_ cby_9__5_ (
    .prog_clk ( { ctsbuf_net_2442226 } ) ,
    .chany_bottom_in ( sb_1__1__91_chany_top_out ) , 
    .chany_top_in ( sb_1__1__92_chany_bottom_out ) , 
    .ccff_head ( grid_clb_100_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__100_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__100_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__100_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__100_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__100_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__100_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__100_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__100_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__100_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__100_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__100_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__100_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__100_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__100_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__100_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__100_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__100_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__100_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__100_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__100_ccff_tail ) ) ;
cby_1__1_ cby_9__6_ (
    .prog_clk ( { ctsbuf_net_2892271 } ) ,
    .chany_bottom_in ( sb_1__1__92_chany_top_out ) , 
    .chany_top_in ( sb_1__1__93_chany_bottom_out ) , 
    .ccff_head ( grid_clb_101_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__101_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__101_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__101_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__101_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__101_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__101_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__101_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__101_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__101_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__101_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__101_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__101_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__101_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__101_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__101_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__101_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__101_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__101_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__101_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__101_ccff_tail ) ) ;
cby_1__1_ cby_9__7_ (
    .prog_clk ( { ctsbuf_net_3102292 } ) ,
    .chany_bottom_in ( sb_1__1__93_chany_top_out ) , 
    .chany_top_in ( sb_1__1__94_chany_bottom_out ) , 
    .ccff_head ( grid_clb_102_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__102_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__102_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__102_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__102_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__102_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__102_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__102_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__102_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__102_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__102_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__102_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__102_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__102_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__102_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__102_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__102_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__102_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__102_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__102_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__102_ccff_tail ) ) ;
cby_1__1_ cby_9__8_ (
    .prog_clk ( { ctsbuf_net_2632245 } ) ,
    .chany_bottom_in ( sb_1__1__94_chany_top_out ) , 
    .chany_top_in ( sb_1__1__95_chany_bottom_out ) , 
    .ccff_head ( grid_clb_103_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__103_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__103_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__103_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__103_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__103_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__103_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__103_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__103_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__103_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__103_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__103_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__103_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__103_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__103_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__103_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__103_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__103_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__103_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__103_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__103_ccff_tail ) ) ;
cby_1__1_ cby_9__9_ (
    .prog_clk ( { ctsbuf_net_2172199 } ) ,
    .chany_bottom_in ( sb_1__1__95_chany_top_out ) , 
    .chany_top_in ( sb_1__1__96_chany_bottom_out ) , 
    .ccff_head ( grid_clb_104_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__104_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__104_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__104_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__104_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__104_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__104_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__104_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__104_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__104_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__104_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__104_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__104_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__104_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__104_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__104_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__104_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__104_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__104_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__104_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__104_ccff_tail ) ) ;
cby_1__1_ cby_9__10_ (
    .prog_clk ( { ctsbuf_net_1712153 } ) ,
    .chany_bottom_in ( sb_1__1__96_chany_top_out ) , 
    .chany_top_in ( sb_1__1__97_chany_bottom_out ) , 
    .ccff_head ( grid_clb_105_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__105_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__105_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__105_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__105_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__105_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__105_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__105_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__105_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__105_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__105_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__105_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__105_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__105_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__105_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__105_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__105_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__105_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__105_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__105_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__105_ccff_tail ) ) ;
cby_1__1_ cby_9__11_ (
    .prog_clk ( { ctsbuf_net_1342116 } ) ,
    .chany_bottom_in ( sb_1__1__97_chany_top_out ) , 
    .chany_top_in ( sb_1__1__98_chany_bottom_out ) , 
    .ccff_head ( grid_clb_106_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__106_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__106_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__106_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__106_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__106_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__106_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__106_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__106_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__106_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__106_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__106_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__106_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__106_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__106_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__106_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__106_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__106_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__106_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__106_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__106_ccff_tail ) ) ;
cby_1__1_ cby_9__12_ (
    .prog_clk ( { ctsbuf_net_1022084 } ) ,
    .chany_bottom_in ( sb_1__1__98_chany_top_out ) , 
    .chany_top_in ( sb_1__12__8_chany_bottom_out ) , 
    .ccff_head ( grid_clb_107_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__107_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__107_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__107_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__107_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__107_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__107_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__107_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__107_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__107_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__107_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__107_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__107_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__107_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__107_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__107_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__107_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__107_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__107_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__107_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__107_ccff_tail ) ) ;
cby_1__1_ cby_10__1_ (
    .prog_clk ( { ctsbuf_net_702052 } ) ,
    .chany_bottom_in ( sb_1__0__9_chany_top_out ) , 
    .chany_top_in ( sb_1__1__99_chany_bottom_out ) , 
    .ccff_head ( grid_clb_108_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__108_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__108_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__108_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__108_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__108_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__108_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__108_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__108_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__108_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__108_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__108_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__108_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__108_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__108_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__108_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__108_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__108_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__108_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__108_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__108_ccff_tail ) ) ;
cby_1__1_ cby_10__2_ (
    .prog_clk ( { ctsbuf_net_952077 } ) ,
    .chany_bottom_in ( sb_1__1__99_chany_top_out ) , 
    .chany_top_in ( sb_1__1__100_chany_bottom_out ) , 
    .ccff_head ( grid_clb_109_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__109_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__109_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__109_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__109_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__109_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__109_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__109_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__109_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__109_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__109_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__109_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__109_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__109_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__109_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__109_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__109_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__109_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__109_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__109_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__109_ccff_tail ) ) ;
cby_1__1_ cby_10__3_ (
    .prog_clk ( { ctsbuf_net_1232105 } ) ,
    .chany_bottom_in ( sb_1__1__100_chany_top_out ) , 
    .chany_top_in ( sb_1__1__101_chany_bottom_out ) , 
    .ccff_head ( grid_clb_110_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__110_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__110_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__110_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__110_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__110_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__110_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__110_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__110_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__110_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__110_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__110_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__110_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__110_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__110_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__110_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__110_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__110_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__110_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__110_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__110_ccff_tail ) ) ;
cby_1__1_ cby_10__4_ (
    .prog_clk ( { ctsbuf_net_1572139 } ) ,
    .chany_bottom_in ( sb_1__1__101_chany_top_out ) , 
    .chany_top_in ( sb_1__1__102_chany_bottom_out ) , 
    .ccff_head ( grid_clb_111_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__111_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__111_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__111_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__111_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__111_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__111_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__111_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__111_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__111_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__111_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__111_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__111_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__111_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__111_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__111_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__111_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__111_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__111_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__111_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__111_ccff_tail ) ) ;
cby_1__1_ cby_10__5_ (
    .prog_clk ( { ctsbuf_net_1982180 } ) ,
    .chany_bottom_in ( sb_1__1__102_chany_top_out ) , 
    .chany_top_in ( sb_1__1__103_chany_bottom_out ) , 
    .ccff_head ( grid_clb_112_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__112_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__112_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__112_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__112_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__112_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__112_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__112_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__112_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__112_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__112_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__112_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__112_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__112_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__112_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__112_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__112_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__112_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__112_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__112_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__112_ccff_tail ) ) ;
cby_1__1_ cby_10__6_ (
    .prog_clk ( { ctsbuf_net_2452227 } ) ,
    .chany_bottom_in ( sb_1__1__103_chany_top_out ) , 
    .chany_top_in ( sb_1__1__104_chany_bottom_out ) , 
    .ccff_head ( grid_clb_113_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__113_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__113_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__113_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__113_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__113_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__113_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__113_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__113_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__113_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__113_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__113_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__113_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__113_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__113_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__113_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__113_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__113_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__113_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__113_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__113_ccff_tail ) ) ;
cby_1__1_ cby_10__7_ (
    .prog_clk ( { ctsbuf_net_2652247 } ) ,
    .chany_bottom_in ( sb_1__1__104_chany_top_out ) , 
    .chany_top_in ( sb_1__1__105_chany_bottom_out ) , 
    .ccff_head ( grid_clb_114_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__114_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__114_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__114_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__114_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__114_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__114_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__114_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__114_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__114_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__114_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__114_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__114_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__114_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__114_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__114_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__114_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__114_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__114_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__114_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__114_ccff_tail ) ) ;
cby_1__1_ cby_10__8_ (
    .prog_clk ( { ctsbuf_net_2182200 } ) ,
    .chany_bottom_in ( sb_1__1__105_chany_top_out ) , 
    .chany_top_in ( sb_1__1__106_chany_bottom_out ) , 
    .ccff_head ( grid_clb_115_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__115_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__115_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__115_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__115_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__115_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__115_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__115_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__115_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__115_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__115_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__115_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__115_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__115_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__115_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__115_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__115_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__115_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__115_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__115_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__115_ccff_tail ) ) ;
cby_1__1_ cby_10__9_ (
    .prog_clk ( { ctsbuf_net_1732155 } ) ,
    .chany_bottom_in ( sb_1__1__106_chany_top_out ) , 
    .chany_top_in ( sb_1__1__107_chany_bottom_out ) , 
    .ccff_head ( grid_clb_116_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__116_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__116_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__116_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__116_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__116_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__116_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__116_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__116_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__116_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__116_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__116_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__116_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__116_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__116_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__116_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__116_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__116_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__116_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__116_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__116_ccff_tail ) ) ;
cby_1__1_ cby_10__10_ (
    .prog_clk ( { ctsbuf_net_1352117 } ) ,
    .chany_bottom_in ( sb_1__1__107_chany_top_out ) , 
    .chany_top_in ( sb_1__1__108_chany_bottom_out ) , 
    .ccff_head ( grid_clb_117_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__117_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__117_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__117_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__117_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__117_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__117_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__117_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__117_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__117_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__117_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__117_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__117_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__117_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__117_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__117_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__117_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__117_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__117_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__117_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__117_ccff_tail ) ) ;
cby_1__1_ cby_10__11_ (
    .prog_clk ( { ctsbuf_net_1042086 } ) ,
    .chany_bottom_in ( sb_1__1__108_chany_top_out ) , 
    .chany_top_in ( sb_1__1__109_chany_bottom_out ) , 
    .ccff_head ( grid_clb_118_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__118_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__118_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__118_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__118_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__118_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__118_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__118_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__118_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__118_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__118_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__118_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__118_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__118_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__118_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__118_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__118_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__118_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__118_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__118_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__118_ccff_tail ) ) ;
cby_1__1_ cby_10__12_ (
    .prog_clk ( { ctsbuf_net_762058 } ) ,
    .chany_bottom_in ( sb_1__1__109_chany_top_out ) , 
    .chany_top_in ( sb_1__12__9_chany_bottom_out ) , 
    .ccff_head ( grid_clb_119_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__119_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__119_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__119_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__119_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__119_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__119_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__119_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__119_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__119_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__119_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__119_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__119_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__119_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__119_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__119_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__119_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__119_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__119_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__119_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__119_ccff_tail ) ) ;
cby_1__1_ cby_11__1_ (
    .prog_clk ( { ctsbuf_net_552037 } ) ,
    .chany_bottom_in ( sb_1__0__10_chany_top_out ) , 
    .chany_top_in ( sb_1__1__110_chany_bottom_out ) , 
    .ccff_head ( grid_clb_120_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__120_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__120_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__120_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__120_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__120_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__120_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__120_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__120_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__120_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__120_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__120_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__120_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__120_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__120_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__120_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__120_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__120_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__120_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__120_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__120_ccff_tail ) ) ;
cby_1__1_ cby_11__2_ (
    .prog_clk ( { ctsbuf_net_712053 } ) ,
    .chany_bottom_in ( sb_1__1__110_chany_top_out ) , 
    .chany_top_in ( sb_1__1__111_chany_bottom_out ) , 
    .ccff_head ( grid_clb_121_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__121_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__121_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__121_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__121_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__121_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__121_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__121_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__121_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__121_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__121_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__121_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__121_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__121_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__121_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__121_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__121_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__121_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__121_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__121_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__121_ccff_tail ) ) ;
cby_1__1_ cby_11__3_ (
    .prog_clk ( { ctsbuf_net_962078 } ) ,
    .chany_bottom_in ( sb_1__1__111_chany_top_out ) , 
    .chany_top_in ( sb_1__1__112_chany_bottom_out ) , 
    .ccff_head ( grid_clb_122_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__122_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__122_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__122_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__122_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__122_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__122_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__122_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__122_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__122_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__122_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__122_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__122_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__122_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__122_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__122_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__122_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__122_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__122_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__122_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__122_ccff_tail ) ) ;
cby_1__1_ cby_11__4_ (
    .prog_clk ( { ctsbuf_net_1242106 } ) ,
    .chany_bottom_in ( sb_1__1__112_chany_top_out ) , 
    .chany_top_in ( sb_1__1__113_chany_bottom_out ) , 
    .ccff_head ( grid_clb_123_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__123_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__123_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__123_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__123_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__123_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__123_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__123_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__123_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__123_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__123_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__123_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__123_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__123_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__123_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__123_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__123_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__123_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__123_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__123_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__123_ccff_tail ) ) ;
cby_1__1_ cby_11__5_ (
    .prog_clk ( { ctsbuf_net_1582140 } ) ,
    .chany_bottom_in ( sb_1__1__113_chany_top_out ) , 
    .chany_top_in ( sb_1__1__114_chany_bottom_out ) , 
    .ccff_head ( grid_clb_124_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__124_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__124_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__124_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__124_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__124_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__124_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__124_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__124_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__124_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__124_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__124_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__124_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__124_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__124_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__124_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__124_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__124_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__124_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__124_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__124_ccff_tail ) ) ;
cby_1__1_ cby_11__6_ (
    .prog_clk ( { ctsbuf_net_1992181 } ) ,
    .chany_bottom_in ( sb_1__1__114_chany_top_out ) , 
    .chany_top_in ( sb_1__1__115_chany_bottom_out ) , 
    .ccff_head ( grid_clb_125_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__125_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__125_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__125_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__125_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__125_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__125_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__125_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__125_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__125_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__125_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__125_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__125_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__125_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__125_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__125_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__125_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__125_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__125_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__125_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__125_ccff_tail ) ) ;
cby_1__1_ cby_11__7_ (
    .prog_clk ( { ctsbuf_net_2202202 } ) ,
    .chany_bottom_in ( sb_1__1__115_chany_top_out ) , 
    .chany_top_in ( sb_1__1__116_chany_bottom_out ) , 
    .ccff_head ( grid_clb_126_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__126_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__126_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__126_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__126_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__126_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__126_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__126_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__126_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__126_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__126_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__126_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__126_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__126_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__126_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__126_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__126_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__126_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__126_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__126_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__126_ccff_tail ) ) ;
cby_1__1_ cby_11__8_ (
    .prog_clk ( { ctsbuf_net_1742156 } ) ,
    .chany_bottom_in ( sb_1__1__116_chany_top_out ) , 
    .chany_top_in ( sb_1__1__117_chany_bottom_out ) , 
    .ccff_head ( grid_clb_127_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__127_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__127_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__127_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__127_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__127_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__127_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__127_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__127_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__127_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__127_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__127_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__127_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__127_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__127_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__127_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__127_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__127_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__127_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__127_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__127_ccff_tail ) ) ;
cby_1__1_ cby_11__9_ (
    .prog_clk ( { ctsbuf_net_1372119 } ) ,
    .chany_bottom_in ( sb_1__1__117_chany_top_out ) , 
    .chany_top_in ( sb_1__1__118_chany_bottom_out ) , 
    .ccff_head ( grid_clb_128_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__128_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__128_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__128_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__128_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__128_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__128_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__128_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__128_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__128_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__128_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__128_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__128_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__128_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__128_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__128_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__128_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__128_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__128_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__128_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__128_ccff_tail ) ) ;
cby_1__1_ cby_11__10_ (
    .prog_clk ( { ctsbuf_net_1062088 } ) ,
    .chany_bottom_in ( sb_1__1__118_chany_top_out ) , 
    .chany_top_in ( sb_1__1__119_chany_bottom_out ) , 
    .ccff_head ( grid_clb_129_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__129_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__129_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__129_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__129_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__129_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__129_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__129_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__129_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__129_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__129_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__129_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__129_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__129_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__129_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__129_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__129_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__129_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__129_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__129_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__129_ccff_tail ) ) ;
cby_1__1_ cby_11__11_ (
    .prog_clk ( { ctsbuf_net_782060 } ) ,
    .chany_bottom_in ( sb_1__1__119_chany_top_out ) , 
    .chany_top_in ( sb_1__1__120_chany_bottom_out ) , 
    .ccff_head ( grid_clb_130_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__130_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__130_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__130_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__130_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__130_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__130_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__130_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__130_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__130_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__130_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__130_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__130_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__130_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__130_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__130_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__130_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__130_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__130_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__130_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__130_ccff_tail ) ) ;
cby_1__1_ cby_11__12_ (
    .prog_clk ( { ctsbuf_net_582040 } ) ,
    .chany_bottom_in ( sb_1__1__120_chany_top_out ) , 
    .chany_top_in ( sb_1__12__10_chany_bottom_out ) , 
    .ccff_head ( grid_clb_131_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__131_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__131_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__131_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__131_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__131_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__131_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__131_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__131_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__131_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__131_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__131_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__131_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__131_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__131_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__131_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__131_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__131_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__131_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__131_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__131_ccff_tail ) ) ;
cby_1__1_ cby_12__1_ (
    .prog_clk ( { ctsbuf_net_452027 } ) ,
    .chany_bottom_in ( sb_12__0__0_chany_top_out ) , 
    .chany_top_in ( sb_12__1__0_chany_bottom_out ) , 
    .ccff_head ( grid_clb_132_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__132_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__132_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__132_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__132_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__132_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__132_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__132_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__132_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__132_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__132_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__132_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__132_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__132_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__132_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__132_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__132_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__132_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__132_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__132_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__132_ccff_tail ) ) ;
cby_1__1_ cby_12__2_ (
    .prog_clk ( { ctsbuf_net_502032 } ) ,
    .chany_bottom_in ( sb_12__1__0_chany_top_out ) , 
    .chany_top_in ( sb_12__1__1_chany_bottom_out ) , 
    .ccff_head ( grid_clb_133_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__133_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__133_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__133_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__133_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__133_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__133_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__133_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__133_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__133_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__133_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__133_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__133_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__133_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__133_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__133_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__133_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__133_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__133_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__133_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__133_ccff_tail ) ) ;
cby_1__1_ cby_12__3_ (
    .prog_clk ( { ctsbuf_net_632045 } ) ,
    .chany_bottom_in ( sb_12__1__1_chany_top_out ) , 
    .chany_top_in ( sb_12__1__2_chany_bottom_out ) , 
    .ccff_head ( grid_clb_134_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__134_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__134_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__134_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__134_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__134_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__134_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__134_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__134_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__134_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__134_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__134_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__134_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__134_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__134_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__134_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__134_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__134_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__134_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__134_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__134_ccff_tail ) ) ;
cby_1__1_ cby_12__4_ (
    .prog_clk ( { ctsbuf_net_832065 } ) ,
    .chany_bottom_in ( sb_12__1__2_chany_top_out ) , 
    .chany_top_in ( sb_12__1__3_chany_bottom_out ) , 
    .ccff_head ( grid_clb_135_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__135_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__135_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__135_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__135_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__135_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__135_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__135_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__135_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__135_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__135_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__135_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__135_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__135_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__135_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__135_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__135_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__135_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__135_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__135_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__135_ccff_tail ) ) ;
cby_1__1_ cby_12__5_ (
    .prog_clk ( { ctsbuf_net_1112093 } ) ,
    .chany_bottom_in ( sb_12__1__3_chany_top_out ) , 
    .chany_top_in ( sb_12__1__4_chany_bottom_out ) , 
    .ccff_head ( grid_clb_136_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__136_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__136_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__136_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__136_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__136_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__136_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__136_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__136_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__136_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__136_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__136_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__136_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__136_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__136_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__136_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__136_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__136_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__136_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__136_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__136_ccff_tail ) ) ;
cby_1__1_ cby_12__6_ (
    .prog_clk ( { ctsbuf_net_1432125 } ) ,
    .chany_bottom_in ( sb_12__1__4_chany_top_out ) , 
    .chany_top_in ( sb_12__1__5_chany_bottom_out ) , 
    .ccff_head ( grid_clb_137_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__137_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__137_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__137_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__137_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__137_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__137_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__137_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__137_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__137_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__137_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__137_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__137_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__137_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__137_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__137_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__137_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__137_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__137_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__137_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__137_ccff_tail ) ) ;
cby_1__1_ cby_12__7_ (
    .prog_clk ( { ctsbuf_net_1762158 } ) ,
    .chany_bottom_in ( sb_12__1__5_chany_top_out ) , 
    .chany_top_in ( sb_12__1__6_chany_bottom_out ) , 
    .ccff_head ( grid_clb_138_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__138_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__138_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__138_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__138_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__138_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__138_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__138_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__138_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__138_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__138_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__138_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__138_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__138_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__138_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__138_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__138_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__138_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__138_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__138_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__138_ccff_tail ) ) ;
cby_1__1_ cby_12__8_ (
    .prog_clk ( { ctsbuf_net_1202102 } ) ,
    .chany_bottom_in ( sb_12__1__6_chany_top_out ) , 
    .chany_top_in ( sb_12__1__7_chany_bottom_out ) , 
    .ccff_head ( grid_clb_139_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__139_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__139_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__139_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__139_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__139_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__139_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__139_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__139_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__139_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__139_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__139_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__139_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__139_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__139_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__139_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__139_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__139_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__139_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__139_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__139_ccff_tail ) ) ;
cby_1__1_ cby_12__9_ (
    .prog_clk ( { ctsbuf_net_912073 } ) ,
    .chany_bottom_in ( sb_12__1__7_chany_top_out ) , 
    .chany_top_in ( sb_12__1__8_chany_bottom_out ) , 
    .ccff_head ( grid_clb_140_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__140_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__140_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__140_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__140_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__140_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__140_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__140_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__140_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__140_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__140_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__140_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__140_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__140_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__140_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__140_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__140_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__140_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__140_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__140_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__140_ccff_tail ) ) ;
cby_1__1_ cby_12__10_ (
    .prog_clk ( { ctsbuf_net_682050 } ) ,
    .chany_bottom_in ( sb_12__1__8_chany_top_out ) , 
    .chany_top_in ( sb_12__1__9_chany_bottom_out ) , 
    .ccff_head ( grid_clb_141_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__141_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__141_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__141_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__141_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__141_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__141_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__141_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__141_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__141_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__141_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__141_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__141_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__141_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__141_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__141_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__141_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__141_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__141_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__141_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__141_ccff_tail ) ) ;
cby_1__1_ cby_12__11_ (
    .prog_clk ( { ctsbuf_net_602042 } ) ,
    .chany_bottom_in ( sb_12__1__9_chany_top_out ) , 
    .chany_top_in ( sb_12__1__10_chany_bottom_out ) , 
    .ccff_head ( grid_clb_142_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__142_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__142_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__142_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__142_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__142_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__142_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__142_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__142_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__142_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__142_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__142_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__142_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__142_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__142_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__142_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__142_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__142_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__142_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__142_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__142_ccff_tail ) ) ;
cby_1__1_ cby_12__12_ (
    .prog_clk ( { ctsbuf_net_462028 } ) ,
    .chany_bottom_in ( sb_12__1__10_chany_top_out ) , 
    .chany_top_in ( sb_12__12__0_chany_bottom_out ) , 
    .ccff_head ( grid_clb_143_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__143_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__143_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__143_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__143_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__143_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__143_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__143_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__143_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__143_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__143_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__143_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__143_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__143_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__143_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__143_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__143_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__143_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__143_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__143_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__143_ccff_tail ) ) ;
direct_interc_0 direct_interc_0_ ( 
    .in ( grid_clb_1_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_0_out ) ) ;
direct_interc_1 direct_interc_1_ ( 
    .in ( grid_clb_2_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_1_out ) ) ;
direct_interc_2 direct_interc_2_ ( 
    .in ( grid_clb_3_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_2_out ) ) ;
direct_interc_3 direct_interc_3_ ( 
    .in ( grid_clb_4_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_3_out ) ) ;
direct_interc_4 direct_interc_4_ ( 
    .in ( grid_clb_5_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_4_out ) ) ;
direct_interc_5 direct_interc_5_ ( 
    .in ( grid_clb_6_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_5_out ) ) ;
direct_interc_6 direct_interc_6_ ( 
    .in ( grid_clb_7_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_6_out ) ) ;
direct_interc_7 direct_interc_7_ ( 
    .in ( grid_clb_8_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_7_out ) ) ;
direct_interc_8 direct_interc_8_ ( 
    .in ( grid_clb_9_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_8_out ) ) ;
direct_interc_9 direct_interc_9_ ( 
    .in ( grid_clb_10_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_9_out ) ) ;
direct_interc_10 direct_interc_10_ ( 
    .in ( grid_clb_11_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_10_out ) ) ;
direct_interc_11 direct_interc_11_ ( 
    .in ( grid_clb_13_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_11_out ) ) ;
direct_interc_12 direct_interc_12_ ( 
    .in ( grid_clb_14_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_12_out ) ) ;
direct_interc_13 direct_interc_13_ ( 
    .in ( grid_clb_15_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_13_out ) ) ;
direct_interc_14 direct_interc_14_ ( 
    .in ( grid_clb_16_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_14_out ) ) ;
direct_interc_15 direct_interc_15_ ( 
    .in ( grid_clb_17_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_15_out ) ) ;
direct_interc_16 direct_interc_16_ ( 
    .in ( grid_clb_18_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_16_out ) ) ;
direct_interc_17 direct_interc_17_ ( 
    .in ( grid_clb_19_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_17_out ) ) ;
direct_interc_18 direct_interc_18_ ( 
    .in ( grid_clb_20_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_18_out ) ) ;
direct_interc_19 direct_interc_19_ ( 
    .in ( grid_clb_21_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_19_out ) ) ;
direct_interc_20 direct_interc_20_ ( 
    .in ( grid_clb_22_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_20_out ) ) ;
direct_interc_21 direct_interc_21_ ( 
    .in ( grid_clb_23_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_21_out ) ) ;
direct_interc_22 direct_interc_22_ ( 
    .in ( grid_clb_25_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_22_out ) ) ;
direct_interc_23 direct_interc_23_ ( 
    .in ( grid_clb_26_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_23_out ) ) ;
direct_interc_24 direct_interc_24_ ( 
    .in ( grid_clb_27_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_24_out ) ) ;
direct_interc_25 direct_interc_25_ ( 
    .in ( grid_clb_28_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_25_out ) ) ;
direct_interc_26 direct_interc_26_ ( 
    .in ( grid_clb_29_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_26_out ) ) ;
direct_interc_27 direct_interc_27_ ( 
    .in ( grid_clb_30_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_27_out ) ) ;
direct_interc_28 direct_interc_28_ ( 
    .in ( grid_clb_31_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_28_out ) ) ;
direct_interc_29 direct_interc_29_ ( 
    .in ( grid_clb_32_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_29_out ) ) ;
direct_interc_30 direct_interc_30_ ( 
    .in ( grid_clb_33_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_30_out ) ) ;
direct_interc_31 direct_interc_31_ ( 
    .in ( grid_clb_34_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_31_out ) ) ;
direct_interc_32 direct_interc_32_ ( 
    .in ( grid_clb_35_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_32_out ) ) ;
direct_interc_33 direct_interc_33_ ( 
    .in ( grid_clb_37_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_33_out ) ) ;
direct_interc_34 direct_interc_34_ ( 
    .in ( grid_clb_38_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_34_out ) ) ;
direct_interc_35 direct_interc_35_ ( 
    .in ( grid_clb_39_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_35_out ) ) ;
direct_interc_36 direct_interc_36_ ( 
    .in ( grid_clb_40_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_36_out ) ) ;
direct_interc_37 direct_interc_37_ ( 
    .in ( grid_clb_41_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_37_out ) ) ;
direct_interc_38 direct_interc_38_ ( 
    .in ( grid_clb_42_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_38_out ) ) ;
direct_interc_39 direct_interc_39_ ( 
    .in ( grid_clb_43_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_39_out ) ) ;
direct_interc_40 direct_interc_40_ ( 
    .in ( grid_clb_44_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_40_out ) ) ;
direct_interc_41 direct_interc_41_ ( 
    .in ( grid_clb_45_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_41_out ) ) ;
direct_interc_42 direct_interc_42_ ( 
    .in ( grid_clb_46_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_42_out ) ) ;
direct_interc_43 direct_interc_43_ ( 
    .in ( grid_clb_47_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_43_out ) ) ;
direct_interc_44 direct_interc_44_ ( 
    .in ( grid_clb_49_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_44_out ) ) ;
direct_interc_45 direct_interc_45_ ( 
    .in ( grid_clb_50_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_45_out ) ) ;
direct_interc_46 direct_interc_46_ ( 
    .in ( grid_clb_51_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_46_out ) ) ;
direct_interc_47 direct_interc_47_ ( 
    .in ( grid_clb_52_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_47_out ) ) ;
direct_interc_48 direct_interc_48_ ( 
    .in ( grid_clb_53_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_48_out ) ) ;
direct_interc_49 direct_interc_49_ ( 
    .in ( grid_clb_54_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_49_out ) ) ;
direct_interc_50 direct_interc_50_ ( 
    .in ( grid_clb_55_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_50_out ) ) ;
direct_interc_51 direct_interc_51_ ( 
    .in ( grid_clb_56_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_51_out ) ) ;
direct_interc_52 direct_interc_52_ ( 
    .in ( grid_clb_57_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_52_out ) ) ;
direct_interc_53 direct_interc_53_ ( 
    .in ( grid_clb_58_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_53_out ) ) ;
direct_interc_54 direct_interc_54_ ( 
    .in ( grid_clb_59_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_54_out ) ) ;
direct_interc_55 direct_interc_55_ ( 
    .in ( grid_clb_61_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_55_out ) ) ;
direct_interc_56 direct_interc_56_ ( 
    .in ( grid_clb_62_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_56_out ) ) ;
direct_interc_57 direct_interc_57_ ( 
    .in ( grid_clb_63_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_57_out ) ) ;
direct_interc_58 direct_interc_58_ ( 
    .in ( grid_clb_64_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_58_out ) ) ;
direct_interc_59 direct_interc_59_ ( 
    .in ( grid_clb_65_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_59_out ) ) ;
direct_interc_60 direct_interc_60_ ( 
    .in ( grid_clb_66_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_60_out ) ) ;
direct_interc_61 direct_interc_61_ ( 
    .in ( grid_clb_67_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_61_out ) ) ;
direct_interc_62 direct_interc_62_ ( 
    .in ( grid_clb_68_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_62_out ) ) ;
direct_interc_63 direct_interc_63_ ( 
    .in ( grid_clb_69_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_63_out ) ) ;
direct_interc_64 direct_interc_64_ ( 
    .in ( grid_clb_70_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_64_out ) ) ;
direct_interc_65 direct_interc_65_ ( 
    .in ( grid_clb_71_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_65_out ) ) ;
direct_interc_66 direct_interc_66_ ( 
    .in ( grid_clb_73_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_66_out ) ) ;
direct_interc_67 direct_interc_67_ ( 
    .in ( grid_clb_74_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_67_out ) ) ;
direct_interc_68 direct_interc_68_ ( 
    .in ( grid_clb_75_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_68_out ) ) ;
direct_interc_69 direct_interc_69_ ( 
    .in ( grid_clb_76_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_69_out ) ) ;
direct_interc_70 direct_interc_70_ ( 
    .in ( grid_clb_77_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_70_out ) ) ;
direct_interc_71 direct_interc_71_ ( 
    .in ( grid_clb_78_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_71_out ) ) ;
direct_interc_72 direct_interc_72_ ( 
    .in ( grid_clb_79_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_72_out ) ) ;
direct_interc_73 direct_interc_73_ ( 
    .in ( grid_clb_80_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_73_out ) ) ;
direct_interc_74 direct_interc_74_ ( 
    .in ( grid_clb_81_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_74_out ) ) ;
direct_interc_75 direct_interc_75_ ( 
    .in ( grid_clb_82_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_75_out ) ) ;
direct_interc_76 direct_interc_76_ ( 
    .in ( grid_clb_83_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_76_out ) ) ;
direct_interc_77 direct_interc_77_ ( 
    .in ( grid_clb_85_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_77_out ) ) ;
direct_interc_78 direct_interc_78_ ( 
    .in ( grid_clb_86_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_78_out ) ) ;
direct_interc_79 direct_interc_79_ ( 
    .in ( grid_clb_87_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_79_out ) ) ;
direct_interc_80 direct_interc_80_ ( 
    .in ( grid_clb_88_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_80_out ) ) ;
direct_interc_81 direct_interc_81_ ( 
    .in ( grid_clb_89_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_81_out ) ) ;
direct_interc_82 direct_interc_82_ ( 
    .in ( grid_clb_90_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_82_out ) ) ;
direct_interc_83 direct_interc_83_ ( 
    .in ( grid_clb_91_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_83_out ) ) ;
direct_interc_84 direct_interc_84_ ( 
    .in ( grid_clb_92_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_84_out ) ) ;
direct_interc_85 direct_interc_85_ ( 
    .in ( grid_clb_93_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_85_out ) ) ;
direct_interc_86 direct_interc_86_ ( 
    .in ( grid_clb_94_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_86_out ) ) ;
direct_interc_87 direct_interc_87_ ( 
    .in ( grid_clb_95_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_87_out ) ) ;
direct_interc_88 direct_interc_88_ ( 
    .in ( grid_clb_97_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_88_out ) ) ;
direct_interc_89 direct_interc_89_ ( 
    .in ( grid_clb_98_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_89_out ) ) ;
direct_interc_90 direct_interc_90_ ( 
    .in ( grid_clb_99_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_90_out ) ) ;
direct_interc_91 direct_interc_91_ ( 
    .in ( grid_clb_100_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_91_out ) ) ;
direct_interc_92 direct_interc_92_ ( 
    .in ( grid_clb_101_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_92_out ) ) ;
direct_interc_93 direct_interc_93_ ( 
    .in ( grid_clb_102_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_93_out ) ) ;
direct_interc_94 direct_interc_94_ ( 
    .in ( grid_clb_103_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_94_out ) ) ;
direct_interc_95 direct_interc_95_ ( 
    .in ( grid_clb_104_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_95_out ) ) ;
direct_interc_96 direct_interc_96_ ( 
    .in ( grid_clb_105_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_96_out ) ) ;
direct_interc_97 direct_interc_97_ ( 
    .in ( grid_clb_106_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_97_out ) ) ;
direct_interc_98 direct_interc_98_ ( 
    .in ( grid_clb_107_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_98_out ) ) ;
direct_interc_99 direct_interc_99_ ( 
    .in ( grid_clb_109_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_99_out ) ) ;
direct_interc_100 direct_interc_100_ ( 
    .in ( grid_clb_110_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_100_out ) ) ;
direct_interc_101 direct_interc_101_ ( 
    .in ( grid_clb_111_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_101_out ) ) ;
direct_interc_102 direct_interc_102_ ( 
    .in ( grid_clb_112_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_102_out ) ) ;
direct_interc_103 direct_interc_103_ ( 
    .in ( grid_clb_113_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_103_out ) ) ;
direct_interc_104 direct_interc_104_ ( 
    .in ( grid_clb_114_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_104_out ) ) ;
direct_interc_105 direct_interc_105_ ( 
    .in ( grid_clb_115_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_105_out ) ) ;
direct_interc_106 direct_interc_106_ ( 
    .in ( grid_clb_116_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_106_out ) ) ;
direct_interc_107 direct_interc_107_ ( 
    .in ( grid_clb_117_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_107_out ) ) ;
direct_interc_108 direct_interc_108_ ( 
    .in ( grid_clb_118_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_108_out ) ) ;
direct_interc_109 direct_interc_109_ ( 
    .in ( grid_clb_119_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_109_out ) ) ;
direct_interc_110 direct_interc_110_ ( 
    .in ( grid_clb_121_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_110_out ) ) ;
direct_interc_111 direct_interc_111_ ( 
    .in ( grid_clb_122_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_111_out ) ) ;
direct_interc_112 direct_interc_112_ ( 
    .in ( grid_clb_123_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_112_out ) ) ;
direct_interc_113 direct_interc_113_ ( 
    .in ( grid_clb_124_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_113_out ) ) ;
direct_interc_114 direct_interc_114_ ( 
    .in ( grid_clb_125_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_114_out ) ) ;
direct_interc_115 direct_interc_115_ ( 
    .in ( grid_clb_126_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_115_out ) ) ;
direct_interc_116 direct_interc_116_ ( 
    .in ( grid_clb_127_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_116_out ) ) ;
direct_interc_117 direct_interc_117_ ( 
    .in ( grid_clb_128_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_117_out ) ) ;
direct_interc_118 direct_interc_118_ ( 
    .in ( grid_clb_129_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_118_out ) ) ;
direct_interc_119 direct_interc_119_ ( 
    .in ( grid_clb_130_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_119_out ) ) ;
direct_interc_120 direct_interc_120_ ( 
    .in ( grid_clb_131_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_120_out ) ) ;
direct_interc_121 direct_interc_121_ ( 
    .in ( grid_clb_133_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_121_out ) ) ;
direct_interc_122 direct_interc_122_ ( 
    .in ( grid_clb_134_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_122_out ) ) ;
direct_interc_123 direct_interc_123_ ( 
    .in ( grid_clb_135_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_123_out ) ) ;
direct_interc_124 direct_interc_124_ ( 
    .in ( grid_clb_136_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_124_out ) ) ;
direct_interc_125 direct_interc_125_ ( 
    .in ( grid_clb_137_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_125_out ) ) ;
direct_interc_126 direct_interc_126_ ( 
    .in ( grid_clb_138_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_126_out ) ) ;
direct_interc_127 direct_interc_127_ ( 
    .in ( grid_clb_139_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_127_out ) ) ;
direct_interc_128 direct_interc_128_ ( 
    .in ( grid_clb_140_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_128_out ) ) ;
direct_interc_129 direct_interc_129_ ( 
    .in ( grid_clb_141_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_129_out ) ) ;
direct_interc_130 direct_interc_130_ ( 
    .in ( grid_clb_142_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_130_out ) ) ;
direct_interc_131 direct_interc_131_ ( 
    .in ( grid_clb_143_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_131_out ) ) ;
direct_interc_132 direct_interc_132_ ( 
    .in ( grid_clb_0_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_132_out ) ) ;
direct_interc_133 direct_interc_133_ ( 
    .in ( grid_clb_12_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_133_out ) ) ;
direct_interc_134 direct_interc_134_ ( 
    .in ( grid_clb_24_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_134_out ) ) ;
direct_interc_135 direct_interc_135_ ( 
    .in ( grid_clb_36_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_135_out ) ) ;
direct_interc_136 direct_interc_136_ ( 
    .in ( grid_clb_48_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_136_out ) ) ;
direct_interc_137 direct_interc_137_ ( 
    .in ( grid_clb_60_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_137_out ) ) ;
direct_interc_138 direct_interc_138_ ( 
    .in ( grid_clb_72_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_138_out ) ) ;
direct_interc_139 direct_interc_139_ ( 
    .in ( grid_clb_84_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_139_out ) ) ;
direct_interc_140 direct_interc_140_ ( 
    .in ( grid_clb_96_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_140_out ) ) ;
direct_interc_141 direct_interc_141_ ( 
    .in ( grid_clb_108_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_141_out ) ) ;
direct_interc_142 direct_interc_142_ ( 
    .in ( grid_clb_120_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_142_out ) ) ;
direct_interc_143 direct_interc_143_ ( 
    .in ( grid_clb_1_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_143_out ) ) ;
direct_interc_144 direct_interc_144_ ( 
    .in ( grid_clb_2_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_144_out ) ) ;
direct_interc_145 direct_interc_145_ ( 
    .in ( grid_clb_3_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_145_out ) ) ;
direct_interc_146 direct_interc_146_ ( 
    .in ( grid_clb_4_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_146_out ) ) ;
direct_interc_147 direct_interc_147_ ( 
    .in ( grid_clb_5_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_147_out ) ) ;
direct_interc_148 direct_interc_148_ ( 
    .in ( grid_clb_6_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_148_out ) ) ;
direct_interc_149 direct_interc_149_ ( 
    .in ( grid_clb_7_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_149_out ) ) ;
direct_interc_150 direct_interc_150_ ( 
    .in ( grid_clb_8_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_150_out ) ) ;
direct_interc_151 direct_interc_151_ ( 
    .in ( grid_clb_9_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_151_out ) ) ;
direct_interc_152 direct_interc_152_ ( 
    .in ( grid_clb_10_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_152_out ) ) ;
direct_interc_153 direct_interc_153_ ( 
    .in ( grid_clb_11_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_153_out ) ) ;
direct_interc_154 direct_interc_154_ ( 
    .in ( grid_clb_13_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_154_out ) ) ;
direct_interc_155 direct_interc_155_ ( 
    .in ( grid_clb_14_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_155_out ) ) ;
direct_interc_156 direct_interc_156_ ( 
    .in ( grid_clb_15_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_156_out ) ) ;
direct_interc_157 direct_interc_157_ ( 
    .in ( grid_clb_16_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_157_out ) ) ;
direct_interc_158 direct_interc_158_ ( 
    .in ( grid_clb_17_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_158_out ) ) ;
direct_interc_159 direct_interc_159_ ( 
    .in ( grid_clb_18_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_159_out ) ) ;
direct_interc_160 direct_interc_160_ ( 
    .in ( grid_clb_19_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_160_out ) ) ;
direct_interc_161 direct_interc_161_ ( 
    .in ( grid_clb_20_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_161_out ) ) ;
direct_interc_162 direct_interc_162_ ( 
    .in ( grid_clb_21_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_162_out ) ) ;
direct_interc_163 direct_interc_163_ ( 
    .in ( grid_clb_22_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_163_out ) ) ;
direct_interc_164 direct_interc_164_ ( 
    .in ( grid_clb_23_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_164_out ) ) ;
direct_interc_165 direct_interc_165_ ( 
    .in ( grid_clb_25_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_165_out ) ) ;
direct_interc_166 direct_interc_166_ ( 
    .in ( grid_clb_26_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_166_out ) ) ;
direct_interc_167 direct_interc_167_ ( 
    .in ( grid_clb_27_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_167_out ) ) ;
direct_interc_168 direct_interc_168_ ( 
    .in ( grid_clb_28_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_168_out ) ) ;
direct_interc_169 direct_interc_169_ ( 
    .in ( grid_clb_29_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_169_out ) ) ;
direct_interc_170 direct_interc_170_ ( 
    .in ( grid_clb_30_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_170_out ) ) ;
direct_interc_171 direct_interc_171_ ( 
    .in ( grid_clb_31_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_171_out ) ) ;
direct_interc_172 direct_interc_172_ ( 
    .in ( grid_clb_32_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_172_out ) ) ;
direct_interc_173 direct_interc_173_ ( 
    .in ( grid_clb_33_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_173_out ) ) ;
direct_interc_174 direct_interc_174_ ( 
    .in ( grid_clb_34_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_174_out ) ) ;
direct_interc_175 direct_interc_175_ ( 
    .in ( grid_clb_35_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_175_out ) ) ;
direct_interc_176 direct_interc_176_ ( 
    .in ( grid_clb_37_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_176_out ) ) ;
direct_interc_177 direct_interc_177_ ( 
    .in ( grid_clb_38_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_177_out ) ) ;
direct_interc_178 direct_interc_178_ ( 
    .in ( grid_clb_39_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_178_out ) ) ;
direct_interc_179 direct_interc_179_ ( 
    .in ( grid_clb_40_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_179_out ) ) ;
direct_interc_180 direct_interc_180_ ( 
    .in ( grid_clb_41_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_180_out ) ) ;
direct_interc_181 direct_interc_181_ ( 
    .in ( grid_clb_42_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_181_out ) ) ;
direct_interc_182 direct_interc_182_ ( 
    .in ( grid_clb_43_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_182_out ) ) ;
direct_interc_183 direct_interc_183_ ( 
    .in ( grid_clb_44_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_183_out ) ) ;
direct_interc_184 direct_interc_184_ ( 
    .in ( grid_clb_45_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_184_out ) ) ;
direct_interc_185 direct_interc_185_ ( 
    .in ( grid_clb_46_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_185_out ) ) ;
direct_interc_186 direct_interc_186_ ( 
    .in ( grid_clb_47_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_186_out ) ) ;
direct_interc_187 direct_interc_187_ ( 
    .in ( grid_clb_49_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_187_out ) ) ;
direct_interc_188 direct_interc_188_ ( 
    .in ( grid_clb_50_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_188_out ) ) ;
direct_interc_189 direct_interc_189_ ( 
    .in ( grid_clb_51_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_189_out ) ) ;
direct_interc_190 direct_interc_190_ ( 
    .in ( grid_clb_52_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_190_out ) ) ;
direct_interc_191 direct_interc_191_ ( 
    .in ( grid_clb_53_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_191_out ) ) ;
direct_interc_192 direct_interc_192_ ( 
    .in ( grid_clb_54_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_192_out ) ) ;
direct_interc_193 direct_interc_193_ ( 
    .in ( grid_clb_55_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_193_out ) ) ;
direct_interc_194 direct_interc_194_ ( 
    .in ( grid_clb_56_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_194_out ) ) ;
direct_interc_195 direct_interc_195_ ( 
    .in ( grid_clb_57_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_195_out ) ) ;
direct_interc_196 direct_interc_196_ ( 
    .in ( grid_clb_58_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_196_out ) ) ;
direct_interc_197 direct_interc_197_ ( 
    .in ( grid_clb_59_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_197_out ) ) ;
direct_interc_198 direct_interc_198_ ( 
    .in ( grid_clb_61_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_198_out ) ) ;
direct_interc_199 direct_interc_199_ ( 
    .in ( grid_clb_62_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_199_out ) ) ;
direct_interc_200 direct_interc_200_ ( 
    .in ( grid_clb_63_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_200_out ) ) ;
direct_interc_201 direct_interc_201_ ( 
    .in ( grid_clb_64_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_201_out ) ) ;
direct_interc_202 direct_interc_202_ ( 
    .in ( grid_clb_65_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_202_out ) ) ;
direct_interc_203 direct_interc_203_ ( 
    .in ( grid_clb_66_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_203_out ) ) ;
direct_interc_204 direct_interc_204_ ( 
    .in ( grid_clb_67_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_204_out ) ) ;
direct_interc_205 direct_interc_205_ ( 
    .in ( grid_clb_68_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_205_out ) ) ;
direct_interc_206 direct_interc_206_ ( 
    .in ( grid_clb_69_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_206_out ) ) ;
direct_interc_207 direct_interc_207_ ( 
    .in ( grid_clb_70_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_207_out ) ) ;
direct_interc_208 direct_interc_208_ ( 
    .in ( grid_clb_71_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_208_out ) ) ;
direct_interc_209 direct_interc_209_ ( 
    .in ( grid_clb_73_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_209_out ) ) ;
direct_interc_210 direct_interc_210_ ( 
    .in ( grid_clb_74_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_210_out ) ) ;
direct_interc_211 direct_interc_211_ ( 
    .in ( grid_clb_75_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_211_out ) ) ;
direct_interc_212 direct_interc_212_ ( 
    .in ( grid_clb_76_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_212_out ) ) ;
direct_interc_213 direct_interc_213_ ( 
    .in ( grid_clb_77_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_213_out ) ) ;
direct_interc_214 direct_interc_214_ ( 
    .in ( grid_clb_78_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_214_out ) ) ;
direct_interc_215 direct_interc_215_ ( 
    .in ( grid_clb_79_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_215_out ) ) ;
direct_interc_216 direct_interc_216_ ( 
    .in ( grid_clb_80_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_216_out ) ) ;
direct_interc_217 direct_interc_217_ ( 
    .in ( grid_clb_81_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_217_out ) ) ;
direct_interc_218 direct_interc_218_ ( 
    .in ( grid_clb_82_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_218_out ) ) ;
direct_interc_219 direct_interc_219_ ( 
    .in ( grid_clb_83_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_219_out ) ) ;
direct_interc_220 direct_interc_220_ ( 
    .in ( grid_clb_85_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_220_out ) ) ;
direct_interc_221 direct_interc_221_ ( 
    .in ( grid_clb_86_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_221_out ) ) ;
direct_interc_222 direct_interc_222_ ( 
    .in ( grid_clb_87_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_222_out ) ) ;
direct_interc_223 direct_interc_223_ ( 
    .in ( grid_clb_88_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_223_out ) ) ;
direct_interc_224 direct_interc_224_ ( 
    .in ( grid_clb_89_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_224_out ) ) ;
direct_interc_225 direct_interc_225_ ( 
    .in ( grid_clb_90_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_225_out ) ) ;
direct_interc_226 direct_interc_226_ ( 
    .in ( grid_clb_91_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_226_out ) ) ;
direct_interc_227 direct_interc_227_ ( 
    .in ( grid_clb_92_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_227_out ) ) ;
direct_interc_228 direct_interc_228_ ( 
    .in ( grid_clb_93_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_228_out ) ) ;
direct_interc_229 direct_interc_229_ ( 
    .in ( grid_clb_94_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_229_out ) ) ;
direct_interc_230 direct_interc_230_ ( 
    .in ( grid_clb_95_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_230_out ) ) ;
direct_interc_231 direct_interc_231_ ( 
    .in ( grid_clb_97_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_231_out ) ) ;
direct_interc_232 direct_interc_232_ ( 
    .in ( grid_clb_98_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_232_out ) ) ;
direct_interc_233 direct_interc_233_ ( 
    .in ( grid_clb_99_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_233_out ) ) ;
direct_interc_234 direct_interc_234_ ( 
    .in ( grid_clb_100_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_234_out ) ) ;
direct_interc_235 direct_interc_235_ ( 
    .in ( grid_clb_101_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_235_out ) ) ;
direct_interc_236 direct_interc_236_ ( 
    .in ( grid_clb_102_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_236_out ) ) ;
direct_interc_237 direct_interc_237_ ( 
    .in ( grid_clb_103_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_237_out ) ) ;
direct_interc_238 direct_interc_238_ ( 
    .in ( grid_clb_104_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_238_out ) ) ;
direct_interc_239 direct_interc_239_ ( 
    .in ( grid_clb_105_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_239_out ) ) ;
direct_interc_240 direct_interc_240_ ( 
    .in ( grid_clb_106_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_240_out ) ) ;
direct_interc_241 direct_interc_241_ ( 
    .in ( grid_clb_107_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_241_out ) ) ;
direct_interc_242 direct_interc_242_ ( 
    .in ( grid_clb_109_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_242_out ) ) ;
direct_interc_243 direct_interc_243_ ( 
    .in ( grid_clb_110_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_243_out ) ) ;
direct_interc_244 direct_interc_244_ ( 
    .in ( grid_clb_111_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_244_out ) ) ;
direct_interc_245 direct_interc_245_ ( 
    .in ( grid_clb_112_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_245_out ) ) ;
direct_interc_246 direct_interc_246_ ( 
    .in ( grid_clb_113_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_246_out ) ) ;
direct_interc_247 direct_interc_247_ ( 
    .in ( grid_clb_114_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_247_out ) ) ;
direct_interc_248 direct_interc_248_ ( 
    .in ( grid_clb_115_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_248_out ) ) ;
direct_interc_249 direct_interc_249_ ( 
    .in ( grid_clb_116_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_249_out ) ) ;
direct_interc_250 direct_interc_250_ ( 
    .in ( grid_clb_117_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_250_out ) ) ;
direct_interc_251 direct_interc_251_ ( 
    .in ( grid_clb_118_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_251_out ) ) ;
direct_interc_252 direct_interc_252_ ( 
    .in ( grid_clb_119_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_252_out ) ) ;
direct_interc_253 direct_interc_253_ ( 
    .in ( grid_clb_121_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_253_out ) ) ;
direct_interc_254 direct_interc_254_ ( 
    .in ( grid_clb_122_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_254_out ) ) ;
direct_interc_255 direct_interc_255_ ( 
    .in ( grid_clb_123_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_255_out ) ) ;
direct_interc_256 direct_interc_256_ ( 
    .in ( grid_clb_124_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_256_out ) ) ;
direct_interc_257 direct_interc_257_ ( 
    .in ( grid_clb_125_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_257_out ) ) ;
direct_interc_258 direct_interc_258_ ( 
    .in ( grid_clb_126_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_258_out ) ) ;
direct_interc_259 direct_interc_259_ ( 
    .in ( grid_clb_127_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_259_out ) ) ;
direct_interc_260 direct_interc_260_ ( 
    .in ( grid_clb_128_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_260_out ) ) ;
direct_interc_261 direct_interc_261_ ( 
    .in ( grid_clb_129_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_261_out ) ) ;
direct_interc_262 direct_interc_262_ ( 
    .in ( grid_clb_130_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_262_out ) ) ;
direct_interc_263 direct_interc_263_ ( 
    .in ( grid_clb_131_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_263_out ) ) ;
direct_interc_264 direct_interc_264_ ( 
    .in ( grid_clb_133_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_264_out ) ) ;
direct_interc_265 direct_interc_265_ ( 
    .in ( grid_clb_134_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_265_out ) ) ;
direct_interc_266 direct_interc_266_ ( 
    .in ( grid_clb_135_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_266_out ) ) ;
direct_interc_267 direct_interc_267_ ( 
    .in ( grid_clb_136_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_267_out ) ) ;
direct_interc_268 direct_interc_268_ ( 
    .in ( grid_clb_137_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_268_out ) ) ;
direct_interc_269 direct_interc_269_ ( 
    .in ( grid_clb_138_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_269_out ) ) ;
direct_interc_270 direct_interc_270_ ( 
    .in ( grid_clb_139_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_270_out ) ) ;
direct_interc_271 direct_interc_271_ ( 
    .in ( grid_clb_140_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_271_out ) ) ;
direct_interc_272 direct_interc_272_ ( 
    .in ( grid_clb_141_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_272_out ) ) ;
direct_interc_273 direct_interc_273_ ( 
    .in ( grid_clb_142_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_273_out ) ) ;
direct_interc_274 direct_interc_274_ ( 
    .in ( grid_clb_143_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_274_out ) ) ;
direct_interc_275 direct_interc_275_ ( 
    .in ( grid_clb_0_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_275_out ) ) ;
direct_interc_276 direct_interc_276_ ( 
    .in ( grid_clb_12_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_276_out ) ) ;
direct_interc_277 direct_interc_277_ ( 
    .in ( grid_clb_24_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_277_out ) ) ;
direct_interc_278 direct_interc_278_ ( 
    .in ( grid_clb_36_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_278_out ) ) ;
direct_interc_279 direct_interc_279_ ( 
    .in ( grid_clb_48_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_279_out ) ) ;
direct_interc_280 direct_interc_280_ ( 
    .in ( grid_clb_60_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_280_out ) ) ;
direct_interc_281 direct_interc_281_ ( 
    .in ( grid_clb_72_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_281_out ) ) ;
direct_interc_282 direct_interc_282_ ( 
    .in ( grid_clb_84_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_282_out ) ) ;
direct_interc_283 direct_interc_283_ ( 
    .in ( grid_clb_96_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_283_out ) ) ;
direct_interc_284 direct_interc_284_ ( 
    .in ( grid_clb_108_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_284_out ) ) ;
direct_interc_285 direct_interc_285_ ( 
    .in ( grid_clb_120_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_285_out ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_440 ( .A ( BUF_net_1175 ) , 
    .X ( BUF_net_440 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_441 ( .A ( BUF_net_842 ) , 
    .X ( BUF_net_441 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_442 ( .A ( BUF_net_713 ) , 
    .X ( BUF_net_442 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_443 ( .A ( BUF_net_841 ) , 
    .X ( BUF_net_443 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_444 ( .A ( BUF_net_711 ) , 
    .X ( BUF_net_444 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_445 ( .A ( BUF_net_844 ) , 
    .X ( BUF_net_445 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_446 ( .A ( BUF_net_960 ) , 
    .X ( BUF_net_446 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_447 ( .A ( BUF_net_843 ) , 
    .X ( BUF_net_447 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_448 ( .A ( BUF_net_1092 ) , 
    .X ( BUF_net_448 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_449 ( .A ( BUF_net_708 ) , 
    .X ( BUF_net_449 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_450 ( .A ( BUF_net_956 ) , 
    .X ( BUF_net_450 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_451 ( .A ( BUF_net_836 ) , 
    .X ( BUF_net_451 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_452 ( .A ( BUF_net_1175 ) , 
    .X ( BUF_net_452 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_846 ( .A ( BUF_net_1253 ) , 
    .X ( BUF_net_846 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_847 ( .A ( BUF_net_1076 ) , 
    .X ( BUF_net_847 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_718 ( .A ( BUF_net_913 ) , 
    .X ( BUF_net_718 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_719 ( .A ( BUF_net_962 ) , 
    .X ( BUF_net_719 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_720 ( .A ( BUF_net_914 ) , 
    .X ( BUF_net_720 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_458 ( .A ( BUF_net_960 ) , 
    .X ( BUF_net_458 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_848 ( .A ( BUF_net_1092 ) , 
    .X ( BUF_net_848 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_849 ( .A ( BUF_net_1034 ) , 
    .X ( BUF_net_849 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_850 ( .A ( BUF_net_1078 ) , 
    .X ( BUF_net_850 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_851 ( .A ( BUF_net_1037 ) , 
    .X ( BUF_net_851 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_463 ( .A ( BUF_net_836 ) , 
    .X ( BUF_net_463 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_464 ( .A ( Test_en[0] ) , 
    .X ( BUF_net_464 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_852 ( .A ( BUF_net_1573 ) , 
    .X ( BUF_net_852 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_726 ( .A ( BUF_net_915 ) , 
    .X ( BUF_net_726 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_727 ( .A ( BUF_net_965 ) , 
    .X ( BUF_net_727 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_853 ( .A ( BUF_net_1035 ) , 
    .X ( BUF_net_853 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_854 ( .A ( BUF_net_1385 ) , 
    .X ( BUF_net_854 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_470 ( .A ( BUF_net_831 ) , 
    .X ( BUF_net_470 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_730 ( .A ( BUF_net_916 ) , 
    .X ( BUF_net_730 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_731 ( .A ( BUF_net_963 ) , 
    .X ( BUF_net_731 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_966 ( .A ( BUF_net_1253 ) , 
    .X ( BUF_net_966 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_967 ( .A ( BUF_net_1177 ) , 
    .X ( BUF_net_967 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_475 ( .A ( BUF_net_955 ) , 
    .X ( BUF_net_475 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_476 ( .A ( Test_en[0] ) , 
    .X ( BUF_net_476 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_857 ( .A ( BUF_net_1083 ) , 
    .X ( BUF_net_857 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_858 ( .A ( BUF_net_1080 ) , 
    .X ( BUF_net_858 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_968 ( .A ( BUF_net_1084 ) , 
    .X ( BUF_net_968 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 ropt_h_inst_50845 ( 
    .A ( direct_interc_175_out[0] ) , .X ( ropt_net_2645 ) ) ;
sky130_fd_sc_hd__inv_4 cts_inv_1595218157 ( .A ( ctsbuf_net_372019 ) , 
    .Y ( ctsbuf_net_11983 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_482 ( .A ( BUF_net_831 ) , 
    .X ( BUF_net_482 ) ) ;
sky130_fd_sc_hd__inv_4 cts_inv_1595318158 ( .A ( ctsbuf_net_392021 ) , 
    .Y ( ctsbuf_net_21984 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_1083 ( .A ( BUF_net_1688 ) , 
    .X ( BUF_net_1083 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_1084 ( .A ( BUF_net_1188 ) , 
    .X ( BUF_net_1084 ) ) ;
sky130_fd_sc_hd__inv_4 cts_inv_1595418159 ( .A ( ctsbuf_net_372019 ) , 
    .Y ( ctsbuf_net_31985 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_487 ( .A ( BUF_net_955 ) , 
    .X ( BUF_net_487 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_488 ( .A ( Test_en[0] ) , 
    .X ( BUF_net_488 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_975 ( .A ( BUF_net_1368 ) , 
    .X ( BUF_net_975 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_976 ( .A ( BUF_net_1176 ) , 
    .X ( BUF_net_976 ) ) ;
sky130_fd_sc_hd__inv_4 cts_inv_1595518160 ( .A ( ctsbuf_net_372019 ) , 
    .Y ( ctsbuf_net_41986 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_1086 ( .A ( BUF_net_1194 ) , 
    .X ( BUF_net_1086 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_979 ( .A ( BUF_net_1086 ) , 
    .X ( BUF_net_979 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_494 ( .A ( BUF_net_822 ) , 
    .X ( BUF_net_494 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_980 ( .A ( BUF_net_1178 ) , 
    .X ( BUF_net_980 ) ) ;
sky130_fd_sc_hd__inv_4 cts_inv_1595618161 ( .A ( ctsbuf_net_382020 ) , 
    .Y ( ctsbuf_net_51987 ) ) ;
sky130_fd_sc_hd__inv_4 cts_inv_1595718162 ( .A ( ctsbuf_net_332015 ) , 
    .Y ( ctsbuf_net_61988 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_1185 ( .A ( BUF_net_1600 ) , 
    .X ( BUF_net_1185 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_499 ( .A ( BUF_net_828 ) , 
    .X ( BUF_net_499 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_500 ( .A ( Test_en[0] ) , 
    .X ( BUF_net_500 ) ) ;
sky130_fd_sc_hd__inv_4 cts_inv_1595818163 ( .A ( ctsbuf_net_332015 ) , 
    .Y ( ctsbuf_net_71989 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_1187 ( .A ( BUF_net_1359 ) , 
    .X ( BUF_net_1187 ) ) ;
sky130_fd_sc_hd__inv_4 cts_inv_1595918164 ( .A ( ctsbuf_net_332015 ) , 
    .Y ( ctsbuf_net_81990 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_1092 ( .A ( BUF_net_1447 ) , 
    .X ( BUF_net_1092 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_505 ( .A ( BUF_net_1608 ) , 
    .X ( BUF_net_505 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_506 ( .A ( BUF_net_822 ) , 
    .X ( BUF_net_506 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_1188 ( .A ( BUF_net_1350 ) , 
    .X ( BUF_net_1188 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_1094 ( .A ( BUF_net_1368 ) , 
    .X ( BUF_net_1094 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_1189 ( .A ( BUF_net_1508 ) , 
    .X ( BUF_net_1189 ) ) ;
sky130_fd_sc_hd__inv_4 cts_inv_1596018165 ( .A ( ctsbuf_net_372019 ) , 
    .Y ( ctsbuf_net_91991 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_511 ( .A ( BUF_net_1267 ) , 
    .X ( BUF_net_511 ) ) ;
sky130_fd_sc_hd__inv_4 cts_inv_1596118166 ( .A ( ctsbuf_net_382020 ) , 
    .Y ( ctsbuf_net_101992 ) ) ;
sky130_fd_sc_hd__inv_4 cts_inv_1596218167 ( .A ( ctsbuf_net_312013 ) , 
    .Y ( ctsbuf_net_111993 ) ) ;
sky130_fd_sc_hd__inv_4 cts_inv_1596318168 ( .A ( ctsbuf_net_382020 ) , 
    .Y ( ctsbuf_net_121994 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_1190 ( .A ( BUF_net_1573 ) , 
    .X ( BUF_net_1190 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_1368 ( .A ( BUF_net_1485 ) , 
    .X ( BUF_net_1368 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_517 ( .A ( BUF_net_1608 ) , 
    .X ( BUF_net_517 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_518 ( .A ( BUF_net_822 ) , 
    .X ( BUF_net_518 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_519 ( .A ( BUF_net_1743 ) , 
    .X ( BUF_net_519 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_1192 ( .A ( BUF_net_1360 ) , 
    .X ( BUF_net_1192 ) ) ;
sky130_fd_sc_hd__inv_4 cts_inv_1596418169 ( .A ( ctsbuf_net_332015 ) , 
    .Y ( ctsbuf_net_131995 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_1194 ( .A ( BUF_net_1351 ) , 
    .X ( BUF_net_1194 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_523 ( .A ( BUF_net_1267 ) , 
    .X ( BUF_net_523 ) ) ;
sky130_fd_sc_hd__inv_4 cts_inv_1596518170 ( .A ( ctsbuf_net_342016 ) , 
    .Y ( ctsbuf_net_141996 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_1195 ( .A ( BUF_net_1361 ) , 
    .X ( BUF_net_1195 ) ) ;
sky130_fd_sc_hd__inv_4 cts_inv_1596618171 ( .A ( ctsbuf_net_382020 ) , 
    .Y ( ctsbuf_net_151997 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_1197 ( .A ( BUF_net_1568 ) , 
    .X ( BUF_net_1197 ) ) ;
sky130_fd_sc_hd__inv_4 cts_inv_1596718172 ( .A ( ctsbuf_net_312013 ) , 
    .Y ( ctsbuf_net_161998 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_1199 ( .A ( BUF_net_1508 ) , 
    .X ( BUF_net_1199 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_530 ( .A ( BUF_net_822 ) , 
    .X ( BUF_net_530 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_1109 ( .A ( BUF_net_1737 ) , 
    .X ( BUF_net_1109 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_1200 ( .A ( BUF_net_1567 ) , 
    .X ( BUF_net_1200 ) ) ;
sky130_fd_sc_hd__inv_4 cts_inv_1596818173 ( .A ( ctsbuf_net_342016 ) , 
    .Y ( ctsbuf_net_171999 ) ) ;
sky130_fd_sc_hd__inv_4 cts_inv_1596918174 ( .A ( ctsbuf_net_312013 ) , 
    .Y ( ctsbuf_net_182000 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_535 ( .A ( BUF_net_1690 ) , 
    .X ( BUF_net_535 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_536 ( .A ( Test_en[0] ) , 
    .X ( BUF_net_536 ) ) ;
sky130_fd_sc_hd__inv_4 cts_inv_1597018175 ( .A ( ctsbuf_net_322014 ) , 
    .Y ( ctsbuf_net_192001 ) ) ;
sky130_fd_sc_hd__inv_4 cts_inv_1597118176 ( .A ( ctsbuf_net_352017 ) , 
    .Y ( ctsbuf_net_202002 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_1288 ( .A ( BUF_net_1373 ) , 
    .X ( BUF_net_1288 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_1206 ( .A ( BUF_net_1485 ) , 
    .X ( BUF_net_1206 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_541 ( .A ( BUF_net_1737 ) , 
    .X ( BUF_net_541 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_542 ( .A ( BUF_net_817 ) , 
    .X ( BUF_net_542 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_1207 ( .A ( BUF_net_1385 ) , 
    .X ( BUF_net_1207 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_1373 ( .A ( BUF_net_1446 ) , 
    .X ( BUF_net_1373 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_1209 ( .A ( BUF_net_1348 ) , 
    .X ( BUF_net_1209 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_1210 ( .A ( BUF_net_1574 ) , 
    .X ( BUF_net_1210 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_547 ( .A ( BUF_net_950 ) , 
    .X ( BUF_net_547 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_548 ( .A ( BUF_net_685 ) , 
    .X ( BUF_net_548 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_1444 ( .A ( BUF_net_1600 ) , 
    .X ( BUF_net_1444 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_1375 ( .A ( BUF_net_1551 ) , 
    .X ( BUF_net_1375 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_1376 ( .A ( BUF_net_1603 ) , 
    .X ( BUF_net_1376 ) ) ;
sky130_fd_sc_hd__inv_4 cts_inv_1597218177 ( .A ( ctsbuf_net_322014 ) , 
    .Y ( ctsbuf_net_212003 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_1445 ( .A ( BUF_net_1568 ) , 
    .X ( BUF_net_1445 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_554 ( .A ( BUF_net_817 ) , 
    .X ( BUF_net_554 ) ) ;
sky130_fd_sc_hd__clkinvlp_4 cts_inv_1597318178 ( .A ( ctsbuf_net_342016 ) , 
    .Y ( ctsbuf_net_222004 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_913 ( .A ( BUF_net_966 ) , 
    .X ( BUF_net_913 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_914 ( .A ( BUF_net_968 ) , 
    .X ( BUF_net_914 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_915 ( .A ( BUF_net_975 ) , 
    .X ( BUF_net_915 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_559 ( .A ( BUF_net_950 ) , 
    .X ( BUF_net_559 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_560 ( .A ( BUF_net_1261 ) , 
    .X ( BUF_net_560 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_916 ( .A ( BUF_net_979 ) , 
    .X ( BUF_net_916 ) ) ;
sky130_fd_sc_hd__inv_4 cts_inv_1597418179 ( .A ( ctsbuf_net_362018 ) , 
    .Y ( ctsbuf_net_232005 ) ) ;
sky130_fd_sc_hd__inv_4 cts_inv_1597518180 ( .A ( ctsbuf_net_342016 ) , 
    .Y ( ctsbuf_net_242006 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_1380 ( .A ( BUF_net_1607 ) , 
    .X ( BUF_net_1380 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_1381 ( .A ( BUF_net_1501 ) , 
    .X ( BUF_net_1381 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_566 ( .A ( BUF_net_813 ) , 
    .X ( BUF_net_566 ) ) ;
sky130_fd_sc_hd__inv_4 cts_inv_1597618181 ( .A ( ctsbuf_net_352017 ) , 
    .Y ( ctsbuf_net_252007 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_1382 ( .A ( BUF_net_1502 ) , 
    .X ( BUF_net_1382 ) ) ;
sky130_fd_sc_hd__inv_4 cts_inv_1597718182 ( .A ( ctsbuf_net_322014 ) , 
    .Y ( ctsbuf_net_262008 ) ) ;
sky130_fd_sc_hd__inv_4 cts_inv_1597818183 ( .A ( ctsbuf_net_362018 ) , 
    .Y ( ctsbuf_net_272009 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_571 ( .A ( BUF_net_948 ) , 
    .X ( BUF_net_571 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_572 ( .A ( BUF_net_802 ) , 
    .X ( BUF_net_572 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_573 ( .A ( BUF_net_1083 ) , 
    .X ( BUF_net_573 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_574 ( .A ( BUF_net_675 ) , 
    .X ( BUF_net_574 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_575 ( .A ( BUF_net_806 ) , 
    .X ( BUF_net_575 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_576 ( .A ( BUF_net_679 ) , 
    .X ( BUF_net_576 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_577 ( .A ( BUF_net_1037 ) , 
    .X ( BUF_net_577 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_578 ( .A ( BUF_net_813 ) , 
    .X ( BUF_net_578 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_579 ( .A ( BUF_net_805 ) , 
    .X ( BUF_net_579 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_580 ( .A ( BUF_net_672 ) , 
    .X ( BUF_net_580 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_581 ( .A ( BUF_net_671 ) , 
    .X ( BUF_net_581 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_582 ( .A ( BUF_net_804 ) , 
    .X ( BUF_net_582 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_583 ( .A ( BUF_net_948 ) , 
    .X ( BUF_net_583 ) ) ;
sky130_fd_sc_hd__inv_4 cts_inv_1597918184 ( .A ( ctsbuf_net_362018 ) , 
    .Y ( ctsbuf_net_282010 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_671 ( .A ( BUF_net_718 ) , 
    .X ( BUF_net_671 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_672 ( .A ( BUF_net_720 ) , 
    .X ( BUF_net_672 ) ) ;
sky130_fd_sc_hd__inv_4 cts_inv_1598018185 ( .A ( ctsbuf_net_362018 ) , 
    .Y ( ctsbuf_net_292011 ) ) ;
sky130_fd_sc_hd__inv_4 cts_inv_1598118186 ( .A ( ctsbuf_net_362018 ) , 
    .Y ( ctsbuf_net_302012 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_675 ( .A ( BUF_net_730 ) , 
    .X ( BUF_net_675 ) ) ;
sky130_fd_sc_hd__clkinvlp_4 cts_inv_1604018245 ( .A ( ctsbuf_net_402022 ) , 
    .Y ( ctsbuf_net_312013 ) ) ;
sky130_fd_sc_hd__clkinvlp_4 cts_inv_1604118246 ( .A ( ctsbuf_net_402022 ) , 
    .Y ( ctsbuf_net_322014 ) ) ;
sky130_fd_sc_hd__clkinvlp_4 cts_inv_1604218247 ( .A ( ctsbuf_net_402022 ) , 
    .Y ( ctsbuf_net_332015 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_679 ( .A ( BUF_net_726 ) , 
    .X ( BUF_net_679 ) ) ;
sky130_fd_sc_hd__inv_2 cts_inv_1604318248 ( .A ( ctsbuf_net_422024 ) , 
    .Y ( ctsbuf_net_342016 ) ) ;
sky130_fd_sc_hd__clkinvlp_2 cts_inv_1604418249 ( .A ( ctsbuf_net_412023 ) , 
    .Y ( ctsbuf_net_352017 ) ) ;
sky130_fd_sc_hd__inv_4 cts_inv_1604518250 ( .A ( ctsbuf_net_422024 ) , 
    .Y ( ctsbuf_net_362018 ) ) ;
sky130_fd_sc_hd__clkinvlp_4 cts_inv_1604618251 ( .A ( ctsbuf_net_402022 ) , 
    .Y ( ctsbuf_net_372019 ) ) ;
sky130_fd_sc_hd__inv_2 cts_inv_1604718252 ( .A ( ctsbuf_net_412023 ) , 
    .Y ( ctsbuf_net_382020 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_685 ( .A ( BUF_net_1261 ) , 
    .X ( BUF_net_685 ) ) ;
sky130_fd_sc_hd__clkinvlp_4 cts_inv_1604818253 ( .A ( ctsbuf_net_402022 ) , 
    .Y ( ctsbuf_net_392021 ) ) ;
sky130_fd_sc_hd__clkinvlp_4 cts_inv_1605918264 ( .A ( ctsbuf_net_432025 ) , 
    .Y ( ctsbuf_net_402022 ) ) ;
sky130_fd_sc_hd__clkinvlp_4 cts_inv_1606018265 ( .A ( ctsbuf_net_442026 ) , 
    .Y ( ctsbuf_net_412023 ) ) ;
sky130_fd_sc_hd__clkinvlp_4 cts_inv_1606118266 ( .A ( ctsbuf_net_432025 ) , 
    .Y ( ctsbuf_net_422024 ) ) ;
sky130_fd_sc_hd__inv_2 cts_inv_1606918274 ( .A ( clk[0] ) , 
    .Y ( ctsbuf_net_432025 ) ) ;
sky130_fd_sc_hd__clkinvlp_2 cts_inv_1607018275 ( .A ( clk[0] ) , 
    .Y ( ctsbuf_net_442026 ) ) ;
sky130_fd_sc_hd__inv_4 cts_inv_4658548790 ( .A ( ctsbuf_net_6172599 ) , 
    .Y ( ctsbuf_net_452027 ) ) ;
sky130_fd_sc_hd__inv_4 cts_inv_4658648791 ( .A ( ctsbuf_net_6082590 ) , 
    .Y ( ctsbuf_net_462028 ) ) ;
sky130_fd_sc_hd__inv_4 cts_inv_4658748792 ( .A ( ctsbuf_net_5842566 ) , 
    .Y ( ctsbuf_net_472029 ) ) ;
sky130_fd_sc_hd__clkinvlp_4 cts_inv_4658848793 ( .A ( ctsbuf_net_6172599 ) , 
    .Y ( ctsbuf_net_482030 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4658948794 ( .A ( ctsbuf_net_6172599 ) , 
    .Y ( ctsbuf_net_492031 ) ) ;
sky130_fd_sc_hd__inv_4 cts_inv_4659048795 ( .A ( ctsbuf_net_6172599 ) , 
    .Y ( ctsbuf_net_502032 ) ) ;
sky130_fd_sc_hd__inv_2 cts_inv_4659148796 ( .A ( ctsbuf_net_6082590 ) , 
    .Y ( ctsbuf_net_512033 ) ) ;
sky130_fd_sc_hd__inv_4 cts_inv_4659348798 ( .A ( ctsbuf_net_6082590 ) , 
    .Y ( ctsbuf_net_532035 ) ) ;
sky130_fd_sc_hd__clkinvlp_4 cts_inv_4659448799 ( .A ( ctsbuf_net_6172599 ) , 
    .Y ( ctsbuf_net_542036 ) ) ;
sky130_fd_sc_hd__clkinvlp_4 cts_inv_4659548800 ( .A ( ctsbuf_net_6312613 ) , 
    .Y ( ctsbuf_net_552037 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4659648801 ( .A ( ctsbuf_net_6082590 ) , 
    .Y ( ctsbuf_net_562038 ) ) ;
sky130_fd_sc_hd__inv_4 cts_inv_4660048805 ( .A ( ctsbuf_net_5842566 ) , 
    .Y ( ctsbuf_net_602042 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_708 ( .A ( BUF_net_719 ) , 
    .X ( BUF_net_708 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4660148806 ( .A ( ctsbuf_net_6172599 ) , 
    .Y ( ctsbuf_net_612043 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4660248807 ( .A ( ctsbuf_net_6172599 ) , 
    .Y ( ctsbuf_net_622044 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_711 ( .A ( BUF_net_727 ) , 
    .X ( BUF_net_711 ) ) ;
sky130_fd_sc_hd__clkinvlp_4 cts_inv_4660348808 ( .A ( ctsbuf_net_6052587 ) , 
    .Y ( ctsbuf_net_632045 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_713 ( .A ( BUF_net_731 ) , 
    .X ( BUF_net_713 ) ) ;
sky130_fd_sc_hd__inv_4 cts_inv_4660548810 ( .A ( ctsbuf_net_6052587 ) , 
    .Y ( ctsbuf_net_652047 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_802 ( .A ( BUF_net_1261 ) , 
    .X ( BUF_net_802 ) ) ;
sky130_fd_sc_hd__inv_8 cts_inv_4660648811 ( .A ( ctsbuf_net_6082590 ) , 
    .Y ( ctsbuf_net_662048 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_804 ( .A ( BUF_net_1600 ) , 
    .X ( BUF_net_804 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_805 ( .A ( BUF_net_1567 ) , 
    .X ( BUF_net_805 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_806 ( .A ( BUF_net_1485 ) , 
    .X ( BUF_net_806 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_1385 ( .A ( BUF_net_1694 ) , 
    .X ( BUF_net_1385 ) ) ;
sky130_fd_sc_hd__clkinvlp_4 cts_inv_4660848813 ( .A ( ctsbuf_net_5842566 ) , 
    .Y ( ctsbuf_net_682050 ) ) ;
sky130_fd_sc_hd__clkinvlp_4 cts_inv_4660948814 ( .A ( ctsbuf_net_6232605 ) , 
    .Y ( ctsbuf_net_692051 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_1446 ( .A ( BUF_net_1550 ) , 
    .X ( BUF_net_1446 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_813 ( .A ( BUF_net_1037 ) , 
    .X ( BUF_net_813 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_1447 ( .A ( BUF_net_1563 ) , 
    .X ( BUF_net_1447 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_1448 ( .A ( BUF_net_1567 ) , 
    .X ( BUF_net_1448 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_817 ( .A ( BUF_net_1737 ) , 
    .X ( BUF_net_817 ) ) ;
sky130_fd_sc_hd__inv_4 cts_inv_4661248817 ( .A ( ctsbuf_net_6082590 ) , 
    .Y ( ctsbuf_net_722054 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_1034 ( .A ( BUF_net_1567 ) , 
    .X ( BUF_net_1034 ) ) ;
sky130_fd_sc_hd__clkinvlp_4 cts_inv_4661348818 ( .A ( ctsbuf_net_6312613 ) , 
    .Y ( ctsbuf_net_732055 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_1035 ( .A ( BUF_net_1485 ) , 
    .X ( BUF_net_1035 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_822 ( .A ( BUF_net_1743 ) , 
    .X ( BUF_net_822 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4661448819 ( .A ( ctsbuf_net_6122594 ) , 
    .Y ( ctsbuf_net_742056 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_1037 ( .A ( BUF_net_1368 ) , 
    .X ( BUF_net_1037 ) ) ;
sky130_fd_sc_hd__inv_2 cts_inv_4661548820 ( .A ( ctsbuf_net_6072589 ) , 
    .Y ( ctsbuf_net_752057 ) ) ;
sky130_fd_sc_hd__clkinvlp_4 cts_inv_4661648821 ( .A ( ctsbuf_net_6082590 ) , 
    .Y ( ctsbuf_net_762058 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_1450 ( .A ( BUF_net_1547 ) , 
    .X ( BUF_net_1450 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_828 ( .A ( BUF_net_1267 ) , 
    .X ( BUF_net_828 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_1451 ( .A ( Test_en[0] ) , 
    .X ( BUF_net_1451 ) ) ;
sky130_fd_sc_hd__clkinvlp_4 cts_inv_4661748822 ( .A ( ctsbuf_net_6082590 ) , 
    .Y ( ctsbuf_net_772059 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_831 ( .A ( BUF_net_1573 ) , 
    .X ( BUF_net_831 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_1567 ( .A ( BUF_net_1716 ) , 
    .X ( BUF_net_1567 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4662048825 ( .A ( ctsbuf_net_6232605 ) , 
    .Y ( ctsbuf_net_802062 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_836 ( .A ( BUF_net_956 ) , 
    .X ( BUF_net_836 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4662148826 ( .A ( ctsbuf_net_6312613 ) , 
    .Y ( ctsbuf_net_812063 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_1568 ( .A ( BUF_net_1757 ) , 
    .X ( BUF_net_1568 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4662248827 ( .A ( ctsbuf_net_6052587 ) , 
    .Y ( ctsbuf_net_822064 ) ) ;
sky130_fd_sc_hd__clkinvlp_4 cts_inv_4662348828 ( .A ( ctsbuf_net_6052587 ) , 
    .Y ( ctsbuf_net_832065 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_841 ( .A ( BUF_net_1385 ) , 
    .X ( BUF_net_841 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_842 ( .A ( BUF_net_1574 ) , 
    .X ( BUF_net_842 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_843 ( .A ( BUF_net_850 ) , 
    .X ( BUF_net_843 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_844 ( .A ( BUF_net_960 ) , 
    .X ( BUF_net_844 ) ) ;
sky130_fd_sc_hd__inv_4 cts_inv_4662448829 ( .A ( ctsbuf_net_6312613 ) , 
    .Y ( ctsbuf_net_842066 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_1514 ( .A ( BUF_net_1607 ) , 
    .X ( BUF_net_1514 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_1515 ( .A ( BUF_net_1723 ) , 
    .X ( BUF_net_1515 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_1569 ( .A ( BUF_net_1768 ) , 
    .X ( BUF_net_1569 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_1570 ( .A ( BUF_net_1681 ) , 
    .X ( BUF_net_1570 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_948 ( .A ( BUF_net_1253 ) , 
    .X ( BUF_net_948 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_1460 ( .A ( BUF_net_1722 ) , 
    .X ( BUF_net_1460 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_950 ( .A ( BUF_net_1600 ) , 
    .X ( BUF_net_950 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_1571 ( .A ( BUF_net_1681 ) , 
    .X ( BUF_net_1571 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_1462 ( .A ( BUF_net_1694 ) , 
    .X ( BUF_net_1462 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_1615 ( .A ( BUF_net_1690 ) , 
    .X ( BUF_net_1615 ) ) ;
sky130_fd_sc_hd__inv_4 cts_inv_4662548830 ( .A ( ctsbuf_net_6312613 ) , 
    .Y ( ctsbuf_net_852067 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_955 ( .A ( BUF_net_1635 ) , 
    .X ( BUF_net_955 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_956 ( .A ( BUF_net_1568 ) , 
    .X ( BUF_net_956 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_1573 ( .A ( BUF_net_1722 ) , 
    .X ( BUF_net_1573 ) ) ;
sky130_fd_sc_hd__inv_4 cts_inv_4662648831 ( .A ( ctsbuf_net_6052587 ) , 
    .Y ( ctsbuf_net_862068 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_1466 ( .A ( BUF_net_1574 ) , 
    .X ( BUF_net_1466 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_960 ( .A ( BUF_net_1573 ) , 
    .X ( BUF_net_960 ) ) ;
sky130_fd_sc_hd__inv_4 cts_inv_4662748832 ( .A ( ctsbuf_net_6082590 ) , 
    .Y ( ctsbuf_net_872069 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_962 ( .A ( BUF_net_967 ) , 
    .X ( BUF_net_962 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_963 ( .A ( BUF_net_980 ) , 
    .X ( BUF_net_963 ) ) ;
sky130_fd_sc_hd__inv_2 cts_inv_4662848833 ( .A ( ctsbuf_net_6232605 ) , 
    .Y ( ctsbuf_net_882070 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_965 ( .A ( BUF_net_976 ) , 
    .X ( BUF_net_965 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_1521 ( .A ( BUF_net_1608 ) , 
    .X ( BUF_net_1521 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_1522 ( .A ( BUF_net_1603 ) , 
    .X ( BUF_net_1522 ) ) ;
sky130_fd_sc_hd__inv_4 cts_inv_4662948834 ( .A ( ctsbuf_net_5842566 ) , 
    .Y ( ctsbuf_net_892071 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_1523 ( .A ( BUF_net_1603 ) , 
    .X ( BUF_net_1523 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_1574 ( .A ( Test_en[0] ) , 
    .X ( BUF_net_1574 ) ) ;
sky130_fd_sc_hd__inv_4 cts_inv_4663048835 ( .A ( ctsbuf_net_5842566 ) , 
    .Y ( ctsbuf_net_902072 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_1253 ( .A ( BUF_net_1288 ) , 
    .X ( BUF_net_1253 ) ) ;
sky130_fd_sc_hd__clkinvlp_4 cts_inv_4663148836 ( .A ( ctsbuf_net_6112593 ) , 
    .Y ( ctsbuf_net_912073 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_1576 ( .A ( BUF_net_1752 ) , 
    .X ( BUF_net_1576 ) ) ;
sky130_fd_sc_hd__inv_12 cts_inv_4663248837 ( .A ( ctsbuf_net_6072589 ) , 
    .Y ( ctsbuf_net_922074 ) ) ;
sky130_fd_sc_hd__clkinvlp_4 cts_inv_4663348838 ( .A ( ctsbuf_net_6242606 ) , 
    .Y ( ctsbuf_net_932075 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_1688 ( .A ( Test_en[0] ) , 
    .X ( BUF_net_1688 ) ) ;
sky130_fd_sc_hd__clkinvlp_4 cts_inv_4663448839 ( .A ( ctsbuf_net_6232605 ) , 
    .Y ( ctsbuf_net_942076 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_1261 ( .A ( Test_en[0] ) , 
    .X ( BUF_net_1261 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4663748842 ( .A ( ctsbuf_net_6072589 ) , 
    .Y ( ctsbuf_net_972079 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_1076 ( .A ( BUF_net_1568 ) , 
    .X ( BUF_net_1076 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4663948844 ( .A ( ctsbuf_net_6122594 ) , 
    .Y ( ctsbuf_net_992081 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_1078 ( .A ( BUF_net_1189 ) , 
    .X ( BUF_net_1078 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_1080 ( .A ( BUF_net_1574 ) , 
    .X ( BUF_net_1080 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_1690 ( .A ( BUF_net_1757 ) , 
    .X ( BUF_net_1690 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_1175 ( .A ( Test_en[0] ) , 
    .X ( BUF_net_1175 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_1176 ( .A ( BUF_net_1192 ) , 
    .X ( BUF_net_1176 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_1177 ( .A ( BUF_net_1187 ) , 
    .X ( BUF_net_1177 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_1178 ( .A ( BUF_net_1195 ) , 
    .X ( BUF_net_1178 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_1657 ( .A ( BUF_net_1768 ) , 
    .X ( BUF_net_1657 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4664148846 ( .A ( ctsbuf_net_5842566 ) , 
    .Y ( ctsbuf_net_1012083 ) ) ;
sky130_fd_sc_hd__clkinvlp_4 cts_inv_4664248847 ( .A ( ctsbuf_net_6072589 ) , 
    .Y ( ctsbuf_net_1022084 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_1267 ( .A ( BUF_net_1607 ) , 
    .X ( BUF_net_1267 ) ) ;
sky130_fd_sc_hd__clkinvlp_4 cts_inv_4664448849 ( .A ( ctsbuf_net_6122594 ) , 
    .Y ( ctsbuf_net_1042086 ) ) ;
sky130_fd_sc_hd__clkinvlp_4 cts_inv_4664548850 ( .A ( ctsbuf_net_5892571 ) , 
    .Y ( ctsbuf_net_1052087 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_1626 ( .A ( Test_en[0] ) , 
    .X ( BUF_net_1626 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_1627 ( .A ( BUF_net_1716 ) , 
    .X ( BUF_net_1627 ) ) ;
sky130_fd_sc_hd__clkinvlp_4 cts_inv_4664648851 ( .A ( ctsbuf_net_5842566 ) , 
    .Y ( ctsbuf_net_1062088 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4664748852 ( .A ( ctsbuf_net_6242606 ) , 
    .Y ( ctsbuf_net_1072089 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4664848853 ( .A ( ctsbuf_net_6232605 ) , 
    .Y ( ctsbuf_net_1082090 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_1348 ( .A ( BUF_net_1688 ) , 
    .X ( BUF_net_1348 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_1485 ( .A ( Test_en[0] ) , 
    .X ( BUF_net_1485 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_1350 ( .A ( BUF_net_1375 ) , 
    .X ( BUF_net_1350 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_1351 ( .A ( BUF_net_1376 ) , 
    .X ( BUF_net_1351 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4664948854 ( .A ( ctsbuf_net_6052587 ) , 
    .Y ( ctsbuf_net_1092091 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_1715 ( .A ( BUF_net_1757 ) , 
    .X ( BUF_net_1715 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4665048855 ( .A ( ctsbuf_net_6052587 ) , 
    .Y ( ctsbuf_net_1102092 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_1631 ( .A ( BUF_net_1694 ) , 
    .X ( BUF_net_1631 ) ) ;
sky130_fd_sc_hd__inv_4 cts_inv_4665148856 ( .A ( ctsbuf_net_5942576 ) , 
    .Y ( ctsbuf_net_1112093 ) ) ;
sky130_fd_sc_hd__inv_6 cts_inv_4665248857 ( .A ( ctsbuf_net_6242606 ) , 
    .Y ( ctsbuf_net_1122094 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_1359 ( .A ( BUF_net_1380 ) , 
    .X ( BUF_net_1359 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_1360 ( .A ( BUF_net_1381 ) , 
    .X ( BUF_net_1360 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_1361 ( .A ( BUF_net_1382 ) , 
    .X ( BUF_net_1361 ) ) ;
sky130_fd_sc_hd__inv_6 cts_inv_4665448859 ( .A ( ctsbuf_net_6372619 ) , 
    .Y ( ctsbuf_net_1142096 ) ) ;
sky130_fd_sc_hd__inv_4 cts_inv_4665648861 ( .A ( ctsbuf_net_6242606 ) , 
    .Y ( ctsbuf_net_1162098 ) ) ;
sky130_fd_sc_hd__inv_6 cts_inv_4665748862 ( .A ( ctsbuf_net_6122594 ) , 
    .Y ( ctsbuf_net_1172099 ) ) ;
sky130_fd_sc_hd__inv_4 cts_inv_4665948864 ( .A ( ctsbuf_net_6112593 ) , 
    .Y ( ctsbuf_net_1192101 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_1694 ( .A ( Test_en[0] ) , 
    .X ( BUF_net_1694 ) ) ;
sky130_fd_sc_hd__inv_4 cts_inv_4666048865 ( .A ( ctsbuf_net_6112593 ) , 
    .Y ( ctsbuf_net_1202102 ) ) ;
sky130_fd_sc_hd__clkinvlp_4 cts_inv_4666148866 ( .A ( ctsbuf_net_6002582 ) , 
    .Y ( ctsbuf_net_1212103 ) ) ;
sky130_fd_sc_hd__clkinvlp_4 cts_inv_4666348868 ( .A ( ctsbuf_net_6372619 ) , 
    .Y ( ctsbuf_net_1232105 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_1547 ( .A ( BUF_net_1576 ) , 
    .X ( BUF_net_1547 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4666548870 ( .A ( ctsbuf_net_6072589 ) , 
    .Y ( ctsbuf_net_1252107 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4666648871 ( .A ( ctsbuf_net_6122594 ) , 
    .Y ( ctsbuf_net_1262108 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_1501 ( .A ( BUF_net_1608 ) , 
    .X ( BUF_net_1501 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_1502 ( .A ( BUF_net_1603 ) , 
    .X ( BUF_net_1502 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_1549 ( .A ( BUF_net_1688 ) , 
    .X ( BUF_net_1549 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_1550 ( .A ( BUF_net_1569 ) , 
    .X ( BUF_net_1550 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_1551 ( .A ( BUF_net_1571 ) , 
    .X ( BUF_net_1551 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_1634 ( .A ( Test_en[0] ) , 
    .X ( BUF_net_1634 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_1635 ( .A ( BUF_net_1685 ) , 
    .X ( BUF_net_1635 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_1508 ( .A ( BUF_net_1723 ) , 
    .X ( BUF_net_1508 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_1716 ( .A ( BUF_net_1737 ) , 
    .X ( BUF_net_1716 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4666848873 ( .A ( ctsbuf_net_5892571 ) , 
    .Y ( ctsbuf_net_1282110 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4666948874 ( .A ( ctsbuf_net_6112593 ) , 
    .Y ( ctsbuf_net_1292111 ) ) ;
sky130_fd_sc_hd__inv_2 cts_inv_4667148876 ( .A ( ctsbuf_net_5992581 ) , 
    .Y ( ctsbuf_net_1312113 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_1563 ( .A ( BUF_net_1570 ) , 
    .X ( BUF_net_1563 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_1600 ( .A ( BUF_net_1690 ) , 
    .X ( BUF_net_1600 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_1665 ( .A ( BUF_net_1722 ) , 
    .X ( BUF_net_1665 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_1603 ( .A ( Test_en[0] ) , 
    .X ( BUF_net_1603 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_1737 ( .A ( BUF_net_1752 ) , 
    .X ( BUF_net_1737 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4667848883 ( .A ( ctsbuf_net_6002582 ) , 
    .Y ( ctsbuf_net_1382120 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4667948884 ( .A ( ctsbuf_net_6242606 ) , 
    .Y ( ctsbuf_net_1392121 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_1607 ( .A ( BUF_net_1681 ) , 
    .X ( BUF_net_1607 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_1608 ( .A ( Test_en[0] ) , 
    .X ( BUF_net_1608 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4668048885 ( .A ( ctsbuf_net_6372619 ) , 
    .Y ( ctsbuf_net_1402122 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4668148886 ( .A ( ctsbuf_net_5942576 ) , 
    .Y ( ctsbuf_net_1412123 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_1722 ( .A ( BUF_net_1743 ) , 
    .X ( BUF_net_1722 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_1723 ( .A ( BUF_net_1762 ) , 
    .X ( BUF_net_1723 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_1724 ( .A ( Test_en[0] ) , 
    .X ( BUF_net_1724 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4668248887 ( .A ( ctsbuf_net_5942576 ) , 
    .Y ( ctsbuf_net_1422124 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_1725 ( .A ( Test_en[0] ) , 
    .X ( BUF_net_1725 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_1726 ( .A ( Test_en[0] ) , 
    .X ( BUF_net_1726 ) ) ;
sky130_fd_sc_hd__inv_4 cts_inv_4668348888 ( .A ( ctsbuf_net_5862568 ) , 
    .Y ( ctsbuf_net_1432125 ) ) ;
sky130_fd_sc_hd__inv_6 cts_inv_4668448889 ( .A ( ctsbuf_net_6412623 ) , 
    .Y ( ctsbuf_net_1442126 ) ) ;
sky130_fd_sc_hd__inv_6 cts_inv_4668648891 ( .A ( ctsbuf_net_6372619 ) , 
    .Y ( ctsbuf_net_1462128 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_1679 ( .A ( BUF_net_1688 ) , 
    .X ( BUF_net_1679 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_1727 ( .A ( BUF_net_1757 ) , 
    .X ( BUF_net_1727 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_1681 ( .A ( BUF_net_1762 ) , 
    .X ( BUF_net_1681 ) ) ;
sky130_fd_sc_hd__inv_4 cts_inv_4668748892 ( .A ( ctsbuf_net_5942576 ) , 
    .Y ( ctsbuf_net_1472129 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_1729 ( .A ( Test_en[0] ) , 
    .X ( BUF_net_1729 ) ) ;
sky130_fd_sc_hd__inv_4 cts_inv_4668848893 ( .A ( ctsbuf_net_6092591 ) , 
    .Y ( ctsbuf_net_1482130 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_1685 ( .A ( BUF_net_1757 ) , 
    .X ( BUF_net_1685 ) ) ;
sky130_fd_sc_hd__inv_4 cts_inv_4668948894 ( .A ( ctsbuf_net_6002582 ) , 
    .Y ( ctsbuf_net_1492131 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_1741 ( .A ( BUF_net_1762 ) , 
    .X ( BUF_net_1741 ) ) ;
sky130_fd_sc_hd__inv_6 cts_inv_4669248897 ( .A ( ctsbuf_net_5952577 ) , 
    .Y ( ctsbuf_net_1522134 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_1714 ( .A ( BUF_net_1723 ) , 
    .X ( BUF_net_1714 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_1743 ( .A ( BUF_net_1762 ) , 
    .X ( BUF_net_1743 ) ) ;
sky130_fd_sc_hd__inv_4 cts_inv_4669348898 ( .A ( ctsbuf_net_5852567 ) , 
    .Y ( ctsbuf_net_1532135 ) ) ;
sky130_fd_sc_hd__clkinvlp_4 cts_inv_4669448899 ( .A ( ctsbuf_net_6002582 ) , 
    .Y ( ctsbuf_net_1542136 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_1752 ( .A ( BUF_net_1786 ) , 
    .X ( BUF_net_1752 ) ) ;
sky130_fd_sc_hd__inv_4 cts_inv_4669948904 ( .A ( ctsbuf_net_5992581 ) , 
    .Y ( ctsbuf_net_1592141 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4670048905 ( .A ( ctsbuf_net_6092591 ) , 
    .Y ( ctsbuf_net_1602142 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_1757 ( .A ( BUF_net_1768 ) , 
    .X ( BUF_net_1757 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_1762 ( .A ( BUF_net_1786 ) , 
    .X ( BUF_net_1762 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_1768 ( .A ( BUF_net_1779 ) , 
    .X ( BUF_net_1768 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_1764 ( .A ( BUF_net_1786 ) , 
    .X ( BUF_net_1764 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4670248907 ( .A ( ctsbuf_net_6012583 ) , 
    .Y ( ctsbuf_net_1622144 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4670348908 ( .A ( ctsbuf_net_5952577 ) , 
    .Y ( ctsbuf_net_1632145 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_1786 ( .A ( Test_en[0] ) , 
    .X ( BUF_net_1786 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_1779 ( .A ( BUF_net_1786 ) , 
    .X ( BUF_net_1779 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4670548910 ( .A ( ctsbuf_net_6112593 ) , 
    .Y ( ctsbuf_net_1652147 ) ) ;
sky130_fd_sc_hd__clkinvlp_4 cts_inv_4670648911 ( .A ( ctsbuf_net_5862568 ) , 
    .Y ( ctsbuf_net_1662148 ) ) ;
sky130_fd_sc_hd__clkinvlp_4 cts_inv_4670948914 ( .A ( ctsbuf_net_6092591 ) , 
    .Y ( ctsbuf_net_1692151 ) ) ;
sky130_fd_sc_hd__bufinv_8 cts_inv_4671248917 ( .A ( ctsbuf_net_6122594 ) , 
    .Y ( ctsbuf_net_1722154 ) ) ;
sky130_fd_sc_hd__inv_4 cts_inv_4671648921 ( .A ( ctsbuf_net_5862568 ) , 
    .Y ( ctsbuf_net_1762158 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4671748922 ( .A ( ctsbuf_net_6002582 ) , 
    .Y ( ctsbuf_net_1772159 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4671848923 ( .A ( ctsbuf_net_6412623 ) , 
    .Y ( ctsbuf_net_1782160 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4671948924 ( .A ( ctsbuf_net_6322614 ) , 
    .Y ( ctsbuf_net_1792161 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4672048925 ( .A ( ctsbuf_net_6372619 ) , 
    .Y ( ctsbuf_net_1802162 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4672148926 ( .A ( ctsbuf_net_5942576 ) , 
    .Y ( ctsbuf_net_1812163 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4672248927 ( .A ( ctsbuf_net_5862568 ) , 
    .Y ( ctsbuf_net_1822164 ) ) ;
sky130_fd_sc_hd__inv_6 cts_inv_4672348928 ( .A ( ctsbuf_net_6002582 ) , 
    .Y ( ctsbuf_net_1832165 ) ) ;
sky130_fd_sc_hd__inv_6 cts_inv_4672548930 ( .A ( ctsbuf_net_6322614 ) , 
    .Y ( ctsbuf_net_1852167 ) ) ;
sky130_fd_sc_hd__inv_4 cts_inv_4672948934 ( .A ( ctsbuf_net_6002582 ) , 
    .Y ( ctsbuf_net_1892171 ) ) ;
sky130_fd_sc_hd__inv_6 cts_inv_4673248937 ( .A ( ctsbuf_net_6012583 ) , 
    .Y ( ctsbuf_net_1922174 ) ) ;
sky130_fd_sc_hd__clkinvlp_4 cts_inv_4673448939 ( .A ( ctsbuf_net_5822564 ) , 
    .Y ( ctsbuf_net_1942176 ) ) ;
sky130_fd_sc_hd__clkinvlp_4 cts_inv_4673748942 ( .A ( ctsbuf_net_6322614 ) , 
    .Y ( ctsbuf_net_1972179 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4674048945 ( .A ( ctsbuf_net_5992581 ) , 
    .Y ( ctsbuf_net_2002182 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4674148946 ( .A ( ctsbuf_net_5992581 ) , 
    .Y ( ctsbuf_net_2012183 ) ) ;
sky130_fd_sc_hd__clkinvlp_4 cts_inv_4674248947 ( .A ( ctsbuf_net_6382620 ) , 
    .Y ( ctsbuf_net_2022184 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4674348948 ( .A ( ctsbuf_net_6092591 ) , 
    .Y ( ctsbuf_net_2032185 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4674448949 ( .A ( ctsbuf_net_6012583 ) , 
    .Y ( ctsbuf_net_2042186 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4674648951 ( .A ( ctsbuf_net_5952577 ) , 
    .Y ( ctsbuf_net_2062188 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4674848953 ( .A ( ctsbuf_net_5862568 ) , 
    .Y ( ctsbuf_net_2082190 ) ) ;
sky130_fd_sc_hd__clkinvlp_4 cts_inv_4674948954 ( .A ( ctsbuf_net_5862568 ) , 
    .Y ( ctsbuf_net_2092191 ) ) ;
sky130_fd_sc_hd__inv_2 cts_inv_4675048955 ( .A ( ctsbuf_net_5852567 ) , 
    .Y ( ctsbuf_net_2102192 ) ) ;
sky130_fd_sc_hd__bufinv_8 cts_inv_4675348958 ( .A ( ctsbuf_net_5992581 ) , 
    .Y ( ctsbuf_net_2132195 ) ) ;
sky130_fd_sc_hd__clkinvlp_4 cts_inv_4675848963 ( .A ( ctsbuf_net_5952577 ) , 
    .Y ( ctsbuf_net_2182200 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4676148966 ( .A ( ctsbuf_net_5822564 ) , 
    .Y ( ctsbuf_net_2212203 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4676248967 ( .A ( ctsbuf_net_6002582 ) , 
    .Y ( ctsbuf_net_2222204 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4676348968 ( .A ( ctsbuf_net_6382620 ) , 
    .Y ( ctsbuf_net_2232205 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4676448969 ( .A ( ctsbuf_net_6322614 ) , 
    .Y ( ctsbuf_net_2242206 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4676548970 ( .A ( ctsbuf_net_5912573 ) , 
    .Y ( ctsbuf_net_2252207 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4676648971 ( .A ( ctsbuf_net_5882570 ) , 
    .Y ( ctsbuf_net_2262208 ) ) ;
sky130_fd_sc_hd__inv_6 cts_inv_4676748972 ( .A ( ctsbuf_net_5982580 ) , 
    .Y ( ctsbuf_net_2272209 ) ) ;
sky130_fd_sc_hd__inv_6 cts_inv_4676948974 ( .A ( ctsbuf_net_6332615 ) , 
    .Y ( ctsbuf_net_2292211 ) ) ;
sky130_fd_sc_hd__inv_4 cts_inv_4677448979 ( .A ( ctsbuf_net_5822564 ) , 
    .Y ( ctsbuf_net_2342216 ) ) ;
sky130_fd_sc_hd__inv_6 cts_inv_4677548980 ( .A ( ctsbuf_net_6152597 ) , 
    .Y ( ctsbuf_net_2352217 ) ) ;
sky130_fd_sc_hd__bufinv_8 cts_inv_4677748982 ( .A ( ctsbuf_net_6012583 ) , 
    .Y ( ctsbuf_net_2372219 ) ) ;
sky130_fd_sc_hd__clkinvlp_2 cts_inv_4677948984 ( .A ( ctsbuf_net_6022584 ) , 
    .Y ( ctsbuf_net_2392221 ) ) ;
sky130_fd_sc_hd__clkinvlp_4 cts_inv_4678048985 ( .A ( ctsbuf_net_5822564 ) , 
    .Y ( ctsbuf_net_2402222 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4678648991 ( .A ( ctsbuf_net_5852567 ) , 
    .Y ( ctsbuf_net_2462228 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4678748992 ( .A ( ctsbuf_net_5902572 ) , 
    .Y ( ctsbuf_net_2472229 ) ) ;
sky130_fd_sc_hd__clkinvlp_4 cts_inv_4678848993 ( .A ( ctsbuf_net_6412623 ) , 
    .Y ( ctsbuf_net_2482230 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4678948994 ( .A ( ctsbuf_net_6152597 ) , 
    .Y ( ctsbuf_net_2492231 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4679048995 ( .A ( ctsbuf_net_6032585 ) , 
    .Y ( ctsbuf_net_2502232 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4679248997 ( .A ( ctsbuf_net_6012583 ) , 
    .Y ( ctsbuf_net_2522234 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4679448999 ( .A ( ctsbuf_net_5872569 ) , 
    .Y ( ctsbuf_net_2542236 ) ) ;
sky130_fd_sc_hd__bufinv_8 cts_inv_4679849003 ( .A ( ctsbuf_net_5902572 ) , 
    .Y ( ctsbuf_net_2582240 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4680649011 ( .A ( ctsbuf_net_5822564 ) , 
    .Y ( ctsbuf_net_2662248 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4680749012 ( .A ( ctsbuf_net_5982580 ) , 
    .Y ( ctsbuf_net_2672249 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4680849013 ( .A ( ctsbuf_net_6342616 ) , 
    .Y ( ctsbuf_net_2682250 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4680949014 ( .A ( ctsbuf_net_6362618 ) , 
    .Y ( ctsbuf_net_2692251 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4681049015 ( .A ( ctsbuf_net_6332615 ) , 
    .Y ( ctsbuf_net_2702252 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4681149016 ( .A ( ctsbuf_net_5912573 ) , 
    .Y ( ctsbuf_net_2712253 ) ) ;
sky130_fd_sc_hd__inv_6 cts_inv_4681249017 ( .A ( ctsbuf_net_5822564 ) , 
    .Y ( ctsbuf_net_2722254 ) ) ;
sky130_fd_sc_hd__inv_6 cts_inv_4681449019 ( .A ( ctsbuf_net_6362618 ) , 
    .Y ( ctsbuf_net_2742256 ) ) ;
sky130_fd_sc_hd__inv_4 cts_inv_4681949024 ( .A ( ctsbuf_net_5822564 ) , 
    .Y ( ctsbuf_net_2792261 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4682049025 ( .A ( ctsbuf_net_5902572 ) , 
    .Y ( ctsbuf_net_2802262 ) ) ;
sky130_fd_sc_hd__clkinvlp_4 cts_inv_4682449029 ( .A ( ctsbuf_net_5822564 ) , 
    .Y ( ctsbuf_net_2842266 ) ) ;
sky130_fd_sc_hd__clkinvlp_4 cts_inv_4682549030 ( .A ( ctsbuf_net_5982580 ) , 
    .Y ( ctsbuf_net_2852267 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4683049035 ( .A ( ctsbuf_net_5852567 ) , 
    .Y ( ctsbuf_net_2902272 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4683149036 ( .A ( ctsbuf_net_5852567 ) , 
    .Y ( ctsbuf_net_2912273 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4683349038 ( .A ( ctsbuf_net_6152597 ) , 
    .Y ( ctsbuf_net_2932275 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4683449039 ( .A ( ctsbuf_net_6222604 ) , 
    .Y ( ctsbuf_net_2942276 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4683649041 ( .A ( ctsbuf_net_6032585 ) , 
    .Y ( ctsbuf_net_2962278 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4683849043 ( .A ( ctsbuf_net_5872569 ) , 
    .Y ( ctsbuf_net_2982280 ) ) ;
sky130_fd_sc_hd__inv_2 cts_inv_4684049045 ( .A ( ctsbuf_net_5832565 ) , 
    .Y ( ctsbuf_net_3002282 ) ) ;
sky130_fd_sc_hd__clkinvlp_4 cts_inv_4684349048 ( .A ( ctsbuf_net_5852567 ) , 
    .Y ( ctsbuf_net_3032285 ) ) ;
sky130_fd_sc_hd__clkinvlp_4 cts_inv_4684849053 ( .A ( ctsbuf_net_6032585 ) , 
    .Y ( ctsbuf_net_3082290 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4685149056 ( .A ( ctsbuf_net_6202602 ) , 
    .Y ( ctsbuf_net_3112293 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4685249057 ( .A ( ctsbuf_net_5822564 ) , 
    .Y ( ctsbuf_net_3122294 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4685349058 ( .A ( ctsbuf_net_6342616 ) , 
    .Y ( ctsbuf_net_3132295 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4685449059 ( .A ( ctsbuf_net_6362618 ) , 
    .Y ( ctsbuf_net_3142296 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4685549060 ( .A ( ctsbuf_net_6332615 ) , 
    .Y ( ctsbuf_net_3152297 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4685649061 ( .A ( ctsbuf_net_5912573 ) , 
    .Y ( ctsbuf_net_3162298 ) ) ;
sky130_fd_sc_hd__inv_6 cts_inv_4685749062 ( .A ( ctsbuf_net_6192601 ) , 
    .Y ( ctsbuf_net_3172299 ) ) ;
sky130_fd_sc_hd__inv_4 cts_inv_4685949064 ( .A ( ctsbuf_net_6402622 ) , 
    .Y ( ctsbuf_net_3192301 ) ) ;
sky130_fd_sc_hd__inv_4 cts_inv_4686249067 ( .A ( ctsbuf_net_5872569 ) , 
    .Y ( ctsbuf_net_3222304 ) ) ;
sky130_fd_sc_hd__inv_4 cts_inv_4686449069 ( .A ( ctsbuf_net_6202602 ) , 
    .Y ( ctsbuf_net_3242306 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4686549070 ( .A ( ctsbuf_net_6432625 ) , 
    .Y ( ctsbuf_net_3252307 ) ) ;
sky130_fd_sc_hd__inv_6 cts_inv_4686749072 ( .A ( ctsbuf_net_6222604 ) , 
    .Y ( ctsbuf_net_3272309 ) ) ;
sky130_fd_sc_hd__inv_4 cts_inv_4686949074 ( .A ( ctsbuf_net_5832565 ) , 
    .Y ( ctsbuf_net_3292311 ) ) ;
sky130_fd_sc_hd__clkinvlp_4 cts_inv_4687049075 ( .A ( ctsbuf_net_6202602 ) , 
    .Y ( ctsbuf_net_3302312 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4687649081 ( .A ( ctsbuf_net_6022584 ) , 
    .Y ( ctsbuf_net_3362318 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4687749082 ( .A ( ctsbuf_net_6432625 ) , 
    .Y ( ctsbuf_net_3372319 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4687949084 ( .A ( ctsbuf_net_5902572 ) , 
    .Y ( ctsbuf_net_3392321 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4688049085 ( .A ( ctsbuf_net_6152597 ) , 
    .Y ( ctsbuf_net_3402322 ) ) ;
sky130_fd_sc_hd__inv_16 cts_inv_4688249087 ( .A ( ctsbuf_net_6222604 ) , 
    .Y ( ctsbuf_net_3422324 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4688449089 ( .A ( ctsbuf_net_6032585 ) , 
    .Y ( ctsbuf_net_3442326 ) ) ;
sky130_fd_sc_hd__clkinvlp_4 cts_inv_4688549090 ( .A ( ctsbuf_net_5872569 ) , 
    .Y ( ctsbuf_net_3452327 ) ) ;
sky130_fd_sc_hd__clkinvlp_4 cts_inv_4688849093 ( .A ( ctsbuf_net_6432625 ) , 
    .Y ( ctsbuf_net_3482330 ) ) ;
sky130_fd_sc_hd__bufinv_8 cts_inv_4689049095 ( .A ( ctsbuf_net_5902572 ) , 
    .Y ( ctsbuf_net_3502332 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4689549100 ( .A ( ctsbuf_net_6202602 ) , 
    .Y ( ctsbuf_net_3552337 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4689649101 ( .A ( ctsbuf_net_6192601 ) , 
    .Y ( ctsbuf_net_3562338 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4689749102 ( .A ( ctsbuf_net_6342616 ) , 
    .Y ( ctsbuf_net_3572339 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4689849103 ( .A ( ctsbuf_net_6402622 ) , 
    .Y ( ctsbuf_net_3582340 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4689949104 ( .A ( ctsbuf_net_6392621 ) , 
    .Y ( ctsbuf_net_3592341 ) ) ;
sky130_fd_sc_hd__inv_4 cts_inv_4690049105 ( .A ( ctsbuf_net_6212603 ) , 
    .Y ( ctsbuf_net_3602342 ) ) ;
sky130_fd_sc_hd__inv_6 cts_inv_4690149106 ( .A ( ctsbuf_net_6202602 ) , 
    .Y ( ctsbuf_net_3612343 ) ) ;
sky130_fd_sc_hd__inv_6 cts_inv_4690349108 ( .A ( ctsbuf_net_6342616 ) , 
    .Y ( ctsbuf_net_3632345 ) ) ;
sky130_fd_sc_hd__inv_6 cts_inv_4690549110 ( .A ( ctsbuf_net_6392621 ) , 
    .Y ( ctsbuf_net_3652347 ) ) ;
sky130_fd_sc_hd__inv_4 cts_inv_4690849113 ( .A ( ctsbuf_net_6062588 ) , 
    .Y ( ctsbuf_net_3682350 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4690949114 ( .A ( ctsbuf_net_6262608 ) , 
    .Y ( ctsbuf_net_3692351 ) ) ;
sky130_fd_sc_hd__inv_6 cts_inv_4691149116 ( .A ( ctsbuf_net_6292611 ) , 
    .Y ( ctsbuf_net_3712353 ) ) ;
sky130_fd_sc_hd__clkinvlp_4 cts_inv_4691349118 ( .A ( ctsbuf_net_6062588 ) , 
    .Y ( ctsbuf_net_3732355 ) ) ;
sky130_fd_sc_hd__clkinvlp_4 cts_inv_4691849123 ( .A ( ctsbuf_net_6212603 ) , 
    .Y ( ctsbuf_net_3782360 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4691949124 ( .A ( ctsbuf_net_5832565 ) , 
    .Y ( ctsbuf_net_3792361 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4692049125 ( .A ( ctsbuf_net_6262608 ) , 
    .Y ( ctsbuf_net_3802362 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4692249127 ( .A ( ctsbuf_net_6432625 ) , 
    .Y ( ctsbuf_net_3822364 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4692349128 ( .A ( ctsbuf_net_6252607 ) , 
    .Y ( ctsbuf_net_3832365 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4692549130 ( .A ( ctsbuf_net_6222604 ) , 
    .Y ( ctsbuf_net_3852367 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4692649131 ( .A ( ctsbuf_net_6212603 ) , 
    .Y ( ctsbuf_net_3862368 ) ) ;
sky130_fd_sc_hd__inv_2 cts_inv_4692849133 ( .A ( ctsbuf_net_5832565 ) , 
    .Y ( ctsbuf_net_3882370 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4693849143 ( .A ( ctsbuf_net_6062588 ) , 
    .Y ( ctsbuf_net_3982380 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4693949144 ( .A ( ctsbuf_net_6192601 ) , 
    .Y ( ctsbuf_net_3992381 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4694049145 ( .A ( ctsbuf_net_6352617 ) , 
    .Y ( ctsbuf_net_4002382 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4694149146 ( .A ( ctsbuf_net_6402622 ) , 
    .Y ( ctsbuf_net_4012383 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4694249147 ( .A ( ctsbuf_net_6402622 ) , 
    .Y ( ctsbuf_net_4022384 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4694349148 ( .A ( ctsbuf_net_6212603 ) , 
    .Y ( ctsbuf_net_4032385 ) ) ;
sky130_fd_sc_hd__inv_6 cts_inv_4694449149 ( .A ( ctsbuf_net_6062588 ) , 
    .Y ( ctsbuf_net_4042386 ) ) ;
sky130_fd_sc_hd__inv_6 cts_inv_4694649151 ( .A ( ctsbuf_net_6352617 ) , 
    .Y ( ctsbuf_net_4062388 ) ) ;
sky130_fd_sc_hd__inv_4 cts_inv_4695149156 ( .A ( ctsbuf_net_6042586 ) , 
    .Y ( ctsbuf_net_4112393 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4695249157 ( .A ( ctsbuf_net_5962578 ) , 
    .Y ( ctsbuf_net_4122394 ) ) ;
sky130_fd_sc_hd__inv_6 cts_inv_4695449159 ( .A ( ctsbuf_net_6252607 ) , 
    .Y ( ctsbuf_net_4142396 ) ) ;
sky130_fd_sc_hd__clkinvlp_4 cts_inv_4695649161 ( .A ( ctsbuf_net_5832565 ) , 
    .Y ( ctsbuf_net_4162398 ) ) ;
sky130_fd_sc_hd__inv_4 cts_inv_4695749162 ( .A ( ctsbuf_net_6042586 ) , 
    .Y ( ctsbuf_net_4172399 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4696349168 ( .A ( ctsbuf_net_5832565 ) , 
    .Y ( ctsbuf_net_4232405 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4696449169 ( .A ( ctsbuf_net_5962578 ) , 
    .Y ( ctsbuf_net_4242406 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4696649171 ( .A ( ctsbuf_net_6262608 ) , 
    .Y ( ctsbuf_net_4262408 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4696749172 ( .A ( ctsbuf_net_6252607 ) , 
    .Y ( ctsbuf_net_4272409 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4696949174 ( .A ( ctsbuf_net_6292611 ) , 
    .Y ( ctsbuf_net_4292411 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4697149176 ( .A ( ctsbuf_net_6292611 ) , 
    .Y ( ctsbuf_net_4312413 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4698249187 ( .A ( ctsbuf_net_6042586 ) , 
    .Y ( ctsbuf_net_4422424 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4698349188 ( .A ( ctsbuf_net_6062588 ) , 
    .Y ( ctsbuf_net_4432425 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4698449189 ( .A ( ctsbuf_net_6352617 ) , 
    .Y ( ctsbuf_net_4442426 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4698549190 ( .A ( ctsbuf_net_6182600 ) , 
    .Y ( ctsbuf_net_4452427 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4698649191 ( .A ( ctsbuf_net_6132595 ) , 
    .Y ( ctsbuf_net_4462428 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4698749192 ( .A ( ctsbuf_net_6132595 ) , 
    .Y ( ctsbuf_net_4472429 ) ) ;
sky130_fd_sc_hd__inv_6 cts_inv_4698849193 ( .A ( ctsbuf_net_6042586 ) , 
    .Y ( ctsbuf_net_4482430 ) ) ;
sky130_fd_sc_hd__clkinvlp_4 cts_inv_4699049195 ( .A ( ctsbuf_net_6352617 ) , 
    .Y ( ctsbuf_net_4502432 ) ) ;
sky130_fd_sc_hd__inv_4 cts_inv_4699149196 ( .A ( ctsbuf_net_6402622 ) , 
    .Y ( ctsbuf_net_4512433 ) ) ;
sky130_fd_sc_hd__inv_4 cts_inv_4699249197 ( .A ( ctsbuf_net_6132595 ) , 
    .Y ( ctsbuf_net_4522434 ) ) ;
sky130_fd_sc_hd__inv_2 cts_inv_4699449199 ( .A ( ctsbuf_net_6042586 ) , 
    .Y ( ctsbuf_net_4542436 ) ) ;
sky130_fd_sc_hd__bufinv_8 cts_inv_4699549200 ( .A ( ctsbuf_net_5962578 ) , 
    .Y ( ctsbuf_net_4552437 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4699649201 ( .A ( ctsbuf_net_5962578 ) , 
    .Y ( ctsbuf_net_4562438 ) ) ;
sky130_fd_sc_hd__inv_4 cts_inv_4699749202 ( .A ( ctsbuf_net_6272609 ) , 
    .Y ( ctsbuf_net_4572439 ) ) ;
sky130_fd_sc_hd__inv_6 cts_inv_4699849203 ( .A ( ctsbuf_net_6252607 ) , 
    .Y ( ctsbuf_net_4582440 ) ) ;
sky130_fd_sc_hd__clkinvlp_4 cts_inv_4700349208 ( .A ( ctsbuf_net_6132595 ) , 
    .Y ( ctsbuf_net_4632445 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4700549210 ( .A ( ctsbuf_net_5832565 ) , 
    .Y ( ctsbuf_net_4652447 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4700649211 ( .A ( ctsbuf_net_5962578 ) , 
    .Y ( ctsbuf_net_4662448 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4700849213 ( .A ( ctsbuf_net_6422624 ) , 
    .Y ( ctsbuf_net_4682450 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4700949214 ( .A ( ctsbuf_net_6272609 ) , 
    .Y ( ctsbuf_net_4692451 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4701149216 ( .A ( ctsbuf_net_6252607 ) , 
    .Y ( ctsbuf_net_4712453 ) ) ;
sky130_fd_sc_hd__clkinvlp_4 cts_inv_4701249217 ( .A ( ctsbuf_net_6132595 ) , 
    .Y ( ctsbuf_net_4722454 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4701349218 ( .A ( ctsbuf_net_6282610 ) , 
    .Y ( ctsbuf_net_4732455 ) ) ;
sky130_fd_sc_hd__inv_4 cts_inv_4701549220 ( .A ( ctsbuf_net_6142596 ) , 
    .Y ( ctsbuf_net_4752457 ) ) ;
sky130_fd_sc_hd__clkinvlp_4 cts_inv_4701649221 ( .A ( ctsbuf_net_5962578 ) , 
    .Y ( ctsbuf_net_4762458 ) ) ;
sky130_fd_sc_hd__bufinv_8 cts_inv_4701849223 ( .A ( ctsbuf_net_6272609 ) , 
    .Y ( ctsbuf_net_4782460 ) ) ;
sky130_fd_sc_hd__clkinvlp_2 cts_inv_4702349228 ( .A ( ctsbuf_net_6142596 ) , 
    .Y ( ctsbuf_net_4832465 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4702449229 ( .A ( ctsbuf_net_6042586 ) , 
    .Y ( ctsbuf_net_4842466 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4702549230 ( .A ( ctsbuf_net_6102592 ) , 
    .Y ( ctsbuf_net_4852467 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4702649231 ( .A ( ctsbuf_net_6352617 ) , 
    .Y ( ctsbuf_net_4862468 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4702749232 ( .A ( ctsbuf_net_6182600 ) , 
    .Y ( ctsbuf_net_4872469 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4702849233 ( .A ( ctsbuf_net_6132595 ) , 
    .Y ( ctsbuf_net_4882470 ) ) ;
sky130_fd_sc_hd__inv_4 cts_inv_4702949234 ( .A ( ctsbuf_net_6042586 ) , 
    .Y ( ctsbuf_net_4892471 ) ) ;
sky130_fd_sc_hd__inv_6 cts_inv_4703049235 ( .A ( ctsbuf_net_6102592 ) , 
    .Y ( ctsbuf_net_4902472 ) ) ;
sky130_fd_sc_hd__inv_6 cts_inv_4703249237 ( .A ( ctsbuf_net_6302612 ) , 
    .Y ( ctsbuf_net_4922474 ) ) ;
sky130_fd_sc_hd__inv_4 cts_inv_4703349238 ( .A ( ctsbuf_net_6132595 ) , 
    .Y ( ctsbuf_net_4932475 ) ) ;
sky130_fd_sc_hd__inv_4 cts_inv_4703449239 ( .A ( ctsbuf_net_6042586 ) , 
    .Y ( ctsbuf_net_4942476 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4703549240 ( .A ( ctsbuf_net_6142596 ) , 
    .Y ( ctsbuf_net_4952477 ) ) ;
sky130_fd_sc_hd__inv_6 cts_inv_4703749242 ( .A ( ctsbuf_net_6252607 ) , 
    .Y ( ctsbuf_net_4972479 ) ) ;
sky130_fd_sc_hd__inv_4 cts_inv_4703849243 ( .A ( ctsbuf_net_6282610 ) , 
    .Y ( ctsbuf_net_4982480 ) ) ;
sky130_fd_sc_hd__clkinvlp_4 cts_inv_4704249247 ( .A ( ctsbuf_net_6132595 ) , 
    .Y ( ctsbuf_net_5022484 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4704349248 ( .A ( ctsbuf_net_6142596 ) , 
    .Y ( ctsbuf_net_5032485 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4704449249 ( .A ( ctsbuf_net_6162598 ) , 
    .Y ( ctsbuf_net_5042486 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4704549250 ( .A ( ctsbuf_net_6422624 ) , 
    .Y ( ctsbuf_net_5052487 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4704749252 ( .A ( ctsbuf_net_6272609 ) , 
    .Y ( ctsbuf_net_5072489 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4704849253 ( .A ( ctsbuf_net_6132595 ) , 
    .Y ( ctsbuf_net_5082490 ) ) ;
sky130_fd_sc_hd__clkinvlp_4 cts_inv_4704949254 ( .A ( ctsbuf_net_6132595 ) , 
    .Y ( ctsbuf_net_5092491 ) ) ;
sky130_fd_sc_hd__clkinvlp_4 cts_inv_4705549260 ( .A ( ctsbuf_net_6132595 ) , 
    .Y ( ctsbuf_net_5152497 ) ) ;
sky130_fd_sc_hd__inv_2 cts_inv_4705649261 ( .A ( ctsbuf_net_6142596 ) , 
    .Y ( ctsbuf_net_5162498 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4705749262 ( .A ( ctsbuf_net_6042586 ) , 
    .Y ( ctsbuf_net_5172499 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4705849263 ( .A ( ctsbuf_net_6102592 ) , 
    .Y ( ctsbuf_net_5182500 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4705949264 ( .A ( ctsbuf_net_6182600 ) , 
    .Y ( ctsbuf_net_5192501 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4706049265 ( .A ( ctsbuf_net_6302612 ) , 
    .Y ( ctsbuf_net_5202502 ) ) ;
sky130_fd_sc_hd__inv_6 cts_inv_4706149266 ( .A ( ctsbuf_net_6102592 ) , 
    .Y ( ctsbuf_net_5212503 ) ) ;
sky130_fd_sc_hd__inv_4 cts_inv_4706249267 ( .A ( ctsbuf_net_6182600 ) , 
    .Y ( ctsbuf_net_5222504 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4706449269 ( .A ( ctsbuf_net_6132595 ) , 
    .Y ( ctsbuf_net_5242506 ) ) ;
sky130_fd_sc_hd__inv_2 cts_inv_4706549270 ( .A ( ctsbuf_net_6102592 ) , 
    .Y ( ctsbuf_net_5252507 ) ) ;
sky130_fd_sc_hd__inv_4 cts_inv_4706649271 ( .A ( ctsbuf_net_6162598 ) , 
    .Y ( ctsbuf_net_5262508 ) ) ;
sky130_fd_sc_hd__inv_6 cts_inv_4706749272 ( .A ( ctsbuf_net_6442626 ) , 
    .Y ( ctsbuf_net_5272509 ) ) ;
sky130_fd_sc_hd__inv_4 cts_inv_4706849273 ( .A ( ctsbuf_net_6272609 ) , 
    .Y ( ctsbuf_net_5282510 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4707249277 ( .A ( ctsbuf_net_6142596 ) , 
    .Y ( ctsbuf_net_5322514 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4707349278 ( .A ( ctsbuf_net_6162598 ) , 
    .Y ( ctsbuf_net_5332515 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4707549280 ( .A ( ctsbuf_net_6422624 ) , 
    .Y ( ctsbuf_net_5352517 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4707749282 ( .A ( ctsbuf_net_6302612 ) , 
    .Y ( ctsbuf_net_5372519 ) ) ;
sky130_fd_sc_hd__clkinvlp_4 cts_inv_4707849283 ( .A ( ctsbuf_net_6302612 ) , 
    .Y ( ctsbuf_net_5382520 ) ) ;
sky130_fd_sc_hd__inv_4 cts_inv_4707949284 ( .A ( ctsbuf_net_6162598 ) , 
    .Y ( ctsbuf_net_5392521 ) ) ;
sky130_fd_sc_hd__clkinvlp_4 cts_inv_4708049285 ( .A ( ctsbuf_net_6162598 ) , 
    .Y ( ctsbuf_net_5402522 ) ) ;
sky130_fd_sc_hd__clkinvlp_2 cts_inv_4708449289 ( .A ( ctsbuf_net_6162598 ) , 
    .Y ( ctsbuf_net_5442526 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4708549290 ( .A ( ctsbuf_net_5972579 ) , 
    .Y ( ctsbuf_net_5452527 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4708649291 ( .A ( ctsbuf_net_6182600 ) , 
    .Y ( ctsbuf_net_5462528 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4708749292 ( .A ( ctsbuf_net_6302612 ) , 
    .Y ( ctsbuf_net_5472529 ) ) ;
sky130_fd_sc_hd__inv_4 cts_inv_4709149296 ( .A ( ctsbuf_net_5972579 ) , 
    .Y ( ctsbuf_net_5512533 ) ) ;
sky130_fd_sc_hd__inv_6 cts_inv_4709249297 ( .A ( ctsbuf_net_6162598 ) , 
    .Y ( ctsbuf_net_5522534 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4709649301 ( .A ( ctsbuf_net_6162598 ) , 
    .Y ( ctsbuf_net_5562538 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4709749302 ( .A ( ctsbuf_net_5922574 ) , 
    .Y ( ctsbuf_net_5572539 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4709949304 ( .A ( ctsbuf_net_6422624 ) , 
    .Y ( ctsbuf_net_5592541 ) ) ;
sky130_fd_sc_hd__inv_2 cts_inv_4710449309 ( .A ( ctsbuf_net_5932575 ) , 
    .Y ( ctsbuf_net_5642546 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4710549310 ( .A ( ctsbuf_net_5972579 ) , 
    .Y ( ctsbuf_net_5652547 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4710649311 ( .A ( ctsbuf_net_5922574 ) , 
    .Y ( ctsbuf_net_5662548 ) ) ;
sky130_fd_sc_hd__inv_4 cts_inv_4710749312 ( .A ( ctsbuf_net_5972579 ) , 
    .Y ( ctsbuf_net_5672549 ) ) ;
sky130_fd_sc_hd__inv_4 cts_inv_4710849313 ( .A ( ctsbuf_net_5922574 ) , 
    .Y ( ctsbuf_net_5682550 ) ) ;
sky130_fd_sc_hd__inv_4 cts_inv_4710949314 ( .A ( ctsbuf_net_5972579 ) , 
    .Y ( ctsbuf_net_5692551 ) ) ;
sky130_fd_sc_hd__inv_4 cts_inv_4711049315 ( .A ( ctsbuf_net_5922574 ) , 
    .Y ( ctsbuf_net_5702552 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4711249317 ( .A ( ctsbuf_net_5932575 ) , 
    .Y ( ctsbuf_net_5722554 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4711349318 ( .A ( ctsbuf_net_5922574 ) , 
    .Y ( ctsbuf_net_5732555 ) ) ;
sky130_fd_sc_hd__inv_4 cts_inv_4711549320 ( .A ( ctsbuf_net_5932575 ) , 
    .Y ( ctsbuf_net_5752557 ) ) ;
sky130_fd_sc_hd__clkinvlp_4 cts_inv_4711649321 ( .A ( ctsbuf_net_5922574 ) , 
    .Y ( ctsbuf_net_5762558 ) ) ;
sky130_fd_sc_hd__clkinvlp_2 cts_inv_4711749322 ( .A ( ctsbuf_net_5932575 ) , 
    .Y ( ctsbuf_net_5772559 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4711849323 ( .A ( ctsbuf_net_5972579 ) , 
    .Y ( ctsbuf_net_5782560 ) ) ;
sky130_fd_sc_hd__inv_4 cts_inv_4711949324 ( .A ( ctsbuf_net_5932575 ) , 
    .Y ( ctsbuf_net_5792561 ) ) ;
sky130_fd_sc_hd__inv_4 cts_inv_4712049325 ( .A ( ctsbuf_net_5932575 ) , 
    .Y ( ctsbuf_net_5802562 ) ) ;
sky130_fd_sc_hd__clkinv_4 cts_inv_4712149326 ( .A ( ctsbuf_net_5932575 ) , 
    .Y ( ctsbuf_net_5812563 ) ) ;
sky130_fd_sc_hd__clkinv_8 cts_inv_4659248797_4712249327 ( 
    .A ( SYNOPSYS_UNCONNECTED_1 ) , .Y ( SYNOPSYS_UNCONNECTED_2 ) ) ;
sky130_fd_sc_hd__clkinv_16 cts_inv_4661148816_4712349328 ( 
    .A ( SYNOPSYS_UNCONNECTED_3 ) , .Y ( p_abuf1 ) ) ;
sky130_fd_sc_hd__clkinv_16 cts_inv_4659848803_4712449329 ( 
    .A ( SYNOPSYS_UNCONNECTED_4 ) , .Y ( p_abuf0 ) ) ;
sky130_fd_sc_hd__inv_12 cts_inv_4660748812_4712549330 ( 
    .A ( SYNOPSYS_UNCONNECTED_5 ) , .Y ( SYNOPSYS_UNCONNECTED_6 ) ) ;
sky130_fd_sc_hd__inv_8 cts_inv_4663848843_4712649331 ( 
    .A ( SYNOPSYS_UNCONNECTED_7 ) , .Y ( SYNOPSYS_UNCONNECTED_8 ) ) ;
sky130_fd_sc_hd__inv_8 cts_inv_4661048815_4712749332 ( 
    .A ( SYNOPSYS_UNCONNECTED_9 ) , .Y ( SYNOPSYS_UNCONNECTED_10 ) ) ;
sky130_fd_sc_hd__inv_8 cts_inv_4661948824_4712849333 ( 
    .A ( SYNOPSYS_UNCONNECTED_11 ) , .Y ( SYNOPSYS_UNCONNECTED_12 ) ) ;
sky130_fd_sc_hd__inv_8 cts_inv_4664048845_4712949334 ( 
    .A ( SYNOPSYS_UNCONNECTED_13 ) , .Y ( SYNOPSYS_UNCONNECTED_14 ) ) ;
sky130_fd_sc_hd__inv_6 cts_inv_4659748802_4713049335 ( 
    .A ( SYNOPSYS_UNCONNECTED_15 ) , .Y ( SYNOPSYS_UNCONNECTED_16 ) ) ;
sky130_fd_sc_hd__inv_8 cts_inv_4663548840_4713149336 ( 
    .A ( SYNOPSYS_UNCONNECTED_17 ) , .Y ( SYNOPSYS_UNCONNECTED_18 ) ) ;
sky130_fd_sc_hd__inv_8 cts_inv_4663648841_4713249337 ( 
    .A ( SYNOPSYS_UNCONNECTED_19 ) , .Y ( SYNOPSYS_UNCONNECTED_20 ) ) ;
sky130_fd_sc_hd__inv_12 cts_inv_4664348848_4713349338 ( 
    .A ( SYNOPSYS_UNCONNECTED_21 ) , .Y ( SYNOPSYS_UNCONNECTED_22 ) ) ;
sky130_fd_sc_hd__inv_12 cts_inv_4659948804_4713449339 ( 
    .A ( SYNOPSYS_UNCONNECTED_23 ) , .Y ( SYNOPSYS_UNCONNECTED_24 ) ) ;
sky130_fd_sc_hd__inv_8 cts_inv_4661848823_4713549340 ( 
    .A ( SYNOPSYS_UNCONNECTED_25 ) , .Y ( SYNOPSYS_UNCONNECTED_26 ) ) ;
sky130_fd_sc_hd__inv_12 cts_inv_4697449179_4713649341 ( 
    .A ( SYNOPSYS_UNCONNECTED_27 ) , .Y ( p_abuf19 ) ) ;
sky130_fd_sc_hd__inv_8 cts_inv_4697349178_4713749342 ( 
    .A ( SYNOPSYS_UNCONNECTED_28 ) , .Y ( SYNOPSYS_UNCONNECTED_29 ) ) ;
sky130_fd_sc_hd__inv_6 cts_inv_4667648881_4713849343 ( 
    .A ( SYNOPSYS_UNCONNECTED_30 ) , .Y ( SYNOPSYS_UNCONNECTED_31 ) ) ;
sky130_fd_sc_hd__inv_8 cts_inv_4705049255_4713949344 ( 
    .A ( SYNOPSYS_UNCONNECTED_32 ) , .Y ( SYNOPSYS_UNCONNECTED_33 ) ) ;
sky130_fd_sc_hd__inv_8 cts_inv_4711149316_4714049345 ( 
    .A ( SYNOPSYS_UNCONNECTED_34 ) , .Y ( SYNOPSYS_UNCONNECTED_35 ) ) ;
sky130_fd_sc_hd__inv_8 cts_inv_4709449299_4714149346 ( 
    .A ( SYNOPSYS_UNCONNECTED_36 ) , .Y ( SYNOPSYS_UNCONNECTED_37 ) ) ;
sky130_fd_sc_hd__clkinv_16 cts_inv_4701949224_4714249347 ( 
    .A ( SYNOPSYS_UNCONNECTED_38 ) , .Y ( SYNOPSYS_UNCONNECTED_39 ) ) ;
sky130_fd_sc_hd__inv_8 cts_inv_4697649181_4714349348 ( 
    .A ( SYNOPSYS_UNCONNECTED_40 ) , .Y ( p_abuf20 ) ) ;
sky130_fd_sc_hd__clkinv_8 cts_inv_4678148986_4714449349 ( 
    .A ( SYNOPSYS_UNCONNECTED_41 ) , .Y ( SYNOPSYS_UNCONNECTED_42 ) ) ;
sky130_fd_sc_hd__inv_8 cts_inv_4710149306_4714549350 ( 
    .A ( SYNOPSYS_UNCONNECTED_43 ) , .Y ( SYNOPSYS_UNCONNECTED_44 ) ) ;
sky130_fd_sc_hd__inv_16 cts_inv_4688749092_4714649351 ( 
    .A ( SYNOPSYS_UNCONNECTED_45 ) , .Y ( SYNOPSYS_UNCONNECTED_46 ) ) ;
sky130_fd_sc_hd__inv_8 cts_inv_4684249047_4714749352 ( 
    .A ( SYNOPSYS_UNCONNECTED_47 ) , .Y ( SYNOPSYS_UNCONNECTED_48 ) ) ;
sky130_fd_sc_hd__inv_8 cts_inv_4669748902_4714849353 ( 
    .A ( SYNOPSYS_UNCONNECTED_49 ) , .Y ( SYNOPSYS_UNCONNECTED_50 ) ) ;
sky130_fd_sc_hd__inv_16 cts_inv_4675648961_4714949354 ( 
    .A ( SYNOPSYS_UNCONNECTED_51 ) , .Y ( SYNOPSYS_UNCONNECTED_52 ) ) ;
sky130_fd_sc_hd__clkinv_16 cts_inv_4666748872_4715049355 ( 
    .A ( SYNOPSYS_UNCONNECTED_53 ) , .Y ( SYNOPSYS_UNCONNECTED_54 ) ) ;
sky130_fd_sc_hd__inv_8 cts_inv_4669648901_4715149356 ( 
    .A ( SYNOPSYS_UNCONNECTED_55 ) , .Y ( SYNOPSYS_UNCONNECTED_56 ) ) ;
sky130_fd_sc_hd__inv_8 cts_inv_4676048965_4715249357 ( 
    .A ( SYNOPSYS_UNCONNECTED_57 ) , .Y ( SYNOPSYS_UNCONNECTED_58 ) ) ;
sky130_fd_sc_hd__inv_8 cts_inv_4667048875_4715349358 ( 
    .A ( SYNOPSYS_UNCONNECTED_59 ) , .Y ( SYNOPSYS_UNCONNECTED_60 ) ) ;
sky130_fd_sc_hd__inv_8 cts_inv_4669848903_4715449359 ( 
    .A ( SYNOPSYS_UNCONNECTED_61 ) , .Y ( SYNOPSYS_UNCONNECTED_62 ) ) ;
sky130_fd_sc_hd__inv_8 cts_inv_4700749212_4715549360 ( 
    .A ( SYNOPSYS_UNCONNECTED_63 ) , .Y ( SYNOPSYS_UNCONNECTED_64 ) ) ;
sky130_fd_sc_hd__inv_8 cts_inv_4700049205_4715649361 ( 
    .A ( SYNOPSYS_UNCONNECTED_65 ) , .Y ( SYNOPSYS_UNCONNECTED_66 ) ) ;
sky130_fd_sc_hd__inv_8 cts_inv_4695849163_4715749362 ( 
    .A ( SYNOPSYS_UNCONNECTED_67 ) , .Y ( SYNOPSYS_UNCONNECTED_68 ) ) ;
sky130_fd_sc_hd__clkinv_16 cts_inv_4684949054_4715849363 ( 
    .A ( SYNOPSYS_UNCONNECTED_69 ) , .Y ( SYNOPSYS_UNCONNECTED_70 ) ) ;
sky130_fd_sc_hd__inv_8 cts_inv_4680149006_4715949364 ( 
    .A ( SYNOPSYS_UNCONNECTED_71 ) , .Y ( SYNOPSYS_UNCONNECTED_72 ) ) ;
sky130_fd_sc_hd__inv_12 cts_inv_4680349008_4716149366 ( 
    .A ( SYNOPSYS_UNCONNECTED_73 ) , .Y ( p_abuf11 ) ) ;
sky130_fd_sc_hd__inv_12 cts_inv_4694549150_4716249367 ( 
    .A ( SYNOPSYS_UNCONNECTED_74 ) , .Y ( SYNOPSYS_UNCONNECTED_75 ) ) ;
sky130_fd_sc_hd__inv_8 cts_inv_4696549170_4716349368 ( 
    .A ( SYNOPSYS_UNCONNECTED_76 ) , .Y ( SYNOPSYS_UNCONNECTED_77 ) ) ;
sky130_fd_sc_hd__inv_8 cts_inv_4695949164_4716449369 ( 
    .A ( SYNOPSYS_UNCONNECTED_78 ) , .Y ( SYNOPSYS_UNCONNECTED_79 ) ) ;
sky130_fd_sc_hd__inv_8 cts_inv_4698049185_4716549370 ( 
    .A ( SYNOPSYS_UNCONNECTED_80 ) , .Y ( SYNOPSYS_UNCONNECTED_81 ) ) ;
sky130_fd_sc_hd__inv_8 cts_inv_4697249177_4716649371 ( 
    .A ( SYNOPSYS_UNCONNECTED_82 ) , .Y ( SYNOPSYS_UNCONNECTED_83 ) ) ;
sky130_fd_sc_hd__inv_8 cts_inv_4670148906_4716749372 ( 
    .A ( SYNOPSYS_UNCONNECTED_84 ) , .Y ( SYNOPSYS_UNCONNECTED_85 ) ) ;
sky130_fd_sc_hd__inv_8 cts_inv_4666248867_4716849373 ( 
    .A ( SYNOPSYS_UNCONNECTED_86 ) , .Y ( SYNOPSYS_UNCONNECTED_87 ) ) ;
sky130_fd_sc_hd__inv_8 cts_inv_4673648941_4716949374 ( 
    .A ( SYNOPSYS_UNCONNECTED_88 ) , .Y ( SYNOPSYS_UNCONNECTED_89 ) ) ;
sky130_fd_sc_hd__clkinv_16 cts_inv_4673548940_4717049375 ( 
    .A ( SYNOPSYS_UNCONNECTED_90 ) , .Y ( p_abuf8 ) ) ;
sky130_fd_sc_hd__inv_8 cts_inv_4675448959_4717149376 ( 
    .A ( SYNOPSYS_UNCONNECTED_91 ) , .Y ( SYNOPSYS_UNCONNECTED_92 ) ) ;
sky130_fd_sc_hd__inv_8 cts_inv_4667348878_4717249377 ( 
    .A ( SYNOPSYS_UNCONNECTED_93 ) , .Y ( p_abuf5 ) ) ;
sky130_fd_sc_hd__inv_16 cts_inv_4675248957_4717349378 ( 
    .A ( SYNOPSYS_UNCONNECTED_94 ) , .Y ( SYNOPSYS_UNCONNECTED_95 ) ) ;
sky130_fd_sc_hd__clkinv_8 cts_inv_4670748912_4717449379 ( 
    .A ( SYNOPSYS_UNCONNECTED_96 ) , .Y ( p_abuf3 ) ) ;
sky130_fd_sc_hd__inv_16 cts_inv_4710249307_4717549380 ( 
    .A ( SYNOPSYS_UNCONNECTED_97 ) , .Y ( SYNOPSYS_UNCONNECTED_98 ) ) ;
sky130_fd_sc_hd__inv_12 cts_inv_4705149256_4717649381 ( 
    .A ( SYNOPSYS_UNCONNECTED_99 ) , .Y ( SYNOPSYS_UNCONNECTED_100 ) ) ;
sky130_fd_sc_hd__inv_8 cts_inv_4705249257_4717749382 ( 
    .A ( SYNOPSYS_UNCONNECTED_101 ) , .Y ( SYNOPSYS_UNCONNECTED_102 ) ) ;
sky130_fd_sc_hd__inv_8 cts_inv_4708149286_4717849383 ( 
    .A ( SYNOPSYS_UNCONNECTED_103 ) , .Y ( SYNOPSYS_UNCONNECTED_104 ) ) ;
sky130_fd_sc_hd__inv_8 cts_inv_4705449259_4717949384 ( 
    .A ( SYNOPSYS_UNCONNECTED_105 ) , .Y ( SYNOPSYS_UNCONNECTED_106 ) ) ;
sky130_fd_sc_hd__inv_8 cts_inv_4705349258_4718049385 ( 
    .A ( SYNOPSYS_UNCONNECTED_107 ) , .Y ( SYNOPSYS_UNCONNECTED_108 ) ) ;
sky130_fd_sc_hd__inv_8 cts_inv_4683949044_4718149386 ( 
    .A ( SYNOPSYS_UNCONNECTED_109 ) , .Y ( SYNOPSYS_UNCONNECTED_110 ) ) ;
sky130_fd_sc_hd__inv_8 cts_inv_4682949034_4718249387 ( 
    .A ( SYNOPSYS_UNCONNECTED_111 ) , .Y ( SYNOPSYS_UNCONNECTED_112 ) ) ;
sky130_fd_sc_hd__inv_8 cts_inv_4703949244_4718349388 ( 
    .A ( SYNOPSYS_UNCONNECTED_113 ) , .Y ( SYNOPSYS_UNCONNECTED_114 ) ) ;
sky130_fd_sc_hd__inv_8 cts_inv_4700149206_4718449389 ( 
    .A ( SYNOPSYS_UNCONNECTED_115 ) , .Y ( SYNOPSYS_UNCONNECTED_116 ) ) ;
sky130_fd_sc_hd__inv_8 cts_inv_4702149226_4718549390 ( 
    .A ( SYNOPSYS_UNCONNECTED_117 ) , .Y ( SYNOPSYS_UNCONNECTED_118 ) ) ;
sky130_fd_sc_hd__inv_8 cts_inv_4679749002_4718649391 ( 
    .A ( SYNOPSYS_UNCONNECTED_119 ) , .Y ( SYNOPSYS_UNCONNECTED_120 ) ) ;
sky130_fd_sc_hd__inv_8 cts_inv_4675148956_4718749392 ( 
    .A ( SYNOPSYS_UNCONNECTED_121 ) , .Y ( p_abuf9 ) ) ;
sky130_fd_sc_hd__inv_8 cts_inv_4675948964_4718849393 ( 
    .A ( SYNOPSYS_UNCONNECTED_122 ) , .Y ( SYNOPSYS_UNCONNECTED_123 ) ) ;
sky130_fd_sc_hd__inv_8 cts_inv_4667748882_4718949394 ( 
    .A ( SYNOPSYS_UNCONNECTED_124 ) , .Y ( SYNOPSYS_UNCONNECTED_125 ) ) ;
sky130_fd_sc_hd__inv_8 cts_inv_4671348918_4719049395 ( 
    .A ( SYNOPSYS_UNCONNECTED_126 ) , .Y ( SYNOPSYS_UNCONNECTED_127 ) ) ;
sky130_fd_sc_hd__inv_8 cts_inv_4671448919_4719149396 ( 
    .A ( SYNOPSYS_UNCONNECTED_128 ) , .Y ( SYNOPSYS_UNCONNECTED_129 ) ) ;
sky130_fd_sc_hd__inv_8 cts_inv_4710049305_4719249397 ( 
    .A ( SYNOPSYS_UNCONNECTED_130 ) , .Y ( SYNOPSYS_UNCONNECTED_131 ) ) ;
sky130_fd_sc_hd__inv_8 cts_inv_4710349308_4719349398 ( 
    .A ( SYNOPSYS_UNCONNECTED_132 ) , .Y ( SYNOPSYS_UNCONNECTED_133 ) ) ;
sky130_fd_sc_hd__inv_6 cts_inv_4708349288_4719449399 ( 
    .A ( SYNOPSYS_UNCONNECTED_134 ) , .Y ( SYNOPSYS_UNCONNECTED_135 ) ) ;
sky130_fd_sc_hd__inv_8 cts_inv_4691649121_4719549400 ( 
    .A ( SYNOPSYS_UNCONNECTED_136 ) , .Y ( SYNOPSYS_UNCONNECTED_137 ) ) ;
sky130_fd_sc_hd__inv_16 cts_inv_4687249077_4719649401 ( 
    .A ( SYNOPSYS_UNCONNECTED_138 ) , .Y ( SYNOPSYS_UNCONNECTED_139 ) ) ;
sky130_fd_sc_hd__inv_8 cts_inv_4679649001_4719749402 ( 
    .A ( SYNOPSYS_UNCONNECTED_140 ) , .Y ( SYNOPSYS_UNCONNECTED_141 ) ) ;
sky130_fd_sc_hd__inv_12 cts_inv_4683549040_4719849403 ( 
    .A ( SYNOPSYS_UNCONNECTED_142 ) , .Y ( SYNOPSYS_UNCONNECTED_143 ) ) ;
sky130_fd_sc_hd__inv_8 cts_inv_4682749032_4719949404 ( 
    .A ( SYNOPSYS_UNCONNECTED_144 ) , .Y ( SYNOPSYS_UNCONNECTED_145 ) ) ;
sky130_fd_sc_hd__inv_8 cts_inv_4687449079_4720049405 ( 
    .A ( SYNOPSYS_UNCONNECTED_146 ) , .Y ( SYNOPSYS_UNCONNECTED_147 ) ) ;
sky130_fd_sc_hd__inv_12 cts_inv_4690649111_4720149406 ( 
    .A ( SYNOPSYS_UNCONNECTED_148 ) , .Y ( SYNOPSYS_UNCONNECTED_149 ) ) ;
sky130_fd_sc_hd__inv_8 cts_inv_4688349088_4720249407 ( 
    .A ( SYNOPSYS_UNCONNECTED_150 ) , .Y ( SYNOPSYS_UNCONNECTED_151 ) ) ;
sky130_fd_sc_hd__inv_8 cts_inv_4689349098_4720349408 ( 
    .A ( SYNOPSYS_UNCONNECTED_152 ) , .Y ( SYNOPSYS_UNCONNECTED_153 ) ) ;
sky130_fd_sc_hd__inv_8 cts_inv_4693749142_4720449409 ( 
    .A ( SYNOPSYS_UNCONNECTED_154 ) , .Y ( SYNOPSYS_UNCONNECTED_155 ) ) ;
sky130_fd_sc_hd__inv_6 cts_inv_4687549080_4720549410 ( 
    .A ( SYNOPSYS_UNCONNECTED_156 ) , .Y ( SYNOPSYS_UNCONNECTED_157 ) ) ;
sky130_fd_sc_hd__inv_8 cts_inv_4707449279_4720649411 ( 
    .A ( SYNOPSYS_UNCONNECTED_158 ) , .Y ( SYNOPSYS_UNCONNECTED_159 ) ) ;
sky130_fd_sc_hd__inv_8 cts_inv_4706949274_4720749412 ( 
    .A ( SYNOPSYS_UNCONNECTED_160 ) , .Y ( SYNOPSYS_UNCONNECTED_161 ) ) ;
sky130_fd_sc_hd__inv_8 cts_inv_4707049275_4720849413 ( 
    .A ( SYNOPSYS_UNCONNECTED_162 ) , .Y ( SYNOPSYS_UNCONNECTED_163 ) ) ;
sky130_fd_sc_hd__inv_16 cts_inv_4671048915_4721049415 ( 
    .A ( SYNOPSYS_UNCONNECTED_164 ) , .Y ( p_abuf4 ) ) ;
sky130_fd_sc_hd__inv_6 cts_inv_4670848913_4721149416 ( 
    .A ( SYNOPSYS_UNCONNECTED_165 ) , .Y ( SYNOPSYS_UNCONNECTED_166 ) ) ;
sky130_fd_sc_hd__inv_8 cts_inv_4667448879_4721249417 ( 
    .A ( SYNOPSYS_UNCONNECTED_167 ) , .Y ( SYNOPSYS_UNCONNECTED_168 ) ) ;
sky130_fd_sc_hd__inv_8 cts_inv_4667248877_4721349418 ( 
    .A ( SYNOPSYS_UNCONNECTED_169 ) , .Y ( SYNOPSYS_UNCONNECTED_170 ) ) ;
sky130_fd_sc_hd__inv_16 cts_inv_4695049155_4721449419 ( 
    .A ( SYNOPSYS_UNCONNECTED_171 ) , .Y ( SYNOPSYS_UNCONNECTED_172 ) ) ;
sky130_fd_sc_hd__inv_8 cts_inv_4693049135_4721549420 ( 
    .A ( SYNOPSYS_UNCONNECTED_173 ) , .Y ( SYNOPSYS_UNCONNECTED_174 ) ) ;
sky130_fd_sc_hd__inv_8 cts_inv_4692949134_4721649421 ( 
    .A ( SYNOPSYS_UNCONNECTED_175 ) , .Y ( SYNOPSYS_UNCONNECTED_176 ) ) ;
sky130_fd_sc_hd__inv_8 cts_inv_4693149136_4721749422 ( 
    .A ( SYNOPSYS_UNCONNECTED_177 ) , .Y ( SYNOPSYS_UNCONNECTED_178 ) ) ;
sky130_fd_sc_hd__inv_8 cts_inv_4701749222_4721849423 ( 
    .A ( SYNOPSYS_UNCONNECTED_179 ) , .Y ( SYNOPSYS_UNCONNECTED_180 ) ) ;
sky130_fd_sc_hd__inv_12 cts_inv_4706349268_4721949424 ( 
    .A ( SYNOPSYS_UNCONNECTED_181 ) , .Y ( SYNOPSYS_UNCONNECTED_182 ) ) ;
sky130_fd_sc_hd__inv_8 cts_inv_4704649251_4722049425 ( 
    .A ( SYNOPSYS_UNCONNECTED_183 ) , .Y ( SYNOPSYS_UNCONNECTED_184 ) ) ;
sky130_fd_sc_hd__inv_8 cts_inv_4709549300_4722149426 ( 
    .A ( SYNOPSYS_UNCONNECTED_185 ) , .Y ( SYNOPSYS_UNCONNECTED_186 ) ) ;
sky130_fd_sc_hd__clkinv_8 cts_inv_4707149276_4722249427 ( 
    .A ( SYNOPSYS_UNCONNECTED_187 ) , .Y ( SYNOPSYS_UNCONNECTED_188 ) ) ;
sky130_fd_sc_hd__inv_16 cts_inv_4704149246_4722349428 ( 
    .A ( SYNOPSYS_UNCONNECTED_189 ) , .Y ( SYNOPSYS_UNCONNECTED_190 ) ) ;
sky130_fd_sc_hd__inv_8 cts_inv_4674548950_4722449429 ( 
    .A ( SYNOPSYS_UNCONNECTED_191 ) , .Y ( SYNOPSYS_UNCONNECTED_192 ) ) ;
sky130_fd_sc_hd__inv_8 cts_inv_4679148996_4722549430 ( 
    .A ( SYNOPSYS_UNCONNECTED_193 ) , .Y ( SYNOPSYS_UNCONNECTED_194 ) ) ;
sky130_fd_sc_hd__inv_16 cts_inv_4678348988_4722649431 ( 
    .A ( SYNOPSYS_UNCONNECTED_195 ) , .Y ( SYNOPSYS_UNCONNECTED_196 ) ) ;
sky130_fd_sc_hd__inv_8 cts_inv_4678448989_4722749432 ( 
    .A ( SYNOPSYS_UNCONNECTED_197 ) , .Y ( SYNOPSYS_UNCONNECTED_198 ) ) ;
sky130_fd_sc_hd__inv_8 cts_inv_4674748952_4722849433 ( 
    .A ( SYNOPSYS_UNCONNECTED_199 ) , .Y ( SYNOPSYS_UNCONNECTED_200 ) ) ;
sky130_fd_sc_hd__inv_8 cts_inv_4673948944_4722949434 ( 
    .A ( SYNOPSYS_UNCONNECTED_201 ) , .Y ( SYNOPSYS_UNCONNECTED_202 ) ) ;
sky130_fd_sc_hd__inv_8 cts_inv_4673848943_4723049435 ( 
    .A ( SYNOPSYS_UNCONNECTED_203 ) , .Y ( SYNOPSYS_UNCONNECTED_204 ) ) ;
sky130_fd_sc_hd__inv_12 cts_inv_4709049295_4723149436 ( 
    .A ( SYNOPSYS_UNCONNECTED_205 ) , .Y ( SYNOPSYS_UNCONNECTED_206 ) ) ;
sky130_fd_sc_hd__inv_8 cts_inv_4707649281_4723249437 ( 
    .A ( SYNOPSYS_UNCONNECTED_207 ) , .Y ( SYNOPSYS_UNCONNECTED_208 ) ) ;
sky130_fd_sc_hd__inv_8 cts_inv_4708249287_4723349438 ( 
    .A ( SYNOPSYS_UNCONNECTED_209 ) , .Y ( SYNOPSYS_UNCONNECTED_210 ) ) ;
sky130_fd_sc_hd__inv_8 cts_inv_4692449129_4723449439 ( 
    .A ( SYNOPSYS_UNCONNECTED_211 ) , .Y ( SYNOPSYS_UNCONNECTED_212 ) ) ;
sky130_fd_sc_hd__inv_8 cts_inv_4687349078_4723549440 ( 
    .A ( SYNOPSYS_UNCONNECTED_213 ) , .Y ( SYNOPSYS_UNCONNECTED_214 ) ) ;
sky130_fd_sc_hd__clkinv_16 cts_inv_4677648981_4723649441 ( 
    .A ( SYNOPSYS_UNCONNECTED_215 ) , .Y ( SYNOPSYS_UNCONNECTED_216 ) ) ;
sky130_fd_sc_hd__clkinv_16 cts_inv_4684749052_4723749442 ( 
    .A ( SYNOPSYS_UNCONNECTED_217 ) , .Y ( SYNOPSYS_UNCONNECTED_218 ) ) ;
sky130_fd_sc_hd__clkinv_16 cts_inv_4684549050_4723849443 ( 
    .A ( SYNOPSYS_UNCONNECTED_219 ) , .Y ( SYNOPSYS_UNCONNECTED_220 ) ) ;
sky130_fd_sc_hd__inv_8 cts_inv_4675548960_4723949444 ( 
    .A ( SYNOPSYS_UNCONNECTED_221 ) , .Y ( SYNOPSYS_UNCONNECTED_222 ) ) ;
sky130_fd_sc_hd__inv_16 cts_inv_4682349028_4724049445 ( 
    .A ( SYNOPSYS_UNCONNECTED_223 ) , .Y ( SYNOPSYS_UNCONNECTED_224 ) ) ;
sky130_fd_sc_hd__inv_8 cts_inv_4680449009_4724149446 ( 
    .A ( SYNOPSYS_UNCONNECTED_225 ) , .Y ( SYNOPSYS_UNCONNECTED_226 ) ) ;
sky130_fd_sc_hd__inv_8 cts_inv_4680249007_4724249447 ( 
    .A ( SYNOPSYS_UNCONNECTED_227 ) , .Y ( SYNOPSYS_UNCONNECTED_228 ) ) ;
sky130_fd_sc_hd__inv_8 cts_inv_4685049055_4724349448 ( 
    .A ( SYNOPSYS_UNCONNECTED_229 ) , .Y ( SYNOPSYS_UNCONNECTED_230 ) ) ;
sky130_fd_sc_hd__clkinv_16 cts_inv_4686849073_4724449449 ( 
    .A ( SYNOPSYS_UNCONNECTED_231 ) , .Y ( p_abuf15 ) ) ;
sky130_fd_sc_hd__inv_8 cts_inv_4680049005_4724549450 ( 
    .A ( SYNOPSYS_UNCONNECTED_232 ) , .Y ( SYNOPSYS_UNCONNECTED_233 ) ) ;
sky130_fd_sc_hd__clkinv_16 cts_inv_4689449099_4724649451 ( 
    .A ( SYNOPSYS_UNCONNECTED_234 ) , .Y ( SYNOPSYS_UNCONNECTED_235 ) ) ;
sky130_fd_sc_hd__inv_16 cts_inv_4692749132_4724749452 ( 
    .A ( SYNOPSYS_UNCONNECTED_236 ) , .Y ( SYNOPSYS_UNCONNECTED_237 ) ) ;
sky130_fd_sc_hd__inv_16 cts_inv_4693649141_4724849453 ( 
    .A ( SYNOPSYS_UNCONNECTED_238 ) , .Y ( SYNOPSYS_UNCONNECTED_239 ) ) ;
sky130_fd_sc_hd__inv_8 cts_inv_4677148976_4724949454 ( 
    .A ( SYNOPSYS_UNCONNECTED_240 ) , .Y ( SYNOPSYS_UNCONNECTED_241 ) ) ;
sky130_fd_sc_hd__inv_8 cts_inv_4670448909_4725049455 ( 
    .A ( SYNOPSYS_UNCONNECTED_242 ) , .Y ( SYNOPSYS_UNCONNECTED_243 ) ) ;
sky130_fd_sc_hd__inv_12 cts_inv_4679549000_4725149456 ( 
    .A ( SYNOPSYS_UNCONNECTED_244 ) , .Y ( SYNOPSYS_UNCONNECTED_245 ) ) ;
sky130_fd_sc_hd__clkinv_8 cts_inv_4679348998_4725249457 ( 
    .A ( SYNOPSYS_UNCONNECTED_246 ) , .Y ( SYNOPSYS_UNCONNECTED_247 ) ) ;
sky130_fd_sc_hd__inv_12 cts_inv_4678548990_4725349458 ( 
    .A ( SYNOPSYS_UNCONNECTED_248 ) , .Y ( SYNOPSYS_UNCONNECTED_249 ) ) ;
sky130_fd_sc_hd__inv_8 cts_inv_4708949294_4725449459 ( 
    .A ( SYNOPSYS_UNCONNECTED_250 ) , .Y ( SYNOPSYS_UNCONNECTED_251 ) ) ;
sky130_fd_sc_hd__inv_8 cts_inv_4709849303_4725549460 ( 
    .A ( SYNOPSYS_UNCONNECTED_252 ) , .Y ( SYNOPSYS_UNCONNECTED_253 ) ) ;
sky130_fd_sc_hd__inv_8 cts_inv_4704049245_4725649461 ( 
    .A ( SYNOPSYS_UNCONNECTED_254 ) , .Y ( SYNOPSYS_UNCONNECTED_255 ) ) ;
sky130_fd_sc_hd__inv_8 cts_inv_4685849063_4725749462 ( 
    .A ( SYNOPSYS_UNCONNECTED_256 ) , .Y ( SYNOPSYS_UNCONNECTED_257 ) ) ;
sky130_fd_sc_hd__inv_12 cts_inv_4691549120_4725849463 ( 
    .A ( SYNOPSYS_UNCONNECTED_258 ) , .Y ( SYNOPSYS_UNCONNECTED_259 ) ) ;
sky130_fd_sc_hd__inv_8 cts_inv_4687849083_4725949464 ( 
    .A ( SYNOPSYS_UNCONNECTED_260 ) , .Y ( SYNOPSYS_UNCONNECTED_261 ) ) ;
sky130_fd_sc_hd__inv_12 cts_inv_4682649031_4726049465 ( 
    .A ( SYNOPSYS_UNCONNECTED_262 ) , .Y ( SYNOPSYS_UNCONNECTED_263 ) ) ;
sky130_fd_sc_hd__inv_16 cts_inv_4681549020_4726149466 ( 
    .A ( SYNOPSYS_UNCONNECTED_264 ) , .Y ( SYNOPSYS_UNCONNECTED_265 ) ) ;
sky130_fd_sc_hd__inv_8 cts_inv_4686049065_4726249467 ( 
    .A ( SYNOPSYS_UNCONNECTED_266 ) , .Y ( SYNOPSYS_UNCONNECTED_267 ) ) ;
sky130_fd_sc_hd__inv_8 cts_inv_4682849033_4726349468 ( 
    .A ( SYNOPSYS_UNCONNECTED_268 ) , .Y ( SYNOPSYS_UNCONNECTED_269 ) ) ;
sky130_fd_sc_hd__inv_8 cts_inv_4688149086_4726449469 ( 
    .A ( SYNOPSYS_UNCONNECTED_270 ) , .Y ( SYNOPSYS_UNCONNECTED_271 ) ) ;
sky130_fd_sc_hd__inv_16 cts_inv_4665848863_4726549470 ( 
    .A ( SYNOPSYS_UNCONNECTED_272 ) , .Y ( SYNOPSYS_UNCONNECTED_273 ) ) ;
sky130_fd_sc_hd__inv_16 cts_inv_4698949194_4726649471 ( 
    .A ( SYNOPSYS_UNCONNECTED_274 ) , .Y ( SYNOPSYS_UNCONNECTED_275 ) ) ;
sky130_fd_sc_hd__inv_8 cts_inv_4691449119_4726749472 ( 
    .A ( SYNOPSYS_UNCONNECTED_276 ) , .Y ( SYNOPSYS_UNCONNECTED_277 ) ) ;
sky130_fd_sc_hd__inv_16 cts_inv_4686649071_4726849473 ( 
    .A ( SYNOPSYS_UNCONNECTED_278 ) , .Y ( SYNOPSYS_UNCONNECTED_279 ) ) ;
sky130_fd_sc_hd__clkinv_16 cts_inv_4693349138_4726949474 ( 
    .A ( SYNOPSYS_UNCONNECTED_280 ) , .Y ( p_abuf17 ) ) ;
sky130_fd_sc_hd__inv_16 cts_inv_4672448929_4727049475 ( 
    .A ( SYNOPSYS_UNCONNECTED_281 ) , .Y ( SYNOPSYS_UNCONNECTED_282 ) ) ;
sky130_fd_sc_hd__inv_16 cts_inv_4668548890_4727149476 ( 
    .A ( SYNOPSYS_UNCONNECTED_283 ) , .Y ( SYNOPSYS_UNCONNECTED_284 ) ) ;
sky130_fd_sc_hd__inv_16 cts_inv_4681649021_4727249477 ( 
    .A ( SYNOPSYS_UNCONNECTED_285 ) , .Y ( SYNOPSYS_UNCONNECTED_286 ) ) ;
sky130_fd_sc_hd__clkinv_16 cts_inv_4672648931_4727349478 ( 
    .A ( SYNOPSYS_UNCONNECTED_287 ) , .Y ( SYNOPSYS_UNCONNECTED_288 ) ) ;
sky130_fd_sc_hd__clkinv_16 cts_inv_4681749022_4727449479 ( 
    .A ( SYNOPSYS_UNCONNECTED_289 ) , .Y ( SYNOPSYS_UNCONNECTED_290 ) ) ;
sky130_fd_sc_hd__inv_12 cts_inv_4672748932_4727549480 ( 
    .A ( SYNOPSYS_UNCONNECTED_291 ) , .Y ( SYNOPSYS_UNCONNECTED_292 ) ) ;
sky130_fd_sc_hd__clkinv_16 cts_inv_4683749042_4727649481 ( 
    .A ( SYNOPSYS_UNCONNECTED_293 ) , .Y ( SYNOPSYS_UNCONNECTED_294 ) ) ;
sky130_fd_sc_hd__inv_12 cts_inv_4680549010_4727749482 ( 
    .A ( SYNOPSYS_UNCONNECTED_295 ) , .Y ( SYNOPSYS_UNCONNECTED_296 ) ) ;
sky130_fd_sc_hd__inv_8 cts_inv_4695549160_4727849483 ( 
    .A ( SYNOPSYS_UNCONNECTED_297 ) , .Y ( SYNOPSYS_UNCONNECTED_298 ) ) ;
sky130_fd_sc_hd__inv_16 cts_inv_4699349198_4727949484 ( 
    .A ( SYNOPSYS_UNCONNECTED_299 ) , .Y ( SYNOPSYS_UNCONNECTED_300 ) ) ;
sky130_fd_sc_hd__inv_16 cts_inv_4699949204_4728049485 ( 
    .A ( SYNOPSYS_UNCONNECTED_301 ) , .Y ( SYNOPSYS_UNCONNECTED_302 ) ) ;
sky130_fd_sc_hd__inv_8 cts_inv_4697049175_4728149486 ( 
    .A ( SYNOPSYS_UNCONNECTED_303 ) , .Y ( SYNOPSYS_UNCONNECTED_304 ) ) ;
sky130_fd_sc_hd__inv_8 cts_inv_4700449209_4728249487 ( 
    .A ( SYNOPSYS_UNCONNECTED_305 ) , .Y ( SYNOPSYS_UNCONNECTED_306 ) ) ;
sky130_fd_sc_hd__inv_8 cts_inv_4673148936_4728349488 ( 
    .A ( SYNOPSYS_UNCONNECTED_307 ) , .Y ( p_abuf7 ) ) ;
sky130_fd_sc_hd__inv_16 cts_inv_4669148896_4728449489 ( 
    .A ( SYNOPSYS_UNCONNECTED_308 ) , .Y ( SYNOPSYS_UNCONNECTED_309 ) ) ;
sky130_fd_sc_hd__inv_8 cts_inv_4671148916_4728649491 ( 
    .A ( SYNOPSYS_UNCONNECTED_310 ) , .Y ( SYNOPSYS_UNCONNECTED_311 ) ) ;
sky130_fd_sc_hd__inv_8 cts_inv_4688649091_4728749492 ( 
    .A ( SYNOPSYS_UNCONNECTED_312 ) , .Y ( p_abuf12 ) ) ;
sky130_fd_sc_hd__inv_8 cts_inv_4691249117_4728849493 ( 
    .A ( SYNOPSYS_UNCONNECTED_313 ) , .Y ( SYNOPSYS_UNCONNECTED_314 ) ) ;
sky130_fd_sc_hd__clkinv_16 cts_inv_4701449219_4728949494 ( 
    .A ( SYNOPSYS_UNCONNECTED_315 ) , .Y ( p_abuf21 ) ) ;
sky130_fd_sc_hd__inv_12 cts_inv_4702249227_4729049495 ( 
    .A ( SYNOPSYS_UNCONNECTED_316 ) , .Y ( SYNOPSYS_UNCONNECTED_317 ) ) ;
sky130_fd_sc_hd__inv_8 cts_inv_4693549140_4729149496 ( 
    .A ( SYNOPSYS_UNCONNECTED_318 ) , .Y ( SYNOPSYS_UNCONNECTED_319 ) ) ;
sky130_fd_sc_hd__inv_8 cts_inv_4677848983_4729249497 ( 
    .A ( SYNOPSYS_UNCONNECTED_320 ) , .Y ( SYNOPSYS_UNCONNECTED_321 ) ) ;
sky130_fd_sc_hd__inv_16 cts_inv_4673348938_4729349498 ( 
    .A ( SYNOPSYS_UNCONNECTED_322 ) , .Y ( SYNOPSYS_UNCONNECTED_323 ) ) ;
sky130_fd_sc_hd__inv_16 cts_inv_4677248977_4729449499 ( 
    .A ( SYNOPSYS_UNCONNECTED_324 ) , .Y ( SYNOPSYS_UNCONNECTED_325 ) ) ;
sky130_fd_sc_hd__inv_16 cts_inv_4671548920_4729549500 ( 
    .A ( SYNOPSYS_UNCONNECTED_326 ) , .Y ( SYNOPSYS_UNCONNECTED_327 ) ) ;
sky130_fd_sc_hd__inv_16 cts_inv_4709349298_4729649501 ( 
    .A ( SYNOPSYS_UNCONNECTED_328 ) , .Y ( SYNOPSYS_UNCONNECTED_329 ) ) ;
sky130_fd_sc_hd__inv_8 cts_inv_4711449319_4729749502 ( 
    .A ( SYNOPSYS_UNCONNECTED_330 ) , .Y ( SYNOPSYS_UNCONNECTED_331 ) ) ;
sky130_fd_sc_hd__inv_16 cts_inv_4703149236_4729849503 ( 
    .A ( SYNOPSYS_UNCONNECTED_332 ) , .Y ( SYNOPSYS_UNCONNECTED_333 ) ) ;
sky130_fd_sc_hd__clkinv_16 cts_inv_4692149126_4729949504 ( 
    .A ( SYNOPSYS_UNCONNECTED_334 ) , .Y ( p_abuf18 ) ) ;
sky130_fd_sc_hd__clkinv_16 cts_inv_4696049165_4730049505 ( 
    .A ( SYNOPSYS_UNCONNECTED_335 ) , .Y ( SYNOPSYS_UNCONNECTED_336 ) ) ;
sky130_fd_sc_hd__inv_16 cts_inv_4686349068_4730149506 ( 
    .A ( SYNOPSYS_UNCONNECTED_337 ) , .Y ( SYNOPSYS_UNCONNECTED_338 ) ) ;
sky130_fd_sc_hd__clkinv_16 cts_inv_4697549180_4730249507 ( 
    .A ( SYNOPSYS_UNCONNECTED_339 ) , .Y ( SYNOPSYS_UNCONNECTED_340 ) ) ;
sky130_fd_sc_hd__inv_8 cts_inv_4684149046_4730349508 ( 
    .A ( SYNOPSYS_UNCONNECTED_341 ) , .Y ( SYNOPSYS_UNCONNECTED_342 ) ) ;
sky130_fd_sc_hd__inv_8 cts_inv_4672848933_4730449509 ( 
    .A ( SYNOPSYS_UNCONNECTED_343 ) , .Y ( SYNOPSYS_UNCONNECTED_344 ) ) ;
sky130_fd_sc_hd__inv_16 cts_inv_4683249037_4730549510 ( 
    .A ( SYNOPSYS_UNCONNECTED_345 ) , .Y ( SYNOPSYS_UNCONNECTED_346 ) ) ;
sky130_fd_sc_hd__clkinv_8 cts_inv_4691749122_4730649511 ( 
    .A ( SYNOPSYS_UNCONNECTED_347 ) , .Y ( SYNOPSYS_UNCONNECTED_348 ) ) ;
sky130_fd_sc_hd__inv_8 cts_inv_4678248987_4730749512 ( 
    .A ( SYNOPSYS_UNCONNECTED_349 ) , .Y ( SYNOPSYS_UNCONNECTED_350 ) ) ;
sky130_fd_sc_hd__inv_8 cts_inv_4703649241_4730849513 ( 
    .A ( SYNOPSYS_UNCONNECTED_351 ) , .Y ( SYNOPSYS_UNCONNECTED_352 ) ) ;
sky130_fd_sc_hd__inv_12 cts_inv_4697749182_4730949514 ( 
    .A ( SYNOPSYS_UNCONNECTED_353 ) , .Y ( SYNOPSYS_UNCONNECTED_354 ) ) ;
sky130_fd_sc_hd__clkinv_8 cts_inv_4702049225_4731049515 ( 
    .A ( SYNOPSYS_UNCONNECTED_355 ) , .Y ( SYNOPSYS_UNCONNECTED_356 ) ) ;
sky130_fd_sc_hd__inv_12 cts_inv_4681349018_4731149516 ( 
    .A ( SYNOPSYS_UNCONNECTED_357 ) , .Y ( SYNOPSYS_UNCONNECTED_358 ) ) ;
sky130_fd_sc_hd__inv_6 cts_inv_4690449109_4731249517 ( 
    .A ( SYNOPSYS_UNCONNECTED_359 ) , .Y ( p_abuf14 ) ) ;
sky130_fd_sc_hd__clkinv_16 cts_inv_4696149166_4731349518 ( 
    .A ( SYNOPSYS_UNCONNECTED_360 ) , .Y ( SYNOPSYS_UNCONNECTED_361 ) ) ;
sky130_fd_sc_hd__inv_8 cts_inv_4673048935_4731449519 ( 
    .A ( SYNOPSYS_UNCONNECTED_362 ) , .Y ( SYNOPSYS_UNCONNECTED_363 ) ) ;
sky130_fd_sc_hd__clkinv_16 cts_inv_4682149026_4731549520 ( 
    .A ( SYNOPSYS_UNCONNECTED_364 ) , .Y ( SYNOPSYS_UNCONNECTED_365 ) ) ;
sky130_fd_sc_hd__inv_16 cts_inv_4677348978_4731649521 ( 
    .A ( SYNOPSYS_UNCONNECTED_366 ) , .Y ( SYNOPSYS_UNCONNECTED_367 ) ) ;
sky130_fd_sc_hd__clkinv_16 cts_inv_4686149066_4731749522 ( 
    .A ( SYNOPSYS_UNCONNECTED_368 ) , .Y ( SYNOPSYS_UNCONNECTED_369 ) ) ;
sky130_fd_sc_hd__clkinv_16 cts_inv_4694949154_4731849523 ( 
    .A ( SYNOPSYS_UNCONNECTED_370 ) , .Y ( SYNOPSYS_UNCONNECTED_371 ) ) ;
sky130_fd_sc_hd__clkinv_8 cts_inv_4696249167_4731949524 ( 
    .A ( SYNOPSYS_UNCONNECTED_372 ) , .Y ( SYNOPSYS_UNCONNECTED_373 ) ) ;
sky130_fd_sc_hd__clkinv_16 cts_inv_4708849293_4732049525 ( 
    .A ( SYNOPSYS_UNCONNECTED_374 ) , .Y ( SYNOPSYS_UNCONNECTED_375 ) ) ;
sky130_fd_sc_hd__inv_8 cts_inv_4700249207_4732149526 ( 
    .A ( SYNOPSYS_UNCONNECTED_376 ) , .Y ( SYNOPSYS_UNCONNECTED_377 ) ) ;
sky130_fd_sc_hd__clkinv_16 cts_inv_4676848973_4732249527 ( 
    .A ( SYNOPSYS_UNCONNECTED_378 ) , .Y ( SYNOPSYS_UNCONNECTED_379 ) ) ;
sky130_fd_sc_hd__clkinv_16 cts_inv_4681849023_4732449529 ( 
    .A ( SYNOPSYS_UNCONNECTED_380 ) , .Y ( p_abuf13 ) ) ;
sky130_fd_sc_hd__clkinv_16 cts_inv_4690749112_4732549530 ( 
    .A ( SYNOPSYS_UNCONNECTED_381 ) , .Y ( SYNOPSYS_UNCONNECTED_382 ) ) ;
sky130_fd_sc_hd__clkinv_16 cts_inv_4694849153_4732749532 ( 
    .A ( SYNOPSYS_UNCONNECTED_383 ) , .Y ( SYNOPSYS_UNCONNECTED_384 ) ) ;
sky130_fd_sc_hd__clkinv_16 cts_inv_4694749152_4733049535 ( 
    .A ( SYNOPSYS_UNCONNECTED_385 ) , .Y ( SYNOPSYS_UNCONNECTED_386 ) ) ;
sky130_fd_sc_hd__inv_8 cts_inv_4690249107_4733349538 ( 
    .A ( SYNOPSYS_UNCONNECTED_387 ) , .Y ( SYNOPSYS_UNCONNECTED_388 ) ) ;
sky130_fd_sc_hd__inv_8 cts_inv_4701049215_4733549540 ( 
    .A ( SYNOPSYS_UNCONNECTED_389 ) , .Y ( SYNOPSYS_UNCONNECTED_390 ) ) ;
sky130_fd_sc_hd__clkinv_8 cts_inv_4697849183_4733749542 ( 
    .A ( SYNOPSYS_UNCONNECTED_391 ) , .Y ( SYNOPSYS_UNCONNECTED_392 ) ) ;
sky130_fd_sc_hd__inv_8 cts_inv_4693449139_4733849543 ( 
    .A ( SYNOPSYS_UNCONNECTED_393 ) , .Y ( SYNOPSYS_UNCONNECTED_394 ) ) ;
sky130_fd_sc_hd__inv_8 cts_inv_4697949184_4733949544 ( 
    .A ( SYNOPSYS_UNCONNECTED_395 ) , .Y ( SYNOPSYS_UNCONNECTED_396 ) ) ;
sky130_fd_sc_hd__inv_8 cts_inv_4689149096_4734149546 ( 
    .A ( SYNOPSYS_UNCONNECTED_397 ) , .Y ( SYNOPSYS_UNCONNECTED_398 ) ) ;
sky130_fd_sc_hd__inv_16 cts_inv_4688949094_4734249547 ( 
    .A ( SYNOPSYS_UNCONNECTED_399 ) , .Y ( SYNOPSYS_UNCONNECTED_400 ) ) ;
sky130_fd_sc_hd__inv_8 cts_inv_4696849173_4734749552 ( 
    .A ( SYNOPSYS_UNCONNECTED_401 ) , .Y ( SYNOPSYS_UNCONNECTED_402 ) ) ;
sky130_fd_sc_hd__clkinvlp_4 cts_inv_4845350658 ( .A ( ctsbuf_net_6532635 ) , 
    .Y ( ctsbuf_net_5822564 ) ) ;
sky130_fd_sc_hd__clkinvlp_4 cts_inv_4845450659 ( .A ( ctsbuf_net_6552637 ) , 
    .Y ( ctsbuf_net_5832565 ) ) ;
sky130_fd_sc_hd__clkinvlp_4 cts_inv_4845550660 ( .A ( ctsbuf_net_6452627 ) , 
    .Y ( ctsbuf_net_5842566 ) ) ;
sky130_fd_sc_hd__clkinvlp_4 cts_inv_4845650661 ( .A ( ctsbuf_net_6512633 ) , 
    .Y ( ctsbuf_net_5852567 ) ) ;
sky130_fd_sc_hd__clkinvlp_4 cts_inv_4845750662 ( .A ( ctsbuf_net_6492631 ) , 
    .Y ( ctsbuf_net_5862568 ) ) ;
sky130_fd_sc_hd__clkinvlp_2 cts_inv_4845850663 ( .A ( ctsbuf_net_6492631 ) , 
    .Y ( ctsbuf_net_5872569 ) ) ;
sky130_fd_sc_hd__clkinvlp_2 cts_inv_4845950664 ( .A ( ctsbuf_net_6492631 ) , 
    .Y ( ctsbuf_net_5882570 ) ) ;
sky130_fd_sc_hd__clkinvlp_2 cts_inv_4846050665 ( .A ( ctsbuf_net_6452627 ) , 
    .Y ( ctsbuf_net_5892571 ) ) ;
sky130_fd_sc_hd__clkinvlp_2 cts_inv_4846150666 ( .A ( ctsbuf_net_6512633 ) , 
    .Y ( ctsbuf_net_5902572 ) ) ;
sky130_fd_sc_hd__clkinvlp_2 cts_inv_4846250667 ( .A ( ctsbuf_net_6492631 ) , 
    .Y ( ctsbuf_net_5912573 ) ) ;
sky130_fd_sc_hd__clkinvlp_4 cts_inv_4846350668 ( .A ( ctsbuf_net_6562638 ) , 
    .Y ( ctsbuf_net_5922574 ) ) ;
sky130_fd_sc_hd__clkinvlp_4 cts_inv_4846450669 ( .A ( ctsbuf_net_6562638 ) , 
    .Y ( ctsbuf_net_5932575 ) ) ;
sky130_fd_sc_hd__clkinvlp_4 cts_inv_4846550670 ( .A ( ctsbuf_net_6492631 ) , 
    .Y ( ctsbuf_net_5942576 ) ) ;
sky130_fd_sc_hd__clkinvlp_2 cts_inv_4846650671 ( .A ( ctsbuf_net_6452627 ) , 
    .Y ( ctsbuf_net_5952577 ) ) ;
sky130_fd_sc_hd__clkinvlp_2 cts_inv_4846750672 ( .A ( ctsbuf_net_6552637 ) , 
    .Y ( ctsbuf_net_5962578 ) ) ;
sky130_fd_sc_hd__clkinvlp_4 cts_inv_4846850673 ( .A ( ctsbuf_net_6562638 ) , 
    .Y ( ctsbuf_net_5972579 ) ) ;
sky130_fd_sc_hd__clkinvlp_2 cts_inv_4846950674 ( .A ( ctsbuf_net_6482630 ) , 
    .Y ( ctsbuf_net_5982580 ) ) ;
sky130_fd_sc_hd__clkinvlp_2 cts_inv_4847050675 ( .A ( ctsbuf_net_6472629 ) , 
    .Y ( ctsbuf_net_5992581 ) ) ;
sky130_fd_sc_hd__clkinvlp_4 cts_inv_4847150676 ( .A ( ctsbuf_net_6482630 ) , 
    .Y ( ctsbuf_net_6002582 ) ) ;
sky130_fd_sc_hd__clkinvlp_2 cts_inv_4847250677 ( .A ( ctsbuf_net_6502632 ) , 
    .Y ( ctsbuf_net_6012583 ) ) ;
sky130_fd_sc_hd__clkinvlp_2 cts_inv_4847350678 ( .A ( ctsbuf_net_6512633 ) , 
    .Y ( ctsbuf_net_6022584 ) ) ;
sky130_fd_sc_hd__clkinvlp_2 cts_inv_4847450679 ( .A ( ctsbuf_net_6472629 ) , 
    .Y ( ctsbuf_net_6032585 ) ) ;
sky130_fd_sc_hd__clkinvlp_4 cts_inv_4847550680 ( .A ( ctsbuf_net_6532635 ) , 
    .Y ( ctsbuf_net_6042586 ) ) ;
sky130_fd_sc_hd__clkinvlp_4 cts_inv_4847650681 ( .A ( ctsbuf_net_6462628 ) , 
    .Y ( ctsbuf_net_6052587 ) ) ;
sky130_fd_sc_hd__clkinvlp_2 cts_inv_4847750682 ( .A ( ctsbuf_net_6532635 ) , 
    .Y ( ctsbuf_net_6062588 ) ) ;
sky130_fd_sc_hd__clkinvlp_4 cts_inv_4847850683 ( .A ( ctsbuf_net_6452627 ) , 
    .Y ( ctsbuf_net_6072589 ) ) ;
sky130_fd_sc_hd__clkinvlp_4 cts_inv_4847950684 ( .A ( ctsbuf_net_6452627 ) , 
    .Y ( ctsbuf_net_6082590 ) ) ;
sky130_fd_sc_hd__clkinvlp_2 cts_inv_4848050685 ( .A ( ctsbuf_net_6472629 ) , 
    .Y ( ctsbuf_net_6092591 ) ) ;
sky130_fd_sc_hd__clkinvlp_2 cts_inv_4848150686 ( .A ( ctsbuf_net_6532635 ) , 
    .Y ( ctsbuf_net_6102592 ) ) ;
sky130_fd_sc_hd__clkinvlp_4 cts_inv_4848250687 ( .A ( ctsbuf_net_6452627 ) , 
    .Y ( ctsbuf_net_6112593 ) ) ;
sky130_fd_sc_hd__clkinvlp_4 cts_inv_4848350688 ( .A ( ctsbuf_net_6452627 ) , 
    .Y ( ctsbuf_net_6122594 ) ) ;
sky130_fd_sc_hd__clkinvlp_4 cts_inv_4848450689 ( .A ( ctsbuf_net_6542636 ) , 
    .Y ( ctsbuf_net_6132595 ) ) ;
sky130_fd_sc_hd__clkinvlp_2 cts_inv_4848550690 ( .A ( ctsbuf_net_6552637 ) , 
    .Y ( ctsbuf_net_6142596 ) ) ;
sky130_fd_sc_hd__clkinvlp_4 cts_inv_4848650691 ( .A ( ctsbuf_net_6472629 ) , 
    .Y ( ctsbuf_net_6152597 ) ) ;
sky130_fd_sc_hd__clkinvlp_4 cts_inv_4848750692 ( .A ( ctsbuf_net_6552637 ) , 
    .Y ( ctsbuf_net_6162598 ) ) ;
sky130_fd_sc_hd__clkinvlp_4 cts_inv_4848850693 ( .A ( ctsbuf_net_6462628 ) , 
    .Y ( ctsbuf_net_6172599 ) ) ;
sky130_fd_sc_hd__clkinvlp_4 cts_inv_4848950694 ( .A ( ctsbuf_net_6572639 ) , 
    .Y ( ctsbuf_net_6182600 ) ) ;
sky130_fd_sc_hd__clkinvlp_2 cts_inv_4849050695 ( .A ( ctsbuf_net_6532635 ) , 
    .Y ( ctsbuf_net_6192601 ) ) ;
sky130_fd_sc_hd__clkinvlp_4 cts_inv_4849150696 ( .A ( ctsbuf_net_6482630 ) , 
    .Y ( ctsbuf_net_6202602 ) ) ;
sky130_fd_sc_hd__clkinvlp_2 cts_inv_4849250697 ( .A ( ctsbuf_net_6502632 ) , 
    .Y ( ctsbuf_net_6212603 ) ) ;
sky130_fd_sc_hd__inv_2 cts_inv_4849350698 ( .A ( ctsbuf_net_6502632 ) , 
    .Y ( ctsbuf_net_6222604 ) ) ;
sky130_fd_sc_hd__clkinvlp_2 cts_inv_4849450699 ( .A ( ctsbuf_net_6462628 ) , 
    .Y ( ctsbuf_net_6232605 ) ) ;
sky130_fd_sc_hd__clkinvlp_4 cts_inv_4849550700 ( .A ( ctsbuf_net_6462628 ) , 
    .Y ( ctsbuf_net_6242606 ) ) ;
sky130_fd_sc_hd__clkinvlp_4 cts_inv_4849650701 ( .A ( ctsbuf_net_6542636 ) , 
    .Y ( ctsbuf_net_6252607 ) ) ;
sky130_fd_sc_hd__clkinvlp_2 cts_inv_4849750702 ( .A ( ctsbuf_net_6512633 ) , 
    .Y ( ctsbuf_net_6262608 ) ) ;
sky130_fd_sc_hd__clkinvlp_2 cts_inv_4849850703 ( .A ( ctsbuf_net_6542636 ) , 
    .Y ( ctsbuf_net_6272609 ) ) ;
sky130_fd_sc_hd__clkinvlp_2 cts_inv_4849950704 ( .A ( ctsbuf_net_6542636 ) , 
    .Y ( ctsbuf_net_6282610 ) ) ;
sky130_fd_sc_hd__clkinvlp_2 cts_inv_4850050705 ( .A ( ctsbuf_net_6502632 ) , 
    .Y ( ctsbuf_net_6292611 ) ) ;
sky130_fd_sc_hd__clkinvlp_4 cts_inv_4850150706 ( .A ( ctsbuf_net_6572639 ) , 
    .Y ( ctsbuf_net_6302612 ) ) ;
sky130_fd_sc_hd__clkinvlp_2 cts_inv_4850250707 ( .A ( ctsbuf_net_6462628 ) , 
    .Y ( ctsbuf_net_6312613 ) ) ;
sky130_fd_sc_hd__clkinvlp_2 cts_inv_4850350708 ( .A ( ctsbuf_net_6462628 ) , 
    .Y ( ctsbuf_net_6322614 ) ) ;
sky130_fd_sc_hd__clkinvlp_2 cts_inv_4850450709 ( .A ( ctsbuf_net_6522634 ) , 
    .Y ( ctsbuf_net_6332615 ) ) ;
sky130_fd_sc_hd__clkinvlp_2 cts_inv_4850550710 ( .A ( ctsbuf_net_6522634 ) , 
    .Y ( ctsbuf_net_6342616 ) ) ;
sky130_fd_sc_hd__clkinvlp_2 cts_inv_4850650711 ( .A ( ctsbuf_net_6532635 ) , 
    .Y ( ctsbuf_net_6352617 ) ) ;
sky130_fd_sc_hd__clkinvlp_2 cts_inv_4850750712 ( .A ( ctsbuf_net_6482630 ) , 
    .Y ( ctsbuf_net_6362618 ) ) ;
sky130_fd_sc_hd__clkinvlp_2 cts_inv_4850850713 ( .A ( ctsbuf_net_6462628 ) , 
    .Y ( ctsbuf_net_6372619 ) ) ;
sky130_fd_sc_hd__clkinvlp_2 cts_inv_4850950714 ( .A ( ctsbuf_net_6482630 ) , 
    .Y ( ctsbuf_net_6382620 ) ) ;
sky130_fd_sc_hd__clkinvlp_2 cts_inv_4851050715 ( .A ( ctsbuf_net_6522634 ) , 
    .Y ( ctsbuf_net_6392621 ) ) ;
sky130_fd_sc_hd__clkinvlp_4 cts_inv_4851150716 ( .A ( ctsbuf_net_6522634 ) , 
    .Y ( ctsbuf_net_6402622 ) ) ;
sky130_fd_sc_hd__clkinvlp_2 cts_inv_4851250717 ( .A ( ctsbuf_net_6482630 ) , 
    .Y ( ctsbuf_net_6412623 ) ) ;
sky130_fd_sc_hd__clkinvlp_4 cts_inv_4851350718 ( .A ( ctsbuf_net_6542636 ) , 
    .Y ( ctsbuf_net_6422624 ) ) ;
sky130_fd_sc_hd__clkinvlp_2 cts_inv_4851450719 ( .A ( ctsbuf_net_6512633 ) , 
    .Y ( ctsbuf_net_6432625 ) ) ;
sky130_fd_sc_hd__clkinvlp_4 cts_inv_4851550720 ( .A ( ctsbuf_net_6502632 ) , 
    .Y ( ctsbuf_net_6442626 ) ) ;
sky130_fd_sc_hd__clkinvlp_4 cts_inv_4858650791 ( .A ( ctsbuf_net_6592641 ) , 
    .Y ( ctsbuf_net_6452627 ) ) ;
sky130_fd_sc_hd__clkinv_1 cts_inv_4858750792 ( .A ( ctsbuf_net_6582640 ) , 
    .Y ( ctsbuf_net_6462628 ) ) ;
sky130_fd_sc_hd__clkinvlp_4 cts_inv_4858850793 ( .A ( ctsbuf_net_6592641 ) , 
    .Y ( ctsbuf_net_6472629 ) ) ;
sky130_fd_sc_hd__clkinv_1 cts_inv_4858950794 ( .A ( ctsbuf_net_6582640 ) , 
    .Y ( ctsbuf_net_6482630 ) ) ;
sky130_fd_sc_hd__clkinvlp_4 cts_inv_4859050795 ( .A ( ctsbuf_net_6592641 ) , 
    .Y ( ctsbuf_net_6492631 ) ) ;
sky130_fd_sc_hd__clkinvlp_4 cts_inv_4859150796 ( .A ( ctsbuf_net_6592641 ) , 
    .Y ( ctsbuf_net_6502632 ) ) ;
sky130_fd_sc_hd__clkinvlp_4 cts_inv_4859250797 ( .A ( ctsbuf_net_6612643 ) , 
    .Y ( ctsbuf_net_6512633 ) ) ;
sky130_fd_sc_hd__clkinvlp_4 cts_inv_4859350798 ( .A ( ctsbuf_net_6582640 ) , 
    .Y ( ctsbuf_net_6522634 ) ) ;
sky130_fd_sc_hd__clkinvlp_4 cts_inv_4859450799 ( .A ( ctsbuf_net_6622644 ) , 
    .Y ( ctsbuf_net_6532635 ) ) ;
sky130_fd_sc_hd__clkinvlp_4 cts_inv_4859550800 ( .A ( ctsbuf_net_6602642 ) , 
    .Y ( ctsbuf_net_6542636 ) ) ;
sky130_fd_sc_hd__clkinv_1 cts_inv_4859650801 ( .A ( ctsbuf_net_6612643 ) , 
    .Y ( ctsbuf_net_6552637 ) ) ;
sky130_fd_sc_hd__clkinvlp_2 cts_inv_4859750802 ( .A ( ctsbuf_net_6612643 ) , 
    .Y ( ctsbuf_net_6562638 ) ) ;
sky130_fd_sc_hd__clkinvlp_2 cts_inv_4859850803 ( .A ( ctsbuf_net_6622644 ) , 
    .Y ( ctsbuf_net_6572639 ) ) ;
sky130_fd_sc_hd__clkinvlp_4 cts_inv_4861850823 ( .A ( prog_clk[0] ) , 
    .Y ( ctsbuf_net_6582640 ) ) ;
sky130_fd_sc_hd__clkinvlp_4 cts_inv_4861950824 ( .A ( prog_clk[0] ) , 
    .Y ( ctsbuf_net_6592641 ) ) ;
sky130_fd_sc_hd__clkinvlp_2 cts_inv_4862050825 ( .A ( prog_clk[0] ) , 
    .Y ( ctsbuf_net_6602642 ) ) ;
sky130_fd_sc_hd__clkinvlp_4 cts_inv_4862150826 ( .A ( prog_clk[0] ) , 
    .Y ( ctsbuf_net_6612643 ) ) ;
sky130_fd_sc_hd__clkinvlp_2 cts_inv_4862250827 ( .A ( prog_clk[0] ) , 
    .Y ( ctsbuf_net_6622644 ) ) ;
endmodule


