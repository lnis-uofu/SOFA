VERSION 5.7 ;
BUSBITCHARS "[]" ;

UNITS
  DATABASE MICRONS 1000 ;
END UNITS

MANUFACTURINGGRID 0.005 ;

LAYER li1
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.46 ;
  WIDTH 0.17 ;
END li1

LAYER mcon
  TYPE CUT ;
END mcon

LAYER met1
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.34 ;
  WIDTH 0.14 ;
END met1

LAYER via
  TYPE CUT ;
END via

LAYER met2
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.46 ;
  WIDTH 0.14 ;
END met2

LAYER via2
  TYPE CUT ;
END via2

LAYER met3
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.68 ;
  WIDTH 0.3 ;
END met3

LAYER via3
  TYPE CUT ;
END via3

LAYER met4
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.92 ;
  WIDTH 0.3 ;
END met4

LAYER via4
  TYPE CUT ;
END via4

LAYER met5
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 3.4 ;
  WIDTH 1.6 ;
END met5

LAYER nwell
  TYPE MASTERSLICE ;
END nwell

LAYER pwell
  TYPE MASTERSLICE ;
END pwell

LAYER OVERLAP
  TYPE OVERLAP ;
END OVERLAP

VIA L1M1_PR
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.145 -0.115 0.145 0.115 ;
END L1M1_PR

VIA L1M1_PR_R
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.115 -0.145 0.115 0.145 ;
END L1M1_PR_R

VIA L1M1_PR_M
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.115 -0.145 0.115 0.145 ;
END L1M1_PR_M

VIA L1M1_PR_MR
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.145 -0.115 0.145 0.115 ;
END L1M1_PR_MR

VIA L1M1_PR_C
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.145 -0.145 0.145 0.145 ;
END L1M1_PR_C

VIA M1M2_PR
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR

VIA M1M2_PR_Enc
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_Enc

VIA M1M2_PR_R
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_R

VIA M1M2_PR_R_Enc
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR_R_Enc

VIA M1M2_PR_M
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_M

VIA M1M2_PR_M_Enc
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR_M_Enc

VIA M1M2_PR_MR
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR_MR

VIA M1M2_PR_MR_Enc
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_MR_Enc

VIA M1M2_PR_C
  LAYER met1 ;
    RECT -0.16 -0.16 0.16 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.16 0.16 0.16 ;
END M1M2_PR_C

VIA M2M3_PR
  LAYER met2 ;
    RECT -0.14 -0.185 0.14 0.185 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR

VIA M2M3_PR_R
  LAYER met2 ;
    RECT -0.185 -0.14 0.185 0.14 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_R

VIA M2M3_PR_M
  LAYER met2 ;
    RECT -0.14 -0.185 0.14 0.185 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_M

VIA M2M3_PR_MR
  LAYER met2 ;
    RECT -0.185 -0.14 0.185 0.14 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_MR

VIA M2M3_PR_C
  LAYER met2 ;
    RECT -0.185 -0.185 0.185 0.185 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_C

VIA M3M4_PR
  LAYER met3 ;
    RECT -0.19 -0.16 0.19 0.16 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR

VIA M3M4_PR_R
  LAYER met3 ;
    RECT -0.16 -0.19 0.16 0.19 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_R

VIA M3M4_PR_M
  LAYER met3 ;
    RECT -0.19 -0.16 0.19 0.16 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_M

VIA M3M4_PR_MR
  LAYER met3 ;
    RECT -0.16 -0.19 0.16 0.19 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_MR

VIA M3M4_PR_C
  LAYER met3 ;
    RECT -0.19 -0.19 0.19 0.19 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_C

VIA M4M5_PR
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR

VIA M4M5_PR_R
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_R

VIA M4M5_PR_M
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_M

VIA M4M5_PR_MR
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_MR

VIA M4M5_PR_C
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_C

SITE unit
  CLASS CORE ;
  SYMMETRY Y ;
  SIZE 0.46 BY 2.72 ;
END unit

SITE unithddbl
  CLASS CORE ;
  SIZE 0.46 BY 5.44 ;
END unithddbl

MACRO sb_1__2_
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  SIZE 103.04 BY 81.6 ;
  SYMMETRY X Y ;
  PIN prog_clk[0]
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER met2 ;
        RECT 20.63 0 20.77 1.36 ;
    END
  END prog_clk[0]
  PIN chanx_right_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 101.66 54.25 103.04 54.55 ;
    END
  END chanx_right_in[0]
  PIN chanx_right_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 101.66 42.01 103.04 42.31 ;
    END
  END chanx_right_in[1]
  PIN chanx_right_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 101.66 56.29 103.04 56.59 ;
    END
  END chanx_right_in[2]
  PIN chanx_right_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 101.66 26.37 103.04 26.67 ;
    END
  END chanx_right_in[3]
  PIN chanx_right_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 101.66 35.89 103.04 36.19 ;
    END
  END chanx_right_in[4]
  PIN chanx_right_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 101.66 69.21 103.04 69.51 ;
    END
  END chanx_right_in[5]
  PIN chanx_right_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 101.66 33.17 103.04 33.47 ;
    END
  END chanx_right_in[6]
  PIN chanx_right_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 101.66 63.77 103.04 64.07 ;
    END
  END chanx_right_in[7]
  PIN chanx_right_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 101.66 43.37 103.04 43.67 ;
    END
  END chanx_right_in[8]
  PIN chanx_right_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 101.66 76.01 103.04 76.31 ;
    END
  END chanx_right_in[9]
  PIN chanx_right_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 101.66 40.65 103.04 40.95 ;
    END
  END chanx_right_in[10]
  PIN chanx_right_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 101.66 77.37 103.04 77.67 ;
    END
  END chanx_right_in[11]
  PIN chanx_right_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 101.66 59.01 103.04 59.31 ;
    END
  END chanx_right_in[12]
  PIN chanx_right_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 101.66 22.97 103.04 23.27 ;
    END
  END chanx_right_in[13]
  PIN chanx_right_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.67 16.32 100.81 17.68 ;
    END
  END chanx_right_in[14]
  PIN chanx_right_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 101.66 67.85 103.04 68.15 ;
    END
  END chanx_right_in[15]
  PIN chanx_right_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 101.66 44.73 103.04 45.03 ;
    END
  END chanx_right_in[16]
  PIN chanx_right_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 101.66 21.61 103.04 21.91 ;
    END
  END chanx_right_in[17]
  PIN chanx_right_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 101.66 61.05 103.04 61.35 ;
    END
  END chanx_right_in[18]
  PIN chanx_right_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 101.66 65.13 103.04 65.43 ;
    END
  END chanx_right_in[19]
  PIN right_top_grid_pin_1_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 101.66 37.25 103.04 37.55 ;
    END
  END right_top_grid_pin_1_[0]
  PIN right_bottom_grid_pin_34_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.91 16.32 98.05 17.68 ;
    END
  END right_bottom_grid_pin_34_[0]
  PIN right_bottom_grid_pin_35_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.75 16.32 99.89 17.68 ;
    END
  END right_bottom_grid_pin_35_[0]
  PIN right_bottom_grid_pin_36_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 97.37 16.32 97.67 17.68 ;
    END
  END right_bottom_grid_pin_36_[0]
  PIN right_bottom_grid_pin_37_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.23 16.32 94.37 17.68 ;
    END
  END right_bottom_grid_pin_37_[0]
  PIN right_bottom_grid_pin_38_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.15 16.32 95.29 17.68 ;
    END
  END right_bottom_grid_pin_38_[0]
  PIN right_bottom_grid_pin_39_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 83.26 5.29 84.64 5.59 ;
    END
  END right_bottom_grid_pin_39_[0]
  PIN right_bottom_grid_pin_40_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.53 16.32 96.67 17.68 ;
    END
  END right_bottom_grid_pin_40_[0]
  PIN right_bottom_grid_pin_41_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.27 0 82.41 1.36 ;
    END
  END right_bottom_grid_pin_41_[0]
  PIN chany_bottom_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.53 0 50.67 1.36 ;
    END
  END chany_bottom_in[0]
  PIN chany_bottom_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.89 0 58.03 1.36 ;
    END
  END chany_bottom_in[1]
  PIN chany_bottom_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.97 0 57.11 1.36 ;
    END
  END chany_bottom_in[2]
  PIN chany_bottom_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.49 0 62.63 1.36 ;
    END
  END chany_bottom_in[3]
  PIN chany_bottom_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.69 0 48.83 1.36 ;
    END
  END chany_bottom_in[4]
  PIN chany_bottom_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.19 0 60.33 1.36 ;
    END
  END chany_bottom_in[5]
  PIN chany_bottom_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.21 0 77.35 1.36 ;
    END
  END chany_bottom_in[6]
  PIN chany_bottom_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.37 0 52.51 1.36 ;
    END
  END chany_bottom_in[7]
  PIN chany_bottom_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.11 0 61.25 1.36 ;
    END
  END chany_bottom_in[8]
  PIN chany_bottom_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.41 0 40.55 1.36 ;
    END
  END chany_bottom_in[9]
  PIN chany_bottom_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.05 0 56.19 1.36 ;
    END
  END chany_bottom_in[10]
  PIN chany_bottom_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.61 0 49.75 1.36 ;
    END
  END chany_bottom_in[11]
  PIN chany_bottom_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.77 0 47.91 1.36 ;
    END
  END chany_bottom_in[12]
  PIN chany_bottom_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.23 0 71.37 1.36 ;
    END
  END chany_bottom_in[13]
  PIN chany_bottom_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.37 0 75.51 1.36 ;
    END
  END chany_bottom_in[14]
  PIN chany_bottom_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.59 0 32.73 1.36 ;
    END
  END chany_bottom_in[15]
  PIN chany_bottom_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.45 0 51.59 1.36 ;
    END
  END chany_bottom_in[16]
  PIN chany_bottom_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.45 0 74.59 1.36 ;
    END
  END chany_bottom_in[17]
  PIN chany_bottom_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.29 0 76.43 1.36 ;
    END
  END chany_bottom_in[18]
  PIN chany_bottom_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.21 0 54.35 1.36 ;
    END
  END chany_bottom_in[19]
  PIN bottom_left_grid_pin_42_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.61 16.32 3.75 17.68 ;
    END
  END bottom_left_grid_pin_42_[0]
  PIN bottom_left_grid_pin_43_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 22.85 0 23.15 1.36 ;
    END
  END bottom_left_grid_pin_43_[0]
  PIN bottom_left_grid_pin_44_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.51 16.32 10.65 17.68 ;
    END
  END bottom_left_grid_pin_44_[0]
  PIN bottom_left_grid_pin_45_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.53 16.32 4.67 17.68 ;
    END
  END bottom_left_grid_pin_45_[0]
  PIN bottom_left_grid_pin_46_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.69 16.32 2.83 17.68 ;
    END
  END bottom_left_grid_pin_46_[0]
  PIN bottom_left_grid_pin_47_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 18.4 12.09 19.78 12.39 ;
    END
  END bottom_left_grid_pin_47_[0]
  PIN bottom_left_grid_pin_48_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.83 16.32 6.97 17.68 ;
    END
  END bottom_left_grid_pin_48_[0]
  PIN bottom_left_grid_pin_49_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.59 16.32 9.73 17.68 ;
    END
  END bottom_left_grid_pin_49_[0]
  PIN chanx_left_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 27.05 1.38 27.35 ;
    END
  END chanx_left_in[0]
  PIN chanx_left_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 67.85 1.38 68.15 ;
    END
  END chanx_left_in[1]
  PIN chanx_left_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 70.57 1.38 70.87 ;
    END
  END chanx_left_in[2]
  PIN chanx_left_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 69.21 1.38 69.51 ;
    END
  END chanx_left_in[3]
  PIN chanx_left_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 37.93 1.38 38.23 ;
    END
  END chanx_left_in[4]
  PIN chanx_left_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 22.97 1.38 23.27 ;
    END
  END chanx_left_in[5]
  PIN chanx_left_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 65.13 1.38 65.43 ;
    END
  END chanx_left_in[6]
  PIN chanx_left_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 25.69 1.38 25.99 ;
    END
  END chanx_left_in[7]
  PIN chanx_left_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 46.09 1.38 46.39 ;
    END
  END chanx_left_in[8]
  PIN chanx_left_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 60.37 1.38 60.67 ;
    END
  END chanx_left_in[9]
  PIN chanx_left_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 63.77 1.38 64.07 ;
    END
  END chanx_left_in[10]
  PIN chanx_left_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 36.57 1.38 36.87 ;
    END
  END chanx_left_in[11]
  PIN chanx_left_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 29.77 1.38 30.07 ;
    END
  END chanx_left_in[12]
  PIN chanx_left_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 20.25 1.38 20.55 ;
    END
  END chanx_left_in[13]
  PIN chanx_left_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 77.37 1.38 77.67 ;
    END
  END chanx_left_in[14]
  PIN chanx_left_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 76.01 1.38 76.31 ;
    END
  END chanx_left_in[15]
  PIN chanx_left_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 59.01 1.38 59.31 ;
    END
  END chanx_left_in[16]
  PIN chanx_left_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 52.21 1.38 52.51 ;
    END
  END chanx_left_in[17]
  PIN chanx_left_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 40.65 1.38 40.95 ;
    END
  END chanx_left_in[18]
  PIN chanx_left_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 24.33 1.38 24.63 ;
    END
  END chanx_left_in[19]
  PIN left_top_grid_pin_1_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 62.41 1.38 62.71 ;
    END
  END left_top_grid_pin_1_[0]
  PIN left_bottom_grid_pin_34_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 18.4 6.65 19.78 6.95 ;
    END
  END left_bottom_grid_pin_34_[0]
  PIN left_bottom_grid_pin_35_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 4.45 16.32 4.75 17.68 ;
    END
  END left_bottom_grid_pin_35_[0]
  PIN left_bottom_grid_pin_36_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 18.4 5.29 19.78 5.59 ;
    END
  END left_bottom_grid_pin_36_[0]
  PIN left_bottom_grid_pin_37_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.45 16.32 5.59 17.68 ;
    END
  END left_bottom_grid_pin_37_[0]
  PIN left_bottom_grid_pin_38_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.01 0 22.15 1.36 ;
    END
  END left_bottom_grid_pin_38_[0]
  PIN left_bottom_grid_pin_39_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.67 16.32 8.81 17.68 ;
    END
  END left_bottom_grid_pin_39_[0]
  PIN left_bottom_grid_pin_40_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.93 0 23.07 1.36 ;
    END
  END left_bottom_grid_pin_40_[0]
  PIN left_bottom_grid_pin_41_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.75 16.32 7.89 17.68 ;
    END
  END left_bottom_grid_pin_41_[0]
  PIN ccff_head[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 101.66 47.45 103.04 47.75 ;
    END
  END ccff_head[0]
  PIN chanx_right_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 101.66 52.89 103.04 53.19 ;
    END
  END chanx_right_out[0]
  PIN chanx_right_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 101.66 29.09 103.04 29.39 ;
    END
  END chanx_right_out[1]
  PIN chanx_right_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 101.66 50.17 103.04 50.47 ;
    END
  END chanx_right_out[2]
  PIN chanx_right_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 101.66 31.81 103.04 32.11 ;
    END
  END chanx_right_out[3]
  PIN chanx_right_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 101.66 70.57 103.04 70.87 ;
    END
  END chanx_right_out[4]
  PIN chanx_right_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 101.66 24.33 103.04 24.63 ;
    END
  END chanx_right_out[5]
  PIN chanx_right_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 101.66 66.49 103.04 66.79 ;
    END
  END chanx_right_out[6]
  PIN chanx_right_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 101.66 51.53 103.04 51.83 ;
    END
  END chanx_right_out[7]
  PIN chanx_right_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 101.66 34.53 103.04 34.83 ;
    END
  END chanx_right_out[8]
  PIN chanx_right_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 101.66 20.25 103.04 20.55 ;
    END
  END chanx_right_out[9]
  PIN chanx_right_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 101.66 71.93 103.04 72.23 ;
    END
  END chanx_right_out[10]
  PIN chanx_right_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 101.66 30.45 103.04 30.75 ;
    END
  END chanx_right_out[11]
  PIN chanx_right_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 101.66 39.29 103.04 39.59 ;
    END
  END chanx_right_out[12]
  PIN chanx_right_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 101.66 27.73 103.04 28.03 ;
    END
  END chanx_right_out[13]
  PIN chanx_right_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 101.66 48.81 103.04 49.11 ;
    END
  END chanx_right_out[14]
  PIN chanx_right_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 101.66 74.65 103.04 74.95 ;
    END
  END chanx_right_out[15]
  PIN chanx_right_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 101.66 57.65 103.04 57.95 ;
    END
  END chanx_right_out[16]
  PIN chanx_right_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 101.66 46.09 103.04 46.39 ;
    END
  END chanx_right_out[17]
  PIN chanx_right_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 101.66 73.29 103.04 73.59 ;
    END
  END chanx_right_out[18]
  PIN chanx_right_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 101.66 62.41 103.04 62.71 ;
    END
  END chanx_right_out[19]
  PIN chany_bottom_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.15 0 72.29 1.36 ;
    END
  END chany_bottom_out[0]
  PIN chany_bottom_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.13 0 55.27 1.36 ;
    END
  END chany_bottom_out[1]
  PIN chany_bottom_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.85 0 46.99 1.36 ;
    END
  END chany_bottom_out[2]
  PIN chany_bottom_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.41 0 63.55 1.36 ;
    END
  END chany_bottom_out[3]
  PIN chany_bottom_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.93 0 46.07 1.36 ;
    END
  END chany_bottom_out[4]
  PIN chany_bottom_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.31 0 70.45 1.36 ;
    END
  END chany_bottom_out[5]
  PIN chany_bottom_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.51 0 33.65 1.36 ;
    END
  END chany_bottom_out[6]
  PIN chany_bottom_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.79 0 64.93 1.36 ;
    END
  END chany_bottom_out[7]
  PIN chany_bottom_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.27 0 59.41 1.36 ;
    END
  END chany_bottom_out[8]
  PIN chany_bottom_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.71 0 65.85 1.36 ;
    END
  END chany_bottom_out[9]
  PIN chany_bottom_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.17 0 43.31 1.36 ;
    END
  END chany_bottom_out[10]
  PIN chany_bottom_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.63 0 66.77 1.36 ;
    END
  END chany_bottom_out[11]
  PIN chany_bottom_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.49 0 39.63 1.36 ;
    END
  END chany_bottom_out[12]
  PIN chany_bottom_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.55 0 67.69 1.36 ;
    END
  END chany_bottom_out[13]
  PIN chany_bottom_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.25 0 42.39 1.36 ;
    END
  END chany_bottom_out[14]
  PIN chany_bottom_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.89 0 81.03 1.36 ;
    END
  END chany_bottom_out[15]
  PIN chany_bottom_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.33 0 41.47 1.36 ;
    END
  END chany_bottom_out[16]
  PIN chany_bottom_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.47 0 68.61 1.36 ;
    END
  END chany_bottom_out[17]
  PIN chany_bottom_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.01 0 45.15 1.36 ;
    END
  END chany_bottom_out[18]
  PIN chany_bottom_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.39 0 69.53 1.36 ;
    END
  END chany_bottom_out[19]
  PIN chanx_left_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 57.65 1.38 57.95 ;
    END
  END chanx_left_out[0]
  PIN chanx_left_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 66.49 1.38 66.79 ;
    END
  END chanx_left_out[1]
  PIN chanx_left_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 55.61 1.38 55.91 ;
    END
  END chanx_left_out[2]
  PIN chanx_left_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 47.45 1.38 47.75 ;
    END
  END chanx_left_out[3]
  PIN chanx_left_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 50.85 1.38 51.15 ;
    END
  END chanx_left_out[4]
  PIN chanx_left_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 28.41 1.38 28.71 ;
    END
  END chanx_left_out[5]
  PIN chanx_left_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 43.37 1.38 43.67 ;
    END
  END chanx_left_out[6]
  PIN chanx_left_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 31.13 1.38 31.43 ;
    END
  END chanx_left_out[7]
  PIN chanx_left_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 73.29 1.38 73.59 ;
    END
  END chanx_left_out[8]
  PIN chanx_left_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 6.29 16.32 6.59 17.68 ;
    END
  END chanx_left_out[9]
  PIN chanx_left_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 74.65 1.38 74.95 ;
    END
  END chanx_left_out[10]
  PIN chanx_left_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 35.21 1.38 35.51 ;
    END
  END chanx_left_out[11]
  PIN chanx_left_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 71.93 1.38 72.23 ;
    END
  END chanx_left_out[12]
  PIN chanx_left_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 53.57 1.38 53.87 ;
    END
  END chanx_left_out[13]
  PIN chanx_left_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 42.01 1.38 42.31 ;
    END
  END chanx_left_out[14]
  PIN chanx_left_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 48.81 1.38 49.11 ;
    END
  END chanx_left_out[15]
  PIN chanx_left_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 33.85 1.38 34.15 ;
    END
  END chanx_left_out[16]
  PIN chanx_left_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 32.49 1.38 32.79 ;
    END
  END chanx_left_out[17]
  PIN chanx_left_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 44.73 1.38 45.03 ;
    END
  END chanx_left_out[18]
  PIN chanx_left_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 39.29 1.38 39.59 ;
    END
  END chanx_left_out[19]
  PIN ccff_tail[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 21.61 1.38 21.91 ;
    END
  END ccff_tail[0]
  PIN SC_IN_TOP
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.21 80.24 54.35 81.6 ;
    END
  END SC_IN_TOP
  PIN SC_IN_BOT
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.29 80.24 53.43 81.6 ;
    END
  END SC_IN_BOT
  PIN SC_OUT_TOP
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.37 80.24 52.51 81.6 ;
    END
  END SC_OUT_TOP
  PIN SC_OUT_BOT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.45 80.24 51.59 81.6 ;
    END
  END SC_OUT_BOT
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 18.4 2.48 18.88 2.96 ;
        RECT 84.16 2.48 84.64 2.96 ;
        RECT 18.4 7.92 18.88 8.4 ;
        RECT 84.16 7.92 84.64 8.4 ;
        RECT 18.4 13.36 18.88 13.84 ;
        RECT 84.16 13.36 84.64 13.84 ;
        RECT 0 18.8 0.48 19.28 ;
        RECT 102.56 18.8 103.04 19.28 ;
        RECT 0 24.24 0.48 24.72 ;
        RECT 102.56 24.24 103.04 24.72 ;
        RECT 0 29.68 0.48 30.16 ;
        RECT 102.56 29.68 103.04 30.16 ;
        RECT 0 35.12 0.48 35.6 ;
        RECT 102.56 35.12 103.04 35.6 ;
        RECT 0 40.56 0.48 41.04 ;
        RECT 102.56 40.56 103.04 41.04 ;
        RECT 0 46 0.48 46.48 ;
        RECT 102.56 46 103.04 46.48 ;
        RECT 0 51.44 0.48 51.92 ;
        RECT 102.56 51.44 103.04 51.92 ;
        RECT 0 56.88 0.48 57.36 ;
        RECT 102.56 56.88 103.04 57.36 ;
        RECT 0 62.32 0.48 62.8 ;
        RECT 102.56 62.32 103.04 62.8 ;
        RECT 0 67.76 0.48 68.24 ;
        RECT 102.56 67.76 103.04 68.24 ;
        RECT 0 73.2 0.48 73.68 ;
        RECT 102.56 73.2 103.04 73.68 ;
        RECT 0 78.64 0.48 79.12 ;
        RECT 102.56 78.64 103.04 79.12 ;
      LAYER met4 ;
        RECT 29.14 0 29.74 0.6 ;
        RECT 58.58 0 59.18 0.6 ;
        RECT 29.14 81 29.74 81.6 ;
        RECT 58.58 81 59.18 81.6 ;
      LAYER met5 ;
        RECT 0 26.96 3.2 30.16 ;
        RECT 99.84 26.96 103.04 30.16 ;
        RECT 0 67.76 3.2 70.96 ;
        RECT 99.84 67.76 103.04 70.96 ;
    END
  END VDD
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 18.4 0 84.64 0.24 ;
        RECT 18.4 5.2 18.88 5.68 ;
        RECT 84.16 5.2 84.64 5.68 ;
        RECT 18.4 10.64 18.88 11.12 ;
        RECT 84.16 10.64 84.64 11.12 ;
        RECT 0 16.08 103.04 16.56 ;
        RECT 0 21.52 0.48 22 ;
        RECT 102.56 21.52 103.04 22 ;
        RECT 0 26.96 0.48 27.44 ;
        RECT 102.56 26.96 103.04 27.44 ;
        RECT 0 32.4 0.48 32.88 ;
        RECT 102.56 32.4 103.04 32.88 ;
        RECT 0 37.84 0.48 38.32 ;
        RECT 102.56 37.84 103.04 38.32 ;
        RECT 0 43.28 0.48 43.76 ;
        RECT 102.56 43.28 103.04 43.76 ;
        RECT 0 48.72 0.48 49.2 ;
        RECT 102.56 48.72 103.04 49.2 ;
        RECT 0 54.16 0.48 54.64 ;
        RECT 102.56 54.16 103.04 54.64 ;
        RECT 0 59.6 0.48 60.08 ;
        RECT 102.56 59.6 103.04 60.08 ;
        RECT 0 65.04 0.48 65.52 ;
        RECT 102.56 65.04 103.04 65.52 ;
        RECT 0 70.48 0.48 70.96 ;
        RECT 102.56 70.48 103.04 70.96 ;
        RECT 0 75.92 0.48 76.4 ;
        RECT 102.56 75.92 103.04 76.4 ;
        RECT 0 81.36 103.04 81.6 ;
      LAYER met4 ;
        RECT 43.86 0 44.46 0.6 ;
        RECT 73.3 0 73.9 0.6 ;
        RECT 43.86 81 44.46 81.6 ;
        RECT 73.3 81 73.9 81.6 ;
      LAYER met5 ;
        RECT 0 47.36 3.2 50.56 ;
        RECT 99.84 47.36 103.04 50.56 ;
    END
  END VSS
  OBS
    LAYER li1 ;
      RECT 0 81.515 103.04 81.685 ;
      RECT 102.12 78.795 103.04 78.965 ;
      RECT 0 78.795 3.68 78.965 ;
      RECT 102.12 76.075 103.04 76.245 ;
      RECT 0 76.075 1.84 76.245 ;
      RECT 99.36 73.355 103.04 73.525 ;
      RECT 0 73.355 1.84 73.525 ;
      RECT 99.36 70.635 103.04 70.805 ;
      RECT 0 70.635 1.84 70.805 ;
      RECT 102.12 67.915 103.04 68.085 ;
      RECT 0 67.915 1.84 68.085 ;
      RECT 102.12 65.195 103.04 65.365 ;
      RECT 0 65.195 1.84 65.365 ;
      RECT 102.12 62.475 103.04 62.645 ;
      RECT 0 62.475 1.84 62.645 ;
      RECT 102.12 59.755 103.04 59.925 ;
      RECT 0 59.755 1.84 59.925 ;
      RECT 102.12 57.035 103.04 57.205 ;
      RECT 0 57.035 1.84 57.205 ;
      RECT 102.12 54.315 103.04 54.485 ;
      RECT 0 54.315 1.84 54.485 ;
      RECT 102.12 51.595 103.04 51.765 ;
      RECT 0 51.595 1.84 51.765 ;
      RECT 102.12 48.875 103.04 49.045 ;
      RECT 0 48.875 1.84 49.045 ;
      RECT 102.12 46.155 103.04 46.325 ;
      RECT 0 46.155 1.84 46.325 ;
      RECT 102.12 43.435 103.04 43.605 ;
      RECT 0 43.435 1.84 43.605 ;
      RECT 102.12 40.715 103.04 40.885 ;
      RECT 0 40.715 1.84 40.885 ;
      RECT 102.12 37.995 103.04 38.165 ;
      RECT 0 37.995 1.84 38.165 ;
      RECT 102.12 35.275 103.04 35.445 ;
      RECT 0 35.275 1.84 35.445 ;
      RECT 102.12 32.555 103.04 32.725 ;
      RECT 0 32.555 1.84 32.725 ;
      RECT 102.12 29.835 103.04 30.005 ;
      RECT 0 29.835 1.84 30.005 ;
      RECT 102.12 27.115 103.04 27.285 ;
      RECT 0 27.115 1.84 27.285 ;
      RECT 102.12 24.395 103.04 24.565 ;
      RECT 0 24.395 1.84 24.565 ;
      RECT 102.12 21.675 103.04 21.845 ;
      RECT 0 21.675 1.84 21.845 ;
      RECT 102.12 18.955 103.04 19.125 ;
      RECT 0 18.955 3.68 19.125 ;
      RECT 82.34 16.235 103.04 16.405 ;
      RECT 0 16.235 22.08 16.405 ;
      RECT 83.72 13.515 84.64 13.685 ;
      RECT 18.4 13.515 22.08 13.685 ;
      RECT 83.72 10.795 84.64 10.965 ;
      RECT 18.4 10.795 22.08 10.965 ;
      RECT 83.72 8.075 84.64 8.245 ;
      RECT 18.4 8.075 22.08 8.245 ;
      RECT 83.72 5.355 84.64 5.525 ;
      RECT 18.4 5.355 22.08 5.525 ;
      RECT 83.72 2.635 84.64 2.805 ;
      RECT 18.4 2.635 22.08 2.805 ;
      RECT 18.4 -0.085 84.64 0.085 ;
    LAYER met2 ;
      RECT 73.46 81.415 73.74 81.785 ;
      RECT 44.02 81.415 44.3 81.785 ;
      RECT 53.69 1.54 53.95 1.86 ;
      RECT 47.25 1.54 47.51 1.86 ;
      RECT 73.46 -0.185 73.74 0.185 ;
      RECT 44.02 -0.185 44.3 0.185 ;
      POLYGON 102.76 81.32 102.76 16.6 101.09 16.6 101.09 17.96 100.39 17.96 100.39 16.6 100.17 16.6 100.17 17.96 99.47 17.96 99.47 16.6 98.33 16.6 98.33 17.96 97.63 17.96 97.63 16.6 96.95 16.6 96.95 17.96 96.25 17.96 96.25 16.6 95.57 16.6 95.57 17.96 94.87 17.96 94.87 16.6 94.65 16.6 94.65 17.96 93.95 17.96 93.95 16.6 84.36 16.6 84.36 0.28 82.69 0.28 82.69 1.64 81.99 1.64 81.99 0.28 81.31 0.28 81.31 1.64 80.61 1.64 80.61 0.28 77.63 0.28 77.63 1.64 76.93 1.64 76.93 0.28 76.71 0.28 76.71 1.64 76.01 1.64 76.01 0.28 75.79 0.28 75.79 1.64 75.09 1.64 75.09 0.28 74.87 0.28 74.87 1.64 74.17 1.64 74.17 0.28 72.57 0.28 72.57 1.64 71.87 1.64 71.87 0.28 71.65 0.28 71.65 1.64 70.95 1.64 70.95 0.28 70.73 0.28 70.73 1.64 70.03 1.64 70.03 0.28 69.81 0.28 69.81 1.64 69.11 1.64 69.11 0.28 68.89 0.28 68.89 1.64 68.19 1.64 68.19 0.28 67.97 0.28 67.97 1.64 67.27 1.64 67.27 0.28 67.05 0.28 67.05 1.64 66.35 1.64 66.35 0.28 66.13 0.28 66.13 1.64 65.43 1.64 65.43 0.28 65.21 0.28 65.21 1.64 64.51 1.64 64.51 0.28 63.83 0.28 63.83 1.64 63.13 1.64 63.13 0.28 62.91 0.28 62.91 1.64 62.21 1.64 62.21 0.28 61.53 0.28 61.53 1.64 60.83 1.64 60.83 0.28 60.61 0.28 60.61 1.64 59.91 1.64 59.91 0.28 59.69 0.28 59.69 1.64 58.99 1.64 58.99 0.28 58.31 0.28 58.31 1.64 57.61 1.64 57.61 0.28 57.39 0.28 57.39 1.64 56.69 1.64 56.69 0.28 56.47 0.28 56.47 1.64 55.77 1.64 55.77 0.28 55.55 0.28 55.55 1.64 54.85 1.64 54.85 0.28 54.63 0.28 54.63 1.64 53.93 1.64 53.93 0.28 52.79 0.28 52.79 1.64 52.09 1.64 52.09 0.28 51.87 0.28 51.87 1.64 51.17 1.64 51.17 0.28 50.95 0.28 50.95 1.64 50.25 1.64 50.25 0.28 50.03 0.28 50.03 1.64 49.33 1.64 49.33 0.28 49.11 0.28 49.11 1.64 48.41 1.64 48.41 0.28 48.19 0.28 48.19 1.64 47.49 1.64 47.49 0.28 47.27 0.28 47.27 1.64 46.57 1.64 46.57 0.28 46.35 0.28 46.35 1.64 45.65 1.64 45.65 0.28 45.43 0.28 45.43 1.64 44.73 1.64 44.73 0.28 43.59 0.28 43.59 1.64 42.89 1.64 42.89 0.28 42.67 0.28 42.67 1.64 41.97 1.64 41.97 0.28 41.75 0.28 41.75 1.64 41.05 1.64 41.05 0.28 40.83 0.28 40.83 1.64 40.13 1.64 40.13 0.28 39.91 0.28 39.91 1.64 39.21 1.64 39.21 0.28 33.93 0.28 33.93 1.64 33.23 1.64 33.23 0.28 33.01 0.28 33.01 1.64 32.31 1.64 32.31 0.28 23.35 0.28 23.35 1.64 22.65 1.64 22.65 0.28 22.43 0.28 22.43 1.64 21.73 1.64 21.73 0.28 21.05 0.28 21.05 1.64 20.35 1.64 20.35 0.28 18.68 0.28 18.68 16.6 10.93 16.6 10.93 17.96 10.23 17.96 10.23 16.6 10.01 16.6 10.01 17.96 9.31 17.96 9.31 16.6 9.09 16.6 9.09 17.96 8.39 17.96 8.39 16.6 8.17 16.6 8.17 17.96 7.47 17.96 7.47 16.6 7.25 16.6 7.25 17.96 6.55 17.96 6.55 16.6 5.87 16.6 5.87 17.96 5.17 17.96 5.17 16.6 4.95 16.6 4.95 17.96 4.25 17.96 4.25 16.6 4.03 16.6 4.03 17.96 3.33 17.96 3.33 16.6 3.11 16.6 3.11 17.96 2.41 17.96 2.41 16.6 0.28 16.6 0.28 81.32 51.17 81.32 51.17 79.96 51.87 79.96 51.87 81.32 52.09 81.32 52.09 79.96 52.79 79.96 52.79 81.32 53.01 81.32 53.01 79.96 53.71 79.96 53.71 81.32 53.93 81.32 53.93 79.96 54.63 79.96 54.63 81.32 ;
    LAYER met3 ;
      POLYGON 73.765 81.765 73.765 81.76 73.98 81.76 73.98 81.44 73.765 81.44 73.765 81.435 73.435 81.435 73.435 81.44 73.22 81.44 73.22 81.76 73.435 81.76 73.435 81.765 ;
      POLYGON 44.325 81.765 44.325 81.76 44.54 81.76 44.54 81.44 44.325 81.44 44.325 81.435 43.995 81.435 43.995 81.44 43.78 81.44 43.78 81.76 43.995 81.76 43.995 81.765 ;
      POLYGON 8.89 72.91 8.89 72.61 1.99 72.61 1.99 71.93 1.78 71.93 1.78 72.63 1.69 72.63 1.69 72.91 ;
      POLYGON 101.81 49.79 101.81 49.51 101.26 49.51 101.26 49.49 99.67 49.49 99.67 49.79 ;
      POLYGON 101.365 38.925 101.365 38.595 101.035 38.595 101.035 38.61 91.85 38.61 91.85 38.91 101.035 38.91 101.035 38.925 ;
      POLYGON 1.545 36.205 1.545 36.2 2.03 36.2 2.03 35.88 1.545 35.88 1.545 35.875 1.215 35.875 1.215 36.205 ;
      POLYGON 2.005 28.045 2.005 28.04 2.03 28.04 2.03 27.72 2.005 27.72 2.005 27.715 1.675 27.715 1.675 27.72 0.97 27.72 0.97 28.04 1.675 28.04 1.675 28.045 ;
      POLYGON 101.81 23.95 101.81 23.67 101.26 23.67 101.26 23.65 51.37 23.65 51.37 23.95 ;
      POLYGON 20.405 13.085 20.405 13.08 20.43 13.08 20.43 12.76 20.405 12.76 20.405 12.755 19.675 12.755 19.675 13.085 ;
      POLYGON 73.765 0.165 73.765 0.16 73.98 0.16 73.98 -0.16 73.765 -0.16 73.765 -0.165 73.435 -0.165 73.435 -0.16 73.22 -0.16 73.22 0.16 73.435 0.16 73.435 0.165 ;
      POLYGON 44.325 0.165 44.325 0.16 44.54 0.16 44.54 -0.16 44.325 -0.16 44.325 -0.165 43.995 -0.165 43.995 -0.16 43.78 -0.16 43.78 0.16 43.995 0.16 43.995 0.165 ;
      POLYGON 102.64 81.2 102.64 78.07 101.26 78.07 101.26 76.97 102.64 76.97 102.64 76.71 101.26 76.71 101.26 75.61 102.64 75.61 102.64 75.35 101.26 75.35 101.26 74.25 102.64 74.25 102.64 73.99 101.26 73.99 101.26 72.89 102.64 72.89 102.64 72.63 101.26 72.63 101.26 71.53 102.64 71.53 102.64 71.27 101.26 71.27 101.26 70.17 102.64 70.17 102.64 69.91 101.26 69.91 101.26 68.81 102.64 68.81 102.64 68.55 101.26 68.55 101.26 67.45 102.64 67.45 102.64 67.19 101.26 67.19 101.26 66.09 102.64 66.09 102.64 65.83 101.26 65.83 101.26 64.73 102.64 64.73 102.64 64.47 101.26 64.47 101.26 63.37 102.64 63.37 102.64 63.11 101.26 63.11 101.26 62.01 102.64 62.01 102.64 61.75 101.26 61.75 101.26 60.65 102.64 60.65 102.64 59.71 101.26 59.71 101.26 58.61 102.64 58.61 102.64 58.35 101.26 58.35 101.26 57.25 102.64 57.25 102.64 56.99 101.26 56.99 101.26 55.89 102.64 55.89 102.64 54.95 101.26 54.95 101.26 53.85 102.64 53.85 102.64 53.59 101.26 53.59 101.26 52.49 102.64 52.49 102.64 52.23 101.26 52.23 101.26 51.13 102.64 51.13 102.64 50.87 101.26 50.87 101.26 49.77 102.64 49.77 102.64 49.51 101.26 49.51 101.26 48.41 102.64 48.41 102.64 48.15 101.26 48.15 101.26 47.05 102.64 47.05 102.64 46.79 101.26 46.79 101.26 45.69 102.64 45.69 102.64 45.43 101.26 45.43 101.26 44.33 102.64 44.33 102.64 44.07 101.26 44.07 101.26 42.97 102.64 42.97 102.64 42.71 101.26 42.71 101.26 41.61 102.64 41.61 102.64 41.35 101.26 41.35 101.26 40.25 102.64 40.25 102.64 39.99 101.26 39.99 101.26 38.89 102.64 38.89 102.64 37.95 101.26 37.95 101.26 36.85 102.64 36.85 102.64 36.59 101.26 36.59 101.26 35.49 102.64 35.49 102.64 35.23 101.26 35.23 101.26 34.13 102.64 34.13 102.64 33.87 101.26 33.87 101.26 32.77 102.64 32.77 102.64 32.51 101.26 32.51 101.26 31.41 102.64 31.41 102.64 31.15 101.26 31.15 101.26 30.05 102.64 30.05 102.64 29.79 101.26 29.79 101.26 28.69 102.64 28.69 102.64 28.43 101.26 28.43 101.26 27.33 102.64 27.33 102.64 27.07 101.26 27.07 101.26 25.97 102.64 25.97 102.64 25.03 101.26 25.03 101.26 23.93 102.64 23.93 102.64 23.67 101.26 23.67 101.26 22.57 102.64 22.57 102.64 22.31 101.26 22.31 101.26 21.21 102.64 21.21 102.64 20.95 101.26 20.95 101.26 19.85 102.64 19.85 102.64 16.72 84.24 16.72 84.24 5.99 82.86 5.99 82.86 4.89 84.24 4.89 84.24 0.4 18.8 0.4 18.8 4.89 20.18 4.89 20.18 5.99 18.8 5.99 18.8 6.25 20.18 6.25 20.18 7.35 18.8 7.35 18.8 11.69 20.18 11.69 20.18 12.79 18.8 12.79 18.8 16.72 0.4 16.72 0.4 19.85 1.78 19.85 1.78 20.95 0.4 20.95 0.4 21.21 1.78 21.21 1.78 22.31 0.4 22.31 0.4 22.57 1.78 22.57 1.78 23.67 0.4 23.67 0.4 23.93 1.78 23.93 1.78 25.03 0.4 25.03 0.4 25.29 1.78 25.29 1.78 26.39 0.4 26.39 0.4 26.65 1.78 26.65 1.78 27.75 0.4 27.75 0.4 28.01 1.78 28.01 1.78 29.11 0.4 29.11 0.4 29.37 1.78 29.37 1.78 30.47 0.4 30.47 0.4 30.73 1.78 30.73 1.78 31.83 0.4 31.83 0.4 32.09 1.78 32.09 1.78 33.19 0.4 33.19 0.4 33.45 1.78 33.45 1.78 34.55 0.4 34.55 0.4 34.81 1.78 34.81 1.78 35.91 0.4 35.91 0.4 36.17 1.78 36.17 1.78 37.27 0.4 37.27 0.4 37.53 1.78 37.53 1.78 38.63 0.4 38.63 0.4 38.89 1.78 38.89 1.78 39.99 0.4 39.99 0.4 40.25 1.78 40.25 1.78 41.35 0.4 41.35 0.4 41.61 1.78 41.61 1.78 42.71 0.4 42.71 0.4 42.97 1.78 42.97 1.78 44.07 0.4 44.07 0.4 44.33 1.78 44.33 1.78 45.43 0.4 45.43 0.4 45.69 1.78 45.69 1.78 46.79 0.4 46.79 0.4 47.05 1.78 47.05 1.78 48.15 0.4 48.15 0.4 48.41 1.78 48.41 1.78 49.51 0.4 49.51 0.4 50.45 1.78 50.45 1.78 51.55 0.4 51.55 0.4 51.81 1.78 51.81 1.78 52.91 0.4 52.91 0.4 53.17 1.78 53.17 1.78 54.27 0.4 54.27 0.4 55.21 1.78 55.21 1.78 56.31 0.4 56.31 0.4 57.25 1.78 57.25 1.78 58.35 0.4 58.35 0.4 58.61 1.78 58.61 1.78 59.71 0.4 59.71 0.4 59.97 1.78 59.97 1.78 61.07 0.4 61.07 0.4 62.01 1.78 62.01 1.78 63.11 0.4 63.11 0.4 63.37 1.78 63.37 1.78 64.47 0.4 64.47 0.4 64.73 1.78 64.73 1.78 65.83 0.4 65.83 0.4 66.09 1.78 66.09 1.78 67.19 0.4 67.19 0.4 67.45 1.78 67.45 1.78 68.55 0.4 68.55 0.4 68.81 1.78 68.81 1.78 69.91 0.4 69.91 0.4 70.17 1.78 70.17 1.78 71.27 0.4 71.27 0.4 71.53 1.78 71.53 1.78 72.63 0.4 72.63 0.4 72.89 1.78 72.89 1.78 73.99 0.4 73.99 0.4 74.25 1.78 74.25 1.78 75.35 0.4 75.35 0.4 75.61 1.78 75.61 1.78 76.71 0.4 76.71 0.4 76.97 1.78 76.97 1.78 78.07 0.4 78.07 0.4 81.2 ;
    LAYER met4 ;
      POLYGON 102.64 81.2 102.64 16.72 98.07 16.72 98.07 18.08 96.97 18.08 96.97 16.72 84.24 16.72 84.24 0.4 74.3 0.4 74.3 1 72.9 1 72.9 0.4 59.58 0.4 59.58 1 58.18 1 58.18 0.4 44.86 0.4 44.86 1 43.46 1 43.46 0.4 30.14 0.4 30.14 1 28.74 1 28.74 0.4 23.55 0.4 23.55 1.76 22.45 1.76 22.45 0.4 18.8 0.4 18.8 16.72 6.99 16.72 6.99 18.08 5.89 18.08 5.89 16.72 5.15 16.72 5.15 18.08 4.05 18.08 4.05 16.72 0.4 16.72 0.4 81.2 28.74 81.2 28.74 80.6 30.14 80.6 30.14 81.2 43.46 81.2 43.46 80.6 44.86 80.6 44.86 81.2 58.18 81.2 58.18 80.6 59.58 80.6 59.58 81.2 72.9 81.2 72.9 80.6 74.3 80.6 74.3 81.2 ;
    LAYER met5 ;
      POLYGON 101.44 80 101.44 72.56 98.24 72.56 98.24 66.16 101.44 66.16 101.44 52.16 98.24 52.16 98.24 45.76 101.44 45.76 101.44 31.76 98.24 31.76 98.24 25.36 101.44 25.36 101.44 17.92 83.04 17.92 83.04 1.6 20 1.6 20 17.92 1.6 17.92 1.6 25.36 4.8 25.36 4.8 31.76 1.6 31.76 1.6 45.76 4.8 45.76 4.8 52.16 1.6 52.16 1.6 66.16 4.8 66.16 4.8 72.56 1.6 72.56 1.6 80 ;
    LAYER met1 ;
      POLYGON 102.76 81.08 102.76 79.4 102.28 79.4 102.28 78.36 102.76 78.36 102.76 76.68 102.28 76.68 102.28 75.64 102.76 75.64 102.76 73.96 102.28 73.96 102.28 72.92 102.76 72.92 102.76 71.24 102.28 71.24 102.28 70.2 102.76 70.2 102.76 68.52 102.28 68.52 102.28 67.48 102.76 67.48 102.76 65.8 102.28 65.8 102.28 64.76 102.76 64.76 102.76 63.08 102.28 63.08 102.28 62.04 102.76 62.04 102.76 60.36 102.28 60.36 102.28 59.32 102.76 59.32 102.76 57.64 102.28 57.64 102.28 56.6 102.76 56.6 102.76 54.92 102.28 54.92 102.28 53.88 102.76 53.88 102.76 52.2 102.28 52.2 102.28 51.16 102.76 51.16 102.76 49.48 102.28 49.48 102.28 48.44 102.76 48.44 102.76 46.76 102.28 46.76 102.28 45.72 102.76 45.72 102.76 44.04 102.28 44.04 102.28 43 102.76 43 102.76 41.32 102.28 41.32 102.28 40.28 102.76 40.28 102.76 38.6 102.28 38.6 102.28 37.56 102.76 37.56 102.76 35.88 102.28 35.88 102.28 34.84 102.76 34.84 102.76 33.16 102.28 33.16 102.28 32.12 102.76 32.12 102.76 30.44 102.28 30.44 102.28 29.4 102.76 29.4 102.76 27.72 102.28 27.72 102.28 26.68 102.76 26.68 102.76 25 102.28 25 102.28 23.96 102.76 23.96 102.76 22.28 102.28 22.28 102.28 21.24 102.76 21.24 102.76 19.56 102.28 19.56 102.28 18.52 102.76 18.52 102.76 16.84 0.28 16.84 0.28 18.52 0.76 18.52 0.76 19.56 0.28 19.56 0.28 21.24 0.76 21.24 0.76 22.28 0.28 22.28 0.28 23.96 0.76 23.96 0.76 25 0.28 25 0.28 26.68 0.76 26.68 0.76 27.72 0.28 27.72 0.28 29.4 0.76 29.4 0.76 30.44 0.28 30.44 0.28 32.12 0.76 32.12 0.76 33.16 0.28 33.16 0.28 34.84 0.76 34.84 0.76 35.88 0.28 35.88 0.28 37.56 0.76 37.56 0.76 38.6 0.28 38.6 0.28 40.28 0.76 40.28 0.76 41.32 0.28 41.32 0.28 43 0.76 43 0.76 44.04 0.28 44.04 0.28 45.72 0.76 45.72 0.76 46.76 0.28 46.76 0.28 48.44 0.76 48.44 0.76 49.48 0.28 49.48 0.28 51.16 0.76 51.16 0.76 52.2 0.28 52.2 0.28 53.88 0.76 53.88 0.76 54.92 0.28 54.92 0.28 56.6 0.76 56.6 0.76 57.64 0.28 57.64 0.28 59.32 0.76 59.32 0.76 60.36 0.28 60.36 0.28 62.04 0.76 62.04 0.76 63.08 0.28 63.08 0.28 64.76 0.76 64.76 0.76 65.8 0.28 65.8 0.28 67.48 0.76 67.48 0.76 68.52 0.28 68.52 0.28 70.2 0.76 70.2 0.76 71.24 0.28 71.24 0.28 72.92 0.76 72.92 0.76 73.96 0.28 73.96 0.28 75.64 0.76 75.64 0.76 76.68 0.28 76.68 0.28 78.36 0.76 78.36 0.76 79.4 0.28 79.4 0.28 81.08 ;
      POLYGON 84.36 15.8 84.36 14.12 83.88 14.12 83.88 13.08 84.36 13.08 84.36 11.4 83.88 11.4 83.88 10.36 84.36 10.36 84.36 8.68 83.88 8.68 83.88 7.64 84.36 7.64 84.36 5.96 83.88 5.96 83.88 4.92 84.36 4.92 84.36 3.24 83.88 3.24 83.88 2.2 84.36 2.2 84.36 0.52 18.68 0.52 18.68 2.2 19.16 2.2 19.16 3.24 18.68 3.24 18.68 4.92 19.16 4.92 19.16 5.96 18.68 5.96 18.68 7.64 19.16 7.64 19.16 8.68 18.68 8.68 18.68 10.36 19.16 10.36 19.16 11.4 18.68 11.4 18.68 13.08 19.16 13.08 19.16 14.12 18.68 14.12 18.68 15.8 ;
    LAYER li1 ;
      POLYGON 102.87 81.43 102.87 16.49 84.47 16.49 84.47 0.17 18.57 0.17 18.57 16.49 0.17 16.49 0.17 81.43 ;
    LAYER mcon ;
      RECT 102.725 81.515 102.895 81.685 ;
      RECT 102.265 81.515 102.435 81.685 ;
      RECT 101.805 81.515 101.975 81.685 ;
      RECT 101.345 81.515 101.515 81.685 ;
      RECT 100.885 81.515 101.055 81.685 ;
      RECT 100.425 81.515 100.595 81.685 ;
      RECT 99.965 81.515 100.135 81.685 ;
      RECT 99.505 81.515 99.675 81.685 ;
      RECT 99.045 81.515 99.215 81.685 ;
      RECT 98.585 81.515 98.755 81.685 ;
      RECT 98.125 81.515 98.295 81.685 ;
      RECT 97.665 81.515 97.835 81.685 ;
      RECT 97.205 81.515 97.375 81.685 ;
      RECT 96.745 81.515 96.915 81.685 ;
      RECT 96.285 81.515 96.455 81.685 ;
      RECT 95.825 81.515 95.995 81.685 ;
      RECT 95.365 81.515 95.535 81.685 ;
      RECT 94.905 81.515 95.075 81.685 ;
      RECT 94.445 81.515 94.615 81.685 ;
      RECT 93.985 81.515 94.155 81.685 ;
      RECT 93.525 81.515 93.695 81.685 ;
      RECT 93.065 81.515 93.235 81.685 ;
      RECT 92.605 81.515 92.775 81.685 ;
      RECT 92.145 81.515 92.315 81.685 ;
      RECT 91.685 81.515 91.855 81.685 ;
      RECT 91.225 81.515 91.395 81.685 ;
      RECT 90.765 81.515 90.935 81.685 ;
      RECT 90.305 81.515 90.475 81.685 ;
      RECT 89.845 81.515 90.015 81.685 ;
      RECT 89.385 81.515 89.555 81.685 ;
      RECT 88.925 81.515 89.095 81.685 ;
      RECT 88.465 81.515 88.635 81.685 ;
      RECT 88.005 81.515 88.175 81.685 ;
      RECT 87.545 81.515 87.715 81.685 ;
      RECT 87.085 81.515 87.255 81.685 ;
      RECT 86.625 81.515 86.795 81.685 ;
      RECT 86.165 81.515 86.335 81.685 ;
      RECT 85.705 81.515 85.875 81.685 ;
      RECT 85.245 81.515 85.415 81.685 ;
      RECT 84.785 81.515 84.955 81.685 ;
      RECT 84.325 81.515 84.495 81.685 ;
      RECT 83.865 81.515 84.035 81.685 ;
      RECT 83.405 81.515 83.575 81.685 ;
      RECT 82.945 81.515 83.115 81.685 ;
      RECT 82.485 81.515 82.655 81.685 ;
      RECT 82.025 81.515 82.195 81.685 ;
      RECT 81.565 81.515 81.735 81.685 ;
      RECT 81.105 81.515 81.275 81.685 ;
      RECT 80.645 81.515 80.815 81.685 ;
      RECT 80.185 81.515 80.355 81.685 ;
      RECT 79.725 81.515 79.895 81.685 ;
      RECT 79.265 81.515 79.435 81.685 ;
      RECT 78.805 81.515 78.975 81.685 ;
      RECT 78.345 81.515 78.515 81.685 ;
      RECT 77.885 81.515 78.055 81.685 ;
      RECT 77.425 81.515 77.595 81.685 ;
      RECT 76.965 81.515 77.135 81.685 ;
      RECT 76.505 81.515 76.675 81.685 ;
      RECT 76.045 81.515 76.215 81.685 ;
      RECT 75.585 81.515 75.755 81.685 ;
      RECT 75.125 81.515 75.295 81.685 ;
      RECT 74.665 81.515 74.835 81.685 ;
      RECT 74.205 81.515 74.375 81.685 ;
      RECT 73.745 81.515 73.915 81.685 ;
      RECT 73.285 81.515 73.455 81.685 ;
      RECT 72.825 81.515 72.995 81.685 ;
      RECT 72.365 81.515 72.535 81.685 ;
      RECT 71.905 81.515 72.075 81.685 ;
      RECT 71.445 81.515 71.615 81.685 ;
      RECT 70.985 81.515 71.155 81.685 ;
      RECT 70.525 81.515 70.695 81.685 ;
      RECT 70.065 81.515 70.235 81.685 ;
      RECT 69.605 81.515 69.775 81.685 ;
      RECT 69.145 81.515 69.315 81.685 ;
      RECT 68.685 81.515 68.855 81.685 ;
      RECT 68.225 81.515 68.395 81.685 ;
      RECT 67.765 81.515 67.935 81.685 ;
      RECT 67.305 81.515 67.475 81.685 ;
      RECT 66.845 81.515 67.015 81.685 ;
      RECT 66.385 81.515 66.555 81.685 ;
      RECT 65.925 81.515 66.095 81.685 ;
      RECT 65.465 81.515 65.635 81.685 ;
      RECT 65.005 81.515 65.175 81.685 ;
      RECT 64.545 81.515 64.715 81.685 ;
      RECT 64.085 81.515 64.255 81.685 ;
      RECT 63.625 81.515 63.795 81.685 ;
      RECT 63.165 81.515 63.335 81.685 ;
      RECT 62.705 81.515 62.875 81.685 ;
      RECT 62.245 81.515 62.415 81.685 ;
      RECT 61.785 81.515 61.955 81.685 ;
      RECT 61.325 81.515 61.495 81.685 ;
      RECT 60.865 81.515 61.035 81.685 ;
      RECT 60.405 81.515 60.575 81.685 ;
      RECT 59.945 81.515 60.115 81.685 ;
      RECT 59.485 81.515 59.655 81.685 ;
      RECT 59.025 81.515 59.195 81.685 ;
      RECT 58.565 81.515 58.735 81.685 ;
      RECT 58.105 81.515 58.275 81.685 ;
      RECT 57.645 81.515 57.815 81.685 ;
      RECT 57.185 81.515 57.355 81.685 ;
      RECT 56.725 81.515 56.895 81.685 ;
      RECT 56.265 81.515 56.435 81.685 ;
      RECT 55.805 81.515 55.975 81.685 ;
      RECT 55.345 81.515 55.515 81.685 ;
      RECT 54.885 81.515 55.055 81.685 ;
      RECT 54.425 81.515 54.595 81.685 ;
      RECT 53.965 81.515 54.135 81.685 ;
      RECT 53.505 81.515 53.675 81.685 ;
      RECT 53.045 81.515 53.215 81.685 ;
      RECT 52.585 81.515 52.755 81.685 ;
      RECT 52.125 81.515 52.295 81.685 ;
      RECT 51.665 81.515 51.835 81.685 ;
      RECT 51.205 81.515 51.375 81.685 ;
      RECT 50.745 81.515 50.915 81.685 ;
      RECT 50.285 81.515 50.455 81.685 ;
      RECT 49.825 81.515 49.995 81.685 ;
      RECT 49.365 81.515 49.535 81.685 ;
      RECT 48.905 81.515 49.075 81.685 ;
      RECT 48.445 81.515 48.615 81.685 ;
      RECT 47.985 81.515 48.155 81.685 ;
      RECT 47.525 81.515 47.695 81.685 ;
      RECT 47.065 81.515 47.235 81.685 ;
      RECT 46.605 81.515 46.775 81.685 ;
      RECT 46.145 81.515 46.315 81.685 ;
      RECT 45.685 81.515 45.855 81.685 ;
      RECT 45.225 81.515 45.395 81.685 ;
      RECT 44.765 81.515 44.935 81.685 ;
      RECT 44.305 81.515 44.475 81.685 ;
      RECT 43.845 81.515 44.015 81.685 ;
      RECT 43.385 81.515 43.555 81.685 ;
      RECT 42.925 81.515 43.095 81.685 ;
      RECT 42.465 81.515 42.635 81.685 ;
      RECT 42.005 81.515 42.175 81.685 ;
      RECT 41.545 81.515 41.715 81.685 ;
      RECT 41.085 81.515 41.255 81.685 ;
      RECT 40.625 81.515 40.795 81.685 ;
      RECT 40.165 81.515 40.335 81.685 ;
      RECT 39.705 81.515 39.875 81.685 ;
      RECT 39.245 81.515 39.415 81.685 ;
      RECT 38.785 81.515 38.955 81.685 ;
      RECT 38.325 81.515 38.495 81.685 ;
      RECT 37.865 81.515 38.035 81.685 ;
      RECT 37.405 81.515 37.575 81.685 ;
      RECT 36.945 81.515 37.115 81.685 ;
      RECT 36.485 81.515 36.655 81.685 ;
      RECT 36.025 81.515 36.195 81.685 ;
      RECT 35.565 81.515 35.735 81.685 ;
      RECT 35.105 81.515 35.275 81.685 ;
      RECT 34.645 81.515 34.815 81.685 ;
      RECT 34.185 81.515 34.355 81.685 ;
      RECT 33.725 81.515 33.895 81.685 ;
      RECT 33.265 81.515 33.435 81.685 ;
      RECT 32.805 81.515 32.975 81.685 ;
      RECT 32.345 81.515 32.515 81.685 ;
      RECT 31.885 81.515 32.055 81.685 ;
      RECT 31.425 81.515 31.595 81.685 ;
      RECT 30.965 81.515 31.135 81.685 ;
      RECT 30.505 81.515 30.675 81.685 ;
      RECT 30.045 81.515 30.215 81.685 ;
      RECT 29.585 81.515 29.755 81.685 ;
      RECT 29.125 81.515 29.295 81.685 ;
      RECT 28.665 81.515 28.835 81.685 ;
      RECT 28.205 81.515 28.375 81.685 ;
      RECT 27.745 81.515 27.915 81.685 ;
      RECT 27.285 81.515 27.455 81.685 ;
      RECT 26.825 81.515 26.995 81.685 ;
      RECT 26.365 81.515 26.535 81.685 ;
      RECT 25.905 81.515 26.075 81.685 ;
      RECT 25.445 81.515 25.615 81.685 ;
      RECT 24.985 81.515 25.155 81.685 ;
      RECT 24.525 81.515 24.695 81.685 ;
      RECT 24.065 81.515 24.235 81.685 ;
      RECT 23.605 81.515 23.775 81.685 ;
      RECT 23.145 81.515 23.315 81.685 ;
      RECT 22.685 81.515 22.855 81.685 ;
      RECT 22.225 81.515 22.395 81.685 ;
      RECT 21.765 81.515 21.935 81.685 ;
      RECT 21.305 81.515 21.475 81.685 ;
      RECT 20.845 81.515 21.015 81.685 ;
      RECT 20.385 81.515 20.555 81.685 ;
      RECT 19.925 81.515 20.095 81.685 ;
      RECT 19.465 81.515 19.635 81.685 ;
      RECT 19.005 81.515 19.175 81.685 ;
      RECT 18.545 81.515 18.715 81.685 ;
      RECT 18.085 81.515 18.255 81.685 ;
      RECT 17.625 81.515 17.795 81.685 ;
      RECT 17.165 81.515 17.335 81.685 ;
      RECT 16.705 81.515 16.875 81.685 ;
      RECT 16.245 81.515 16.415 81.685 ;
      RECT 15.785 81.515 15.955 81.685 ;
      RECT 15.325 81.515 15.495 81.685 ;
      RECT 14.865 81.515 15.035 81.685 ;
      RECT 14.405 81.515 14.575 81.685 ;
      RECT 13.945 81.515 14.115 81.685 ;
      RECT 13.485 81.515 13.655 81.685 ;
      RECT 13.025 81.515 13.195 81.685 ;
      RECT 12.565 81.515 12.735 81.685 ;
      RECT 12.105 81.515 12.275 81.685 ;
      RECT 11.645 81.515 11.815 81.685 ;
      RECT 11.185 81.515 11.355 81.685 ;
      RECT 10.725 81.515 10.895 81.685 ;
      RECT 10.265 81.515 10.435 81.685 ;
      RECT 9.805 81.515 9.975 81.685 ;
      RECT 9.345 81.515 9.515 81.685 ;
      RECT 8.885 81.515 9.055 81.685 ;
      RECT 8.425 81.515 8.595 81.685 ;
      RECT 7.965 81.515 8.135 81.685 ;
      RECT 7.505 81.515 7.675 81.685 ;
      RECT 7.045 81.515 7.215 81.685 ;
      RECT 6.585 81.515 6.755 81.685 ;
      RECT 6.125 81.515 6.295 81.685 ;
      RECT 5.665 81.515 5.835 81.685 ;
      RECT 5.205 81.515 5.375 81.685 ;
      RECT 4.745 81.515 4.915 81.685 ;
      RECT 4.285 81.515 4.455 81.685 ;
      RECT 3.825 81.515 3.995 81.685 ;
      RECT 3.365 81.515 3.535 81.685 ;
      RECT 2.905 81.515 3.075 81.685 ;
      RECT 2.445 81.515 2.615 81.685 ;
      RECT 1.985 81.515 2.155 81.685 ;
      RECT 1.525 81.515 1.695 81.685 ;
      RECT 1.065 81.515 1.235 81.685 ;
      RECT 0.605 81.515 0.775 81.685 ;
      RECT 0.145 81.515 0.315 81.685 ;
      RECT 102.725 78.795 102.895 78.965 ;
      RECT 102.265 78.795 102.435 78.965 ;
      RECT 0.605 78.795 0.775 78.965 ;
      RECT 0.145 78.795 0.315 78.965 ;
      RECT 102.725 76.075 102.895 76.245 ;
      RECT 102.265 76.075 102.435 76.245 ;
      RECT 0.605 76.075 0.775 76.245 ;
      RECT 0.145 76.075 0.315 76.245 ;
      RECT 102.725 73.355 102.895 73.525 ;
      RECT 102.265 73.355 102.435 73.525 ;
      RECT 0.605 73.355 0.775 73.525 ;
      RECT 0.145 73.355 0.315 73.525 ;
      RECT 102.725 70.635 102.895 70.805 ;
      RECT 102.265 70.635 102.435 70.805 ;
      RECT 0.605 70.635 0.775 70.805 ;
      RECT 0.145 70.635 0.315 70.805 ;
      RECT 102.725 67.915 102.895 68.085 ;
      RECT 102.265 67.915 102.435 68.085 ;
      RECT 0.605 67.915 0.775 68.085 ;
      RECT 0.145 67.915 0.315 68.085 ;
      RECT 102.725 65.195 102.895 65.365 ;
      RECT 102.265 65.195 102.435 65.365 ;
      RECT 0.605 65.195 0.775 65.365 ;
      RECT 0.145 65.195 0.315 65.365 ;
      RECT 102.725 62.475 102.895 62.645 ;
      RECT 102.265 62.475 102.435 62.645 ;
      RECT 0.605 62.475 0.775 62.645 ;
      RECT 0.145 62.475 0.315 62.645 ;
      RECT 102.725 59.755 102.895 59.925 ;
      RECT 102.265 59.755 102.435 59.925 ;
      RECT 0.605 59.755 0.775 59.925 ;
      RECT 0.145 59.755 0.315 59.925 ;
      RECT 102.725 57.035 102.895 57.205 ;
      RECT 102.265 57.035 102.435 57.205 ;
      RECT 0.605 57.035 0.775 57.205 ;
      RECT 0.145 57.035 0.315 57.205 ;
      RECT 102.725 54.315 102.895 54.485 ;
      RECT 102.265 54.315 102.435 54.485 ;
      RECT 0.605 54.315 0.775 54.485 ;
      RECT 0.145 54.315 0.315 54.485 ;
      RECT 102.725 51.595 102.895 51.765 ;
      RECT 102.265 51.595 102.435 51.765 ;
      RECT 0.605 51.595 0.775 51.765 ;
      RECT 0.145 51.595 0.315 51.765 ;
      RECT 102.725 48.875 102.895 49.045 ;
      RECT 102.265 48.875 102.435 49.045 ;
      RECT 0.605 48.875 0.775 49.045 ;
      RECT 0.145 48.875 0.315 49.045 ;
      RECT 102.725 46.155 102.895 46.325 ;
      RECT 102.265 46.155 102.435 46.325 ;
      RECT 0.605 46.155 0.775 46.325 ;
      RECT 0.145 46.155 0.315 46.325 ;
      RECT 102.725 43.435 102.895 43.605 ;
      RECT 102.265 43.435 102.435 43.605 ;
      RECT 0.605 43.435 0.775 43.605 ;
      RECT 0.145 43.435 0.315 43.605 ;
      RECT 102.725 40.715 102.895 40.885 ;
      RECT 102.265 40.715 102.435 40.885 ;
      RECT 0.605 40.715 0.775 40.885 ;
      RECT 0.145 40.715 0.315 40.885 ;
      RECT 102.725 37.995 102.895 38.165 ;
      RECT 102.265 37.995 102.435 38.165 ;
      RECT 0.605 37.995 0.775 38.165 ;
      RECT 0.145 37.995 0.315 38.165 ;
      RECT 102.725 35.275 102.895 35.445 ;
      RECT 102.265 35.275 102.435 35.445 ;
      RECT 0.605 35.275 0.775 35.445 ;
      RECT 0.145 35.275 0.315 35.445 ;
      RECT 102.725 32.555 102.895 32.725 ;
      RECT 102.265 32.555 102.435 32.725 ;
      RECT 0.605 32.555 0.775 32.725 ;
      RECT 0.145 32.555 0.315 32.725 ;
      RECT 102.725 29.835 102.895 30.005 ;
      RECT 102.265 29.835 102.435 30.005 ;
      RECT 0.605 29.835 0.775 30.005 ;
      RECT 0.145 29.835 0.315 30.005 ;
      RECT 102.725 27.115 102.895 27.285 ;
      RECT 102.265 27.115 102.435 27.285 ;
      RECT 0.605 27.115 0.775 27.285 ;
      RECT 0.145 27.115 0.315 27.285 ;
      RECT 102.725 24.395 102.895 24.565 ;
      RECT 102.265 24.395 102.435 24.565 ;
      RECT 0.605 24.395 0.775 24.565 ;
      RECT 0.145 24.395 0.315 24.565 ;
      RECT 102.725 21.675 102.895 21.845 ;
      RECT 102.265 21.675 102.435 21.845 ;
      RECT 0.605 21.675 0.775 21.845 ;
      RECT 0.145 21.675 0.315 21.845 ;
      RECT 102.725 18.955 102.895 19.125 ;
      RECT 102.265 18.955 102.435 19.125 ;
      RECT 0.605 18.955 0.775 19.125 ;
      RECT 0.145 18.955 0.315 19.125 ;
      RECT 102.725 16.235 102.895 16.405 ;
      RECT 102.265 16.235 102.435 16.405 ;
      RECT 101.805 16.235 101.975 16.405 ;
      RECT 101.345 16.235 101.515 16.405 ;
      RECT 100.885 16.235 101.055 16.405 ;
      RECT 100.425 16.235 100.595 16.405 ;
      RECT 99.965 16.235 100.135 16.405 ;
      RECT 99.505 16.235 99.675 16.405 ;
      RECT 99.045 16.235 99.215 16.405 ;
      RECT 98.585 16.235 98.755 16.405 ;
      RECT 98.125 16.235 98.295 16.405 ;
      RECT 97.665 16.235 97.835 16.405 ;
      RECT 97.205 16.235 97.375 16.405 ;
      RECT 96.745 16.235 96.915 16.405 ;
      RECT 96.285 16.235 96.455 16.405 ;
      RECT 95.825 16.235 95.995 16.405 ;
      RECT 95.365 16.235 95.535 16.405 ;
      RECT 94.905 16.235 95.075 16.405 ;
      RECT 94.445 16.235 94.615 16.405 ;
      RECT 93.985 16.235 94.155 16.405 ;
      RECT 93.525 16.235 93.695 16.405 ;
      RECT 93.065 16.235 93.235 16.405 ;
      RECT 92.605 16.235 92.775 16.405 ;
      RECT 92.145 16.235 92.315 16.405 ;
      RECT 91.685 16.235 91.855 16.405 ;
      RECT 91.225 16.235 91.395 16.405 ;
      RECT 90.765 16.235 90.935 16.405 ;
      RECT 90.305 16.235 90.475 16.405 ;
      RECT 89.845 16.235 90.015 16.405 ;
      RECT 89.385 16.235 89.555 16.405 ;
      RECT 88.925 16.235 89.095 16.405 ;
      RECT 88.465 16.235 88.635 16.405 ;
      RECT 88.005 16.235 88.175 16.405 ;
      RECT 87.545 16.235 87.715 16.405 ;
      RECT 87.085 16.235 87.255 16.405 ;
      RECT 86.625 16.235 86.795 16.405 ;
      RECT 86.165 16.235 86.335 16.405 ;
      RECT 85.705 16.235 85.875 16.405 ;
      RECT 85.245 16.235 85.415 16.405 ;
      RECT 84.785 16.235 84.955 16.405 ;
      RECT 84.325 16.235 84.495 16.405 ;
      RECT 83.865 16.235 84.035 16.405 ;
      RECT 83.405 16.235 83.575 16.405 ;
      RECT 82.945 16.235 83.115 16.405 ;
      RECT 82.485 16.235 82.655 16.405 ;
      RECT 82.025 16.235 82.195 16.405 ;
      RECT 81.565 16.235 81.735 16.405 ;
      RECT 81.105 16.235 81.275 16.405 ;
      RECT 80.645 16.235 80.815 16.405 ;
      RECT 80.185 16.235 80.355 16.405 ;
      RECT 79.725 16.235 79.895 16.405 ;
      RECT 79.265 16.235 79.435 16.405 ;
      RECT 78.805 16.235 78.975 16.405 ;
      RECT 78.345 16.235 78.515 16.405 ;
      RECT 77.885 16.235 78.055 16.405 ;
      RECT 77.425 16.235 77.595 16.405 ;
      RECT 76.965 16.235 77.135 16.405 ;
      RECT 76.505 16.235 76.675 16.405 ;
      RECT 76.045 16.235 76.215 16.405 ;
      RECT 75.585 16.235 75.755 16.405 ;
      RECT 75.125 16.235 75.295 16.405 ;
      RECT 74.665 16.235 74.835 16.405 ;
      RECT 74.205 16.235 74.375 16.405 ;
      RECT 73.745 16.235 73.915 16.405 ;
      RECT 73.285 16.235 73.455 16.405 ;
      RECT 72.825 16.235 72.995 16.405 ;
      RECT 72.365 16.235 72.535 16.405 ;
      RECT 71.905 16.235 72.075 16.405 ;
      RECT 71.445 16.235 71.615 16.405 ;
      RECT 70.985 16.235 71.155 16.405 ;
      RECT 70.525 16.235 70.695 16.405 ;
      RECT 70.065 16.235 70.235 16.405 ;
      RECT 69.605 16.235 69.775 16.405 ;
      RECT 69.145 16.235 69.315 16.405 ;
      RECT 68.685 16.235 68.855 16.405 ;
      RECT 68.225 16.235 68.395 16.405 ;
      RECT 67.765 16.235 67.935 16.405 ;
      RECT 67.305 16.235 67.475 16.405 ;
      RECT 66.845 16.235 67.015 16.405 ;
      RECT 66.385 16.235 66.555 16.405 ;
      RECT 65.925 16.235 66.095 16.405 ;
      RECT 65.465 16.235 65.635 16.405 ;
      RECT 65.005 16.235 65.175 16.405 ;
      RECT 64.545 16.235 64.715 16.405 ;
      RECT 64.085 16.235 64.255 16.405 ;
      RECT 63.625 16.235 63.795 16.405 ;
      RECT 63.165 16.235 63.335 16.405 ;
      RECT 62.705 16.235 62.875 16.405 ;
      RECT 62.245 16.235 62.415 16.405 ;
      RECT 61.785 16.235 61.955 16.405 ;
      RECT 61.325 16.235 61.495 16.405 ;
      RECT 60.865 16.235 61.035 16.405 ;
      RECT 60.405 16.235 60.575 16.405 ;
      RECT 59.945 16.235 60.115 16.405 ;
      RECT 59.485 16.235 59.655 16.405 ;
      RECT 59.025 16.235 59.195 16.405 ;
      RECT 58.565 16.235 58.735 16.405 ;
      RECT 58.105 16.235 58.275 16.405 ;
      RECT 57.645 16.235 57.815 16.405 ;
      RECT 57.185 16.235 57.355 16.405 ;
      RECT 56.725 16.235 56.895 16.405 ;
      RECT 56.265 16.235 56.435 16.405 ;
      RECT 55.805 16.235 55.975 16.405 ;
      RECT 55.345 16.235 55.515 16.405 ;
      RECT 54.885 16.235 55.055 16.405 ;
      RECT 54.425 16.235 54.595 16.405 ;
      RECT 53.965 16.235 54.135 16.405 ;
      RECT 53.505 16.235 53.675 16.405 ;
      RECT 53.045 16.235 53.215 16.405 ;
      RECT 52.585 16.235 52.755 16.405 ;
      RECT 52.125 16.235 52.295 16.405 ;
      RECT 51.665 16.235 51.835 16.405 ;
      RECT 51.205 16.235 51.375 16.405 ;
      RECT 50.745 16.235 50.915 16.405 ;
      RECT 50.285 16.235 50.455 16.405 ;
      RECT 49.825 16.235 49.995 16.405 ;
      RECT 49.365 16.235 49.535 16.405 ;
      RECT 48.905 16.235 49.075 16.405 ;
      RECT 48.445 16.235 48.615 16.405 ;
      RECT 47.985 16.235 48.155 16.405 ;
      RECT 47.525 16.235 47.695 16.405 ;
      RECT 47.065 16.235 47.235 16.405 ;
      RECT 46.605 16.235 46.775 16.405 ;
      RECT 46.145 16.235 46.315 16.405 ;
      RECT 45.685 16.235 45.855 16.405 ;
      RECT 45.225 16.235 45.395 16.405 ;
      RECT 44.765 16.235 44.935 16.405 ;
      RECT 44.305 16.235 44.475 16.405 ;
      RECT 43.845 16.235 44.015 16.405 ;
      RECT 43.385 16.235 43.555 16.405 ;
      RECT 42.925 16.235 43.095 16.405 ;
      RECT 42.465 16.235 42.635 16.405 ;
      RECT 42.005 16.235 42.175 16.405 ;
      RECT 41.545 16.235 41.715 16.405 ;
      RECT 41.085 16.235 41.255 16.405 ;
      RECT 40.625 16.235 40.795 16.405 ;
      RECT 40.165 16.235 40.335 16.405 ;
      RECT 39.705 16.235 39.875 16.405 ;
      RECT 39.245 16.235 39.415 16.405 ;
      RECT 38.785 16.235 38.955 16.405 ;
      RECT 38.325 16.235 38.495 16.405 ;
      RECT 37.865 16.235 38.035 16.405 ;
      RECT 37.405 16.235 37.575 16.405 ;
      RECT 36.945 16.235 37.115 16.405 ;
      RECT 36.485 16.235 36.655 16.405 ;
      RECT 36.025 16.235 36.195 16.405 ;
      RECT 35.565 16.235 35.735 16.405 ;
      RECT 35.105 16.235 35.275 16.405 ;
      RECT 34.645 16.235 34.815 16.405 ;
      RECT 34.185 16.235 34.355 16.405 ;
      RECT 33.725 16.235 33.895 16.405 ;
      RECT 33.265 16.235 33.435 16.405 ;
      RECT 32.805 16.235 32.975 16.405 ;
      RECT 32.345 16.235 32.515 16.405 ;
      RECT 31.885 16.235 32.055 16.405 ;
      RECT 31.425 16.235 31.595 16.405 ;
      RECT 30.965 16.235 31.135 16.405 ;
      RECT 30.505 16.235 30.675 16.405 ;
      RECT 30.045 16.235 30.215 16.405 ;
      RECT 29.585 16.235 29.755 16.405 ;
      RECT 29.125 16.235 29.295 16.405 ;
      RECT 28.665 16.235 28.835 16.405 ;
      RECT 28.205 16.235 28.375 16.405 ;
      RECT 27.745 16.235 27.915 16.405 ;
      RECT 27.285 16.235 27.455 16.405 ;
      RECT 26.825 16.235 26.995 16.405 ;
      RECT 26.365 16.235 26.535 16.405 ;
      RECT 25.905 16.235 26.075 16.405 ;
      RECT 25.445 16.235 25.615 16.405 ;
      RECT 24.985 16.235 25.155 16.405 ;
      RECT 24.525 16.235 24.695 16.405 ;
      RECT 24.065 16.235 24.235 16.405 ;
      RECT 23.605 16.235 23.775 16.405 ;
      RECT 23.145 16.235 23.315 16.405 ;
      RECT 22.685 16.235 22.855 16.405 ;
      RECT 22.225 16.235 22.395 16.405 ;
      RECT 21.765 16.235 21.935 16.405 ;
      RECT 21.305 16.235 21.475 16.405 ;
      RECT 20.845 16.235 21.015 16.405 ;
      RECT 20.385 16.235 20.555 16.405 ;
      RECT 19.925 16.235 20.095 16.405 ;
      RECT 19.465 16.235 19.635 16.405 ;
      RECT 19.005 16.235 19.175 16.405 ;
      RECT 18.545 16.235 18.715 16.405 ;
      RECT 18.085 16.235 18.255 16.405 ;
      RECT 17.625 16.235 17.795 16.405 ;
      RECT 17.165 16.235 17.335 16.405 ;
      RECT 16.705 16.235 16.875 16.405 ;
      RECT 16.245 16.235 16.415 16.405 ;
      RECT 15.785 16.235 15.955 16.405 ;
      RECT 15.325 16.235 15.495 16.405 ;
      RECT 14.865 16.235 15.035 16.405 ;
      RECT 14.405 16.235 14.575 16.405 ;
      RECT 13.945 16.235 14.115 16.405 ;
      RECT 13.485 16.235 13.655 16.405 ;
      RECT 13.025 16.235 13.195 16.405 ;
      RECT 12.565 16.235 12.735 16.405 ;
      RECT 12.105 16.235 12.275 16.405 ;
      RECT 11.645 16.235 11.815 16.405 ;
      RECT 11.185 16.235 11.355 16.405 ;
      RECT 10.725 16.235 10.895 16.405 ;
      RECT 10.265 16.235 10.435 16.405 ;
      RECT 9.805 16.235 9.975 16.405 ;
      RECT 9.345 16.235 9.515 16.405 ;
      RECT 8.885 16.235 9.055 16.405 ;
      RECT 8.425 16.235 8.595 16.405 ;
      RECT 7.965 16.235 8.135 16.405 ;
      RECT 7.505 16.235 7.675 16.405 ;
      RECT 7.045 16.235 7.215 16.405 ;
      RECT 6.585 16.235 6.755 16.405 ;
      RECT 6.125 16.235 6.295 16.405 ;
      RECT 5.665 16.235 5.835 16.405 ;
      RECT 5.205 16.235 5.375 16.405 ;
      RECT 4.745 16.235 4.915 16.405 ;
      RECT 4.285 16.235 4.455 16.405 ;
      RECT 3.825 16.235 3.995 16.405 ;
      RECT 3.365 16.235 3.535 16.405 ;
      RECT 2.905 16.235 3.075 16.405 ;
      RECT 2.445 16.235 2.615 16.405 ;
      RECT 1.985 16.235 2.155 16.405 ;
      RECT 1.525 16.235 1.695 16.405 ;
      RECT 1.065 16.235 1.235 16.405 ;
      RECT 0.605 16.235 0.775 16.405 ;
      RECT 0.145 16.235 0.315 16.405 ;
      RECT 84.325 13.515 84.495 13.685 ;
      RECT 83.865 13.515 84.035 13.685 ;
      RECT 19.005 13.515 19.175 13.685 ;
      RECT 18.545 13.515 18.715 13.685 ;
      RECT 84.325 10.795 84.495 10.965 ;
      RECT 83.865 10.795 84.035 10.965 ;
      RECT 19.005 10.795 19.175 10.965 ;
      RECT 18.545 10.795 18.715 10.965 ;
      RECT 84.325 8.075 84.495 8.245 ;
      RECT 83.865 8.075 84.035 8.245 ;
      RECT 19.005 8.075 19.175 8.245 ;
      RECT 18.545 8.075 18.715 8.245 ;
      RECT 84.325 5.355 84.495 5.525 ;
      RECT 83.865 5.355 84.035 5.525 ;
      RECT 19.005 5.355 19.175 5.525 ;
      RECT 18.545 5.355 18.715 5.525 ;
      RECT 84.325 2.635 84.495 2.805 ;
      RECT 83.865 2.635 84.035 2.805 ;
      RECT 19.005 2.635 19.175 2.805 ;
      RECT 18.545 2.635 18.715 2.805 ;
      RECT 84.325 -0.085 84.495 0.085 ;
      RECT 83.865 -0.085 84.035 0.085 ;
      RECT 83.405 -0.085 83.575 0.085 ;
      RECT 82.945 -0.085 83.115 0.085 ;
      RECT 82.485 -0.085 82.655 0.085 ;
      RECT 82.025 -0.085 82.195 0.085 ;
      RECT 81.565 -0.085 81.735 0.085 ;
      RECT 81.105 -0.085 81.275 0.085 ;
      RECT 80.645 -0.085 80.815 0.085 ;
      RECT 80.185 -0.085 80.355 0.085 ;
      RECT 79.725 -0.085 79.895 0.085 ;
      RECT 79.265 -0.085 79.435 0.085 ;
      RECT 78.805 -0.085 78.975 0.085 ;
      RECT 78.345 -0.085 78.515 0.085 ;
      RECT 77.885 -0.085 78.055 0.085 ;
      RECT 77.425 -0.085 77.595 0.085 ;
      RECT 76.965 -0.085 77.135 0.085 ;
      RECT 76.505 -0.085 76.675 0.085 ;
      RECT 76.045 -0.085 76.215 0.085 ;
      RECT 75.585 -0.085 75.755 0.085 ;
      RECT 75.125 -0.085 75.295 0.085 ;
      RECT 74.665 -0.085 74.835 0.085 ;
      RECT 74.205 -0.085 74.375 0.085 ;
      RECT 73.745 -0.085 73.915 0.085 ;
      RECT 73.285 -0.085 73.455 0.085 ;
      RECT 72.825 -0.085 72.995 0.085 ;
      RECT 72.365 -0.085 72.535 0.085 ;
      RECT 71.905 -0.085 72.075 0.085 ;
      RECT 71.445 -0.085 71.615 0.085 ;
      RECT 70.985 -0.085 71.155 0.085 ;
      RECT 70.525 -0.085 70.695 0.085 ;
      RECT 70.065 -0.085 70.235 0.085 ;
      RECT 69.605 -0.085 69.775 0.085 ;
      RECT 69.145 -0.085 69.315 0.085 ;
      RECT 68.685 -0.085 68.855 0.085 ;
      RECT 68.225 -0.085 68.395 0.085 ;
      RECT 67.765 -0.085 67.935 0.085 ;
      RECT 67.305 -0.085 67.475 0.085 ;
      RECT 66.845 -0.085 67.015 0.085 ;
      RECT 66.385 -0.085 66.555 0.085 ;
      RECT 65.925 -0.085 66.095 0.085 ;
      RECT 65.465 -0.085 65.635 0.085 ;
      RECT 65.005 -0.085 65.175 0.085 ;
      RECT 64.545 -0.085 64.715 0.085 ;
      RECT 64.085 -0.085 64.255 0.085 ;
      RECT 63.625 -0.085 63.795 0.085 ;
      RECT 63.165 -0.085 63.335 0.085 ;
      RECT 62.705 -0.085 62.875 0.085 ;
      RECT 62.245 -0.085 62.415 0.085 ;
      RECT 61.785 -0.085 61.955 0.085 ;
      RECT 61.325 -0.085 61.495 0.085 ;
      RECT 60.865 -0.085 61.035 0.085 ;
      RECT 60.405 -0.085 60.575 0.085 ;
      RECT 59.945 -0.085 60.115 0.085 ;
      RECT 59.485 -0.085 59.655 0.085 ;
      RECT 59.025 -0.085 59.195 0.085 ;
      RECT 58.565 -0.085 58.735 0.085 ;
      RECT 58.105 -0.085 58.275 0.085 ;
      RECT 57.645 -0.085 57.815 0.085 ;
      RECT 57.185 -0.085 57.355 0.085 ;
      RECT 56.725 -0.085 56.895 0.085 ;
      RECT 56.265 -0.085 56.435 0.085 ;
      RECT 55.805 -0.085 55.975 0.085 ;
      RECT 55.345 -0.085 55.515 0.085 ;
      RECT 54.885 -0.085 55.055 0.085 ;
      RECT 54.425 -0.085 54.595 0.085 ;
      RECT 53.965 -0.085 54.135 0.085 ;
      RECT 53.505 -0.085 53.675 0.085 ;
      RECT 53.045 -0.085 53.215 0.085 ;
      RECT 52.585 -0.085 52.755 0.085 ;
      RECT 52.125 -0.085 52.295 0.085 ;
      RECT 51.665 -0.085 51.835 0.085 ;
      RECT 51.205 -0.085 51.375 0.085 ;
      RECT 50.745 -0.085 50.915 0.085 ;
      RECT 50.285 -0.085 50.455 0.085 ;
      RECT 49.825 -0.085 49.995 0.085 ;
      RECT 49.365 -0.085 49.535 0.085 ;
      RECT 48.905 -0.085 49.075 0.085 ;
      RECT 48.445 -0.085 48.615 0.085 ;
      RECT 47.985 -0.085 48.155 0.085 ;
      RECT 47.525 -0.085 47.695 0.085 ;
      RECT 47.065 -0.085 47.235 0.085 ;
      RECT 46.605 -0.085 46.775 0.085 ;
      RECT 46.145 -0.085 46.315 0.085 ;
      RECT 45.685 -0.085 45.855 0.085 ;
      RECT 45.225 -0.085 45.395 0.085 ;
      RECT 44.765 -0.085 44.935 0.085 ;
      RECT 44.305 -0.085 44.475 0.085 ;
      RECT 43.845 -0.085 44.015 0.085 ;
      RECT 43.385 -0.085 43.555 0.085 ;
      RECT 42.925 -0.085 43.095 0.085 ;
      RECT 42.465 -0.085 42.635 0.085 ;
      RECT 42.005 -0.085 42.175 0.085 ;
      RECT 41.545 -0.085 41.715 0.085 ;
      RECT 41.085 -0.085 41.255 0.085 ;
      RECT 40.625 -0.085 40.795 0.085 ;
      RECT 40.165 -0.085 40.335 0.085 ;
      RECT 39.705 -0.085 39.875 0.085 ;
      RECT 39.245 -0.085 39.415 0.085 ;
      RECT 38.785 -0.085 38.955 0.085 ;
      RECT 38.325 -0.085 38.495 0.085 ;
      RECT 37.865 -0.085 38.035 0.085 ;
      RECT 37.405 -0.085 37.575 0.085 ;
      RECT 36.945 -0.085 37.115 0.085 ;
      RECT 36.485 -0.085 36.655 0.085 ;
      RECT 36.025 -0.085 36.195 0.085 ;
      RECT 35.565 -0.085 35.735 0.085 ;
      RECT 35.105 -0.085 35.275 0.085 ;
      RECT 34.645 -0.085 34.815 0.085 ;
      RECT 34.185 -0.085 34.355 0.085 ;
      RECT 33.725 -0.085 33.895 0.085 ;
      RECT 33.265 -0.085 33.435 0.085 ;
      RECT 32.805 -0.085 32.975 0.085 ;
      RECT 32.345 -0.085 32.515 0.085 ;
      RECT 31.885 -0.085 32.055 0.085 ;
      RECT 31.425 -0.085 31.595 0.085 ;
      RECT 30.965 -0.085 31.135 0.085 ;
      RECT 30.505 -0.085 30.675 0.085 ;
      RECT 30.045 -0.085 30.215 0.085 ;
      RECT 29.585 -0.085 29.755 0.085 ;
      RECT 29.125 -0.085 29.295 0.085 ;
      RECT 28.665 -0.085 28.835 0.085 ;
      RECT 28.205 -0.085 28.375 0.085 ;
      RECT 27.745 -0.085 27.915 0.085 ;
      RECT 27.285 -0.085 27.455 0.085 ;
      RECT 26.825 -0.085 26.995 0.085 ;
      RECT 26.365 -0.085 26.535 0.085 ;
      RECT 25.905 -0.085 26.075 0.085 ;
      RECT 25.445 -0.085 25.615 0.085 ;
      RECT 24.985 -0.085 25.155 0.085 ;
      RECT 24.525 -0.085 24.695 0.085 ;
      RECT 24.065 -0.085 24.235 0.085 ;
      RECT 23.605 -0.085 23.775 0.085 ;
      RECT 23.145 -0.085 23.315 0.085 ;
      RECT 22.685 -0.085 22.855 0.085 ;
      RECT 22.225 -0.085 22.395 0.085 ;
      RECT 21.765 -0.085 21.935 0.085 ;
      RECT 21.305 -0.085 21.475 0.085 ;
      RECT 20.845 -0.085 21.015 0.085 ;
      RECT 20.385 -0.085 20.555 0.085 ;
      RECT 19.925 -0.085 20.095 0.085 ;
      RECT 19.465 -0.085 19.635 0.085 ;
      RECT 19.005 -0.085 19.175 0.085 ;
      RECT 18.545 -0.085 18.715 0.085 ;
    LAYER via ;
      RECT 73.525 81.525 73.675 81.675 ;
      RECT 44.085 81.525 44.235 81.675 ;
      RECT 96.525 17.945 96.675 18.095 ;
      RECT 10.505 17.945 10.655 18.095 ;
      RECT 4.525 17.945 4.675 18.095 ;
      RECT 73.525 16.245 73.675 16.395 ;
      RECT 44.085 16.245 44.235 16.395 ;
      RECT 48.685 1.625 48.835 1.775 ;
      RECT 46.845 1.625 46.995 1.775 ;
      RECT 73.525 -0.075 73.675 0.075 ;
      RECT 44.085 -0.075 44.235 0.075 ;
    LAYER via2 ;
      RECT 73.5 81.5 73.7 81.7 ;
      RECT 44.06 81.5 44.26 81.7 ;
      RECT 1.28 77.42 1.48 77.62 ;
      RECT 101.1 66.54 101.3 66.74 ;
      RECT 1.28 57.7 1.48 57.9 ;
      RECT 101.1 52.94 101.3 53.14 ;
      RECT 1.74 46.14 1.94 46.34 ;
      RECT 1.74 39.34 1.94 39.54 ;
      RECT 101.56 31.86 101.76 32.06 ;
      RECT 1.74 31.18 1.94 31.38 ;
      RECT 1.74 25.74 1.94 25.94 ;
      RECT 101.56 24.38 101.76 24.58 ;
      RECT 1.74 24.38 1.94 24.58 ;
      RECT 19.68 12.14 19.88 12.34 ;
      RECT 73.5 -0.1 73.7 0.1 ;
      RECT 44.06 -0.1 44.26 0.1 ;
    LAYER via3 ;
      RECT 73.5 81.5 73.7 81.7 ;
      RECT 44.06 81.5 44.26 81.7 ;
      RECT 101.1 40.7 101.3 40.9 ;
      RECT 20.14 6.7 20.34 6.9 ;
      RECT 73.5 -0.1 73.7 0.1 ;
      RECT 44.06 -0.1 44.26 0.1 ;
    LAYER OVERLAP ;
      POLYGON 18.4 0 18.4 16.32 0 16.32 0 81.6 103.04 81.6 103.04 16.32 84.64 16.32 84.64 0 ;
  END
END sb_1__2_

END LIBRARY
