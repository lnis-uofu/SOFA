VERSION 5.7 ;
BUSBITCHARS "[]" ;

UNITS
  DATABASE MICRONS 1000 ;
END UNITS

MANUFACTURINGGRID 0.005 ;

LAYER li1
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.46 ;
  WIDTH 0.17 ;
END li1

LAYER mcon
  TYPE CUT ;
END mcon

LAYER met1
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.34 ;
  WIDTH 0.14 ;
END met1

LAYER via
  TYPE CUT ;
END via

LAYER met2
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.46 ;
  WIDTH 0.14 ;
END met2

LAYER via2
  TYPE CUT ;
END via2

LAYER met3
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.68 ;
  WIDTH 0.3 ;
END met3

LAYER via3
  TYPE CUT ;
END via3

LAYER met4
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.92 ;
  WIDTH 0.3 ;
END met4

LAYER via4
  TYPE CUT ;
END via4

LAYER met5
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 3.4 ;
  WIDTH 1.6 ;
END met5

LAYER nwell
  TYPE MASTERSLICE ;
END nwell

LAYER pwell
  TYPE MASTERSLICE ;
END pwell

LAYER OVERLAP
  TYPE OVERLAP ;
END OVERLAP

VIA L1M1_PR
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.145 -0.115 0.145 0.115 ;
END L1M1_PR

VIA L1M1_PR_R
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.115 -0.145 0.115 0.145 ;
END L1M1_PR_R

VIA L1M1_PR_M
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.115 -0.145 0.115 0.145 ;
END L1M1_PR_M

VIA L1M1_PR_MR
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.145 -0.115 0.145 0.115 ;
END L1M1_PR_MR

VIA L1M1_PR_C
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.145 -0.145 0.145 0.145 ;
END L1M1_PR_C

VIA M1M2_PR
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR

VIA M1M2_PR_Enc
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_Enc

VIA M1M2_PR_R
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_R

VIA M1M2_PR_R_Enc
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR_R_Enc

VIA M1M2_PR_M
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_M

VIA M1M2_PR_M_Enc
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR_M_Enc

VIA M1M2_PR_MR
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR_MR

VIA M1M2_PR_MR_Enc
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_MR_Enc

VIA M1M2_PR_C
  LAYER met1 ;
    RECT -0.16 -0.16 0.16 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.16 0.16 0.16 ;
END M1M2_PR_C

VIA M2M3_PR
  LAYER met2 ;
    RECT -0.14 -0.185 0.14 0.185 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR

VIA M2M3_PR_R
  LAYER met2 ;
    RECT -0.185 -0.14 0.185 0.14 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_R

VIA M2M3_PR_M
  LAYER met2 ;
    RECT -0.14 -0.185 0.14 0.185 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_M

VIA M2M3_PR_MR
  LAYER met2 ;
    RECT -0.185 -0.14 0.185 0.14 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_MR

VIA M2M3_PR_C
  LAYER met2 ;
    RECT -0.185 -0.185 0.185 0.185 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_C

VIA M3M4_PR
  LAYER met3 ;
    RECT -0.19 -0.16 0.19 0.16 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR

VIA M3M4_PR_R
  LAYER met3 ;
    RECT -0.16 -0.19 0.16 0.19 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_R

VIA M3M4_PR_M
  LAYER met3 ;
    RECT -0.19 -0.16 0.19 0.16 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_M

VIA M3M4_PR_MR
  LAYER met3 ;
    RECT -0.16 -0.19 0.16 0.19 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_MR

VIA M3M4_PR_C
  LAYER met3 ;
    RECT -0.19 -0.19 0.19 0.19 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_C

VIA M4M5_PR
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR

VIA M4M5_PR_R
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_R

VIA M4M5_PR_M
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_M

VIA M4M5_PR_MR
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_MR

VIA M4M5_PR_C
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_C

SITE unit
  CLASS CORE ;
  SYMMETRY Y ;
  SIZE 0.46 BY 2.72 ;
END unit

SITE unithddbl
  CLASS CORE ;
  SIZE 0.46 BY 5.44 ;
END unithddbl

MACRO sb_0__2_
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  SIZE 103.96 BY 87.04 ;
  SYMMETRY X Y ;
  PIN pReset[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.14 86.555 52.28 87.04 ;
    END
  END pReset[0]
  PIN chanx_right_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 103.16 43.03 103.96 43.33 ;
    END
  END chanx_right_in[0]
  PIN chanx_right_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 77.28 103.96 77.42 ;
    END
  END chanx_right_in[1]
  PIN chanx_right_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 61.3 103.96 61.44 ;
    END
  END chanx_right_in[2]
  PIN chanx_right_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 50.42 103.96 50.56 ;
    END
  END chanx_right_in[3]
  PIN chanx_right_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 103.16 55.27 103.96 55.57 ;
    END
  END chanx_right_in[4]
  PIN chanx_right_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 53.48 103.96 53.62 ;
    END
  END chanx_right_in[5]
  PIN chanx_right_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 103.16 56.63 103.96 56.93 ;
    END
  END chanx_right_in[6]
  PIN chanx_right_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 18.12 103.96 18.26 ;
    END
  END chanx_right_in[7]
  PIN chanx_right_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 103.16 36.23 103.96 36.53 ;
    END
  END chanx_right_in[8]
  PIN chanx_right_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 52.46 103.96 52.6 ;
    END
  END chanx_right_in[9]
  PIN chanx_right_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 103.16 32.15 103.96 32.45 ;
    END
  END chanx_right_in[10]
  PIN chanx_right_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 103.16 34.87 103.96 35.17 ;
    END
  END chanx_right_in[11]
  PIN chanx_right_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 36.14 103.96 36.28 ;
    END
  END chanx_right_in[12]
  PIN chanx_right_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 49.74 103.96 49.88 ;
    END
  END chanx_right_in[13]
  PIN chanx_right_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 60.62 103.96 60.76 ;
    END
  END chanx_right_in[14]
  PIN chanx_right_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 103.16 33.51 103.96 33.81 ;
    END
  END chanx_right_in[15]
  PIN chanx_right_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 103.16 53.91 103.96 54.21 ;
    END
  END chanx_right_in[16]
  PIN chanx_right_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 23.56 103.96 23.7 ;
    END
  END chanx_right_in[17]
  PIN chanx_right_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 31.72 103.96 31.86 ;
    END
  END chanx_right_in[18]
  PIN chanx_right_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 55.86 103.96 56 ;
    END
  END chanx_right_in[19]
  PIN chanx_right_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 68.78 103.96 68.92 ;
    END
  END chanx_right_in[20]
  PIN chanx_right_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 37.16 103.96 37.3 ;
    END
  END chanx_right_in[21]
  PIN chanx_right_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 103.16 52.55 103.96 52.85 ;
    END
  END chanx_right_in[22]
  PIN chanx_right_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 33.76 103.96 33.9 ;
    END
  END chanx_right_in[23]
  PIN chanx_right_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 57.9 103.96 58.04 ;
    END
  END chanx_right_in[24]
  PIN chanx_right_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 103.16 45.75 103.96 46.05 ;
    END
  END chanx_right_in[25]
  PIN chanx_right_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 34.44 103.96 34.58 ;
    END
  END chanx_right_in[26]
  PIN chanx_right_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 71.5 103.96 71.64 ;
    END
  END chanx_right_in[27]
  PIN chanx_right_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 41.58 103.96 41.72 ;
    END
  END chanx_right_in[28]
  PIN chanx_right_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 69.46 103.96 69.6 ;
    END
  END chanx_right_in[29]
  PIN right_top_grid_pin_1_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 42.26 103.96 42.4 ;
    END
  END right_top_grid_pin_1_[0]
  PIN right_bottom_grid_pin_36_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.52 10.88 99.66 11.365 ;
    END
  END right_bottom_grid_pin_36_[0]
  PIN right_bottom_grid_pin_37_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 12.68 103.96 12.82 ;
    END
  END right_bottom_grid_pin_37_[0]
  PIN right_bottom_grid_pin_38_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.78 10.88 90.92 11.365 ;
    END
  END right_bottom_grid_pin_38_[0]
  PIN right_bottom_grid_pin_39_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 14.38 103.96 14.52 ;
    END
  END right_bottom_grid_pin_39_[0]
  PIN right_bottom_grid_pin_40_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.54 10.88 93.68 11.365 ;
    END
  END right_bottom_grid_pin_40_[0]
  PIN right_bottom_grid_pin_41_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 73.005 1.8 73.6 1.94 ;
    END
  END right_bottom_grid_pin_41_[0]
  PIN right_bottom_grid_pin_42_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.56 10.88 87.7 11.365 ;
    END
  END right_bottom_grid_pin_42_[0]
  PIN right_bottom_grid_pin_43_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.46 10.88 94.6 11.365 ;
    END
  END right_bottom_grid_pin_43_[0]
  PIN chany_bottom_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.24 0 68.38 0.485 ;
    END
  END chany_bottom_in[0]
  PIN chany_bottom_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.52 0 53.66 0.485 ;
    END
  END chany_bottom_in[1]
  PIN chany_bottom_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.44 0 54.58 0.485 ;
    END
  END chany_bottom_in[2]
  PIN chany_bottom_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 17.79 0 18.09 0.8 ;
    END
  END chany_bottom_in[3]
  PIN chany_bottom_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.64 0 63.78 0.485 ;
    END
  END chany_bottom_in[4]
  PIN chany_bottom_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.96 0 60.1 0.485 ;
    END
  END chany_bottom_in[5]
  PIN chany_bottom_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.52 0 30.66 0.485 ;
    END
  END chany_bottom_in[6]
  PIN chany_bottom_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.48 0 42.62 0.485 ;
    END
  END chany_bottom_in[7]
  PIN chany_bottom_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.96 0 37.1 0.485 ;
    END
  END chany_bottom_in[8]
  PIN chany_bottom_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.36 0 55.5 0.485 ;
    END
  END chany_bottom_in[9]
  PIN chany_bottom_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.68 0 5.82 0.485 ;
    END
  END chany_bottom_in[10]
  PIN chany_bottom_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.2 0 34.34 0.485 ;
    END
  END chany_bottom_in[11]
  PIN chany_bottom_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.76 0 50.9 0.485 ;
    END
  END chany_bottom_in[12]
  PIN chany_bottom_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.12 0 58.26 0.485 ;
    END
  END chany_bottom_in[13]
  PIN chany_bottom_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.56 0 64.7 0.485 ;
    END
  END chany_bottom_in[14]
  PIN chany_bottom_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.54 0 70.68 0.485 ;
    END
  END chany_bottom_in[15]
  PIN chany_bottom_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.62 0 69.76 0.485 ;
    END
  END chany_bottom_in[16]
  PIN chany_bottom_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 19.63 0 19.93 0.8 ;
    END
  END chany_bottom_in[17]
  PIN chany_bottom_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.24 0 45.38 0.485 ;
    END
  END chany_bottom_in[18]
  PIN chany_bottom_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.12 0 12.26 0.485 ;
    END
  END chany_bottom_in[19]
  PIN chany_bottom_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.32 0 44.46 0.485 ;
    END
  END chany_bottom_in[20]
  PIN chany_bottom_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.4 0 66.54 0.485 ;
    END
  END chany_bottom_in[21]
  PIN chany_bottom_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.12 0 35.26 0.485 ;
    END
  END chany_bottom_in[22]
  PIN chany_bottom_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.44 0 8.58 0.485 ;
    END
  END chany_bottom_in[23]
  PIN chany_bottom_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 21.47 0 21.77 0.8 ;
    END
  END chany_bottom_in[24]
  PIN chany_bottom_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.48 0 65.62 0.485 ;
    END
  END chany_bottom_in[25]
  PIN chany_bottom_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.4 0 43.54 0.485 ;
    END
  END chany_bottom_in[26]
  PIN chany_bottom_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.88 0 61.02 0.485 ;
    END
  END chany_bottom_in[27]
  PIN chany_bottom_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.28 0 56.42 0.485 ;
    END
  END chany_bottom_in[28]
  PIN chany_bottom_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.2 0 57.34 0.485 ;
    END
  END chany_bottom_in[29]
  PIN bottom_left_grid_pin_1_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.6 0 52.74 0.485 ;
    END
  END bottom_left_grid_pin_1_[0]
  PIN ccff_head[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 17.44 103.96 17.58 ;
    END
  END ccff_head[0]
  PIN chanx_right_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 103.16 47.11 103.96 47.41 ;
    END
  END chanx_right_out[0]
  PIN chanx_right_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 44.98 103.96 45.12 ;
    END
  END chanx_right_out[1]
  PIN chanx_right_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 47.7 103.96 47.84 ;
    END
  END chanx_right_out[2]
  PIN chanx_right_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 103.16 48.47 103.96 48.77 ;
    END
  END chanx_right_out[3]
  PIN chanx_right_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 103.16 23.99 103.96 24.29 ;
    END
  END chanx_right_out[4]
  PIN chanx_right_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 103.16 38.95 103.96 39.25 ;
    END
  END chanx_right_out[5]
  PIN chanx_right_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 103.16 25.35 103.96 25.65 ;
    END
  END chanx_right_out[6]
  PIN chanx_right_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 103.16 16.51 103.96 16.81 ;
    END
  END chanx_right_out[7]
  PIN chanx_right_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 30.7 103.96 30.84 ;
    END
  END chanx_right_out[8]
  PIN chanx_right_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 38.86 103.96 39 ;
    END
  END chanx_right_out[9]
  PIN chanx_right_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 103.16 26.71 103.96 27.01 ;
    END
  END chanx_right_out[10]
  PIN chanx_right_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 25.94 103.96 26.08 ;
    END
  END chanx_right_out[11]
  PIN chanx_right_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 29 103.96 29.14 ;
    END
  END chanx_right_out[12]
  PIN chanx_right_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 103.16 22.63 103.96 22.93 ;
    END
  END chanx_right_out[13]
  PIN chanx_right_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 103.16 41.67 103.96 41.97 ;
    END
  END chanx_right_out[14]
  PIN chanx_right_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 103.16 40.31 103.96 40.61 ;
    END
  END chanx_right_out[15]
  PIN chanx_right_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 103.16 17.87 103.96 18.17 ;
    END
  END chanx_right_out[16]
  PIN chanx_right_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 28.32 103.96 28.46 ;
    END
  END chanx_right_out[17]
  PIN chanx_right_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 103.16 44.39 103.96 44.69 ;
    END
  END chanx_right_out[18]
  PIN chanx_right_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 103.16 20.59 103.96 20.89 ;
    END
  END chanx_right_out[19]
  PIN chanx_right_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 103.16 28.07 103.96 28.37 ;
    END
  END chanx_right_out[20]
  PIN chanx_right_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 103.16 37.59 103.96 37.89 ;
    END
  END chanx_right_out[21]
  PIN chanx_right_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 44.3 103.96 44.44 ;
    END
  END chanx_right_out[22]
  PIN chanx_right_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 103.16 30.79 103.96 31.09 ;
    END
  END chanx_right_out[23]
  PIN chanx_right_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 103.16 51.19 103.96 51.49 ;
    END
  END chanx_right_out[24]
  PIN chanx_right_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 103.16 49.83 103.96 50.13 ;
    END
  END chanx_right_out[25]
  PIN chanx_right_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 58.58 103.96 58.72 ;
    END
  END chanx_right_out[26]
  PIN chanx_right_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 55.18 103.96 55.32 ;
    END
  END chanx_right_out[27]
  PIN chanx_right_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 103.16 19.23 103.96 19.53 ;
    END
  END chanx_right_out[28]
  PIN chanx_right_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 103.16 29.43 103.96 29.73 ;
    END
  END chanx_right_out[29]
  PIN chany_bottom_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.36 0 9.5 0.485 ;
    END
  END chany_bottom_out[0]
  PIN chany_bottom_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.72 0 62.86 0.485 ;
    END
  END chany_bottom_out[1]
  PIN chany_bottom_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.56 0 41.7 0.485 ;
    END
  END chany_bottom_out[2]
  PIN chany_bottom_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.52 0 7.66 0.485 ;
    END
  END chany_bottom_out[3]
  PIN chany_bottom_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.16 0 23.3 0.485 ;
    END
  END chany_bottom_out[4]
  PIN chany_bottom_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.88 0 38.02 0.485 ;
    END
  END chany_bottom_out[5]
  PIN chany_bottom_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.6 0 6.74 0.485 ;
    END
  END chany_bottom_out[6]
  PIN chany_bottom_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.04 0 13.18 0.485 ;
    END
  END chany_bottom_out[7]
  PIN chany_bottom_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.24 0 22.38 0.485 ;
    END
  END chany_bottom_out[8]
  PIN chany_bottom_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.8 0 61.94 0.485 ;
    END
  END chany_bottom_out[9]
  PIN chany_bottom_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.64 0 40.78 0.485 ;
    END
  END chany_bottom_out[10]
  PIN chany_bottom_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.8 0 38.94 0.485 ;
    END
  END chany_bottom_out[11]
  PIN chany_bottom_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.2 0 11.34 0.485 ;
    END
  END chany_bottom_out[12]
  PIN chany_bottom_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.96 0 14.1 0.485 ;
    END
  END chany_bottom_out[13]
  PIN chany_bottom_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.32 0 67.46 0.485 ;
    END
  END chany_bottom_out[14]
  PIN chany_bottom_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.32 0 21.46 0.485 ;
    END
  END chany_bottom_out[15]
  PIN chany_bottom_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.46 0 2.6 0.485 ;
    END
  END chany_bottom_out[16]
  PIN chany_bottom_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.88 0 15.02 0.485 ;
    END
  END chany_bottom_out[17]
  PIN chany_bottom_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.04 0 36.18 0.485 ;
    END
  END chany_bottom_out[18]
  PIN chany_bottom_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.4 0 20.54 0.485 ;
    END
  END chany_bottom_out[19]
  PIN chany_bottom_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.8 0 15.94 0.485 ;
    END
  END chany_bottom_out[20]
  PIN chany_bottom_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.48 0 19.62 0.485 ;
    END
  END chany_bottom_out[21]
  PIN chany_bottom_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.28 0 10.42 0.485 ;
    END
  END chany_bottom_out[22]
  PIN chany_bottom_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.72 0 16.86 0.485 ;
    END
  END chany_bottom_out[23]
  PIN chany_bottom_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25 0 25.14 0.485 ;
    END
  END chany_bottom_out[24]
  PIN chany_bottom_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.56 0 18.7 0.485 ;
    END
  END chany_bottom_out[25]
  PIN chany_bottom_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.72 0 39.86 0.485 ;
    END
  END chany_bottom_out[26]
  PIN chany_bottom_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.64 0 17.78 0.485 ;
    END
  END chany_bottom_out[27]
  PIN chany_bottom_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.3 0 4.44 0.485 ;
    END
  END chany_bottom_out[28]
  PIN chany_bottom_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.38 0 3.52 0.485 ;
    END
  END chany_bottom_out[29]
  PIN ccff_tail[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.08 0 24.22 0.485 ;
    END
  END ccff_tail[0]
  PIN SC_IN_TOP
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.06 10.88 76.2 11.365 ;
    END
  END SC_IN_TOP
  PIN SC_OUT_BOT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 22.54 103.96 22.68 ;
    END
  END SC_OUT_BOT
  PIN pReset_E_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.365 39.88 103.96 40.02 ;
    END
  END pReset_E_in
  PIN pReset_S_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.68 0 28.82 0.485 ;
    END
  END pReset_S_out
  PIN prog_clk_0_E_in
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER met1 ;
        RECT 103.365 25.26 103.96 25.4 ;
    END
  END prog_clk_0_E_in
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0 26.96 3.2 30.16 ;
        RECT 100.76 26.96 103.96 30.16 ;
        RECT 0 67.76 3.2 70.96 ;
        RECT 100.76 67.76 103.96 70.96 ;
      LAYER met4 ;
        RECT 14.42 0 15.02 0.6 ;
        RECT 43.86 0 44.46 0.6 ;
        RECT 89.86 10.88 90.46 11.48 ;
        RECT 14.42 86.44 15.02 87.04 ;
        RECT 43.86 86.44 44.46 87.04 ;
        RECT 89.86 86.44 90.46 87.04 ;
      LAYER met1 ;
        RECT 0 2.48 0.48 2.96 ;
        RECT 73.12 2.48 73.6 2.96 ;
        RECT 0 7.92 0.48 8.4 ;
        RECT 73.12 7.92 73.6 8.4 ;
        RECT 0 13.36 0.48 13.84 ;
        RECT 103.48 13.36 103.96 13.84 ;
        RECT 0 18.8 0.48 19.28 ;
        RECT 103.48 18.8 103.96 19.28 ;
        RECT 0 24.24 0.48 24.72 ;
        RECT 103.48 24.24 103.96 24.72 ;
        RECT 0 29.68 0.48 30.16 ;
        RECT 103.48 29.68 103.96 30.16 ;
        RECT 0 35.12 0.48 35.6 ;
        RECT 103.48 35.12 103.96 35.6 ;
        RECT 0 40.56 0.48 41.04 ;
        RECT 103.48 40.56 103.96 41.04 ;
        RECT 0 46 0.48 46.48 ;
        RECT 103.48 46 103.96 46.48 ;
        RECT 0 51.44 0.48 51.92 ;
        RECT 103.48 51.44 103.96 51.92 ;
        RECT 0 56.88 0.48 57.36 ;
        RECT 103.48 56.88 103.96 57.36 ;
        RECT 0 62.32 0.48 62.8 ;
        RECT 103.48 62.32 103.96 62.8 ;
        RECT 0 67.76 0.48 68.24 ;
        RECT 103.48 67.76 103.96 68.24 ;
        RECT 0 73.2 0.48 73.68 ;
        RECT 103.48 73.2 103.96 73.68 ;
        RECT 0 78.64 0.48 79.12 ;
        RECT 103.48 78.64 103.96 79.12 ;
        RECT 0 84.08 0.48 84.56 ;
        RECT 103.48 84.08 103.96 84.56 ;
    END
  END VDD
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0 47.36 3.2 50.56 ;
        RECT 100.76 47.36 103.96 50.56 ;
      LAYER met4 ;
        RECT 29.14 0 29.74 0.6 ;
        RECT 58.58 0 59.18 0.6 ;
        RECT 29.14 86.44 29.74 87.04 ;
        RECT 58.58 86.44 59.18 87.04 ;
      LAYER met1 ;
        RECT 0 -0.24 0.48 0.24 ;
        RECT 73.12 -0.24 73.6 0.24 ;
        RECT 0 5.2 0.48 5.68 ;
        RECT 73.12 5.2 73.6 5.68 ;
        RECT 0 10.64 0.48 11.12 ;
        RECT 103.48 10.64 103.96 11.12 ;
        RECT 0 16.08 0.48 16.56 ;
        RECT 103.48 16.08 103.96 16.56 ;
        RECT 0 21.52 0.48 22 ;
        RECT 103.48 21.52 103.96 22 ;
        RECT 0 26.96 0.48 27.44 ;
        RECT 103.48 26.96 103.96 27.44 ;
        RECT 0 32.4 0.48 32.88 ;
        RECT 103.48 32.4 103.96 32.88 ;
        RECT 0 37.84 0.48 38.32 ;
        RECT 103.48 37.84 103.96 38.32 ;
        RECT 0 43.28 0.48 43.76 ;
        RECT 103.48 43.28 103.96 43.76 ;
        RECT 0 48.72 0.48 49.2 ;
        RECT 103.48 48.72 103.96 49.2 ;
        RECT 0 54.16 0.48 54.64 ;
        RECT 103.48 54.16 103.96 54.64 ;
        RECT 0 59.6 0.48 60.08 ;
        RECT 103.48 59.6 103.96 60.08 ;
        RECT 0 65.04 0.48 65.52 ;
        RECT 103.48 65.04 103.96 65.52 ;
        RECT 0 70.48 0.48 70.96 ;
        RECT 103.48 70.48 103.96 70.96 ;
        RECT 0 75.92 0.48 76.4 ;
        RECT 103.48 75.92 103.96 76.4 ;
        RECT 0 81.36 0.48 81.84 ;
        RECT 103.48 81.36 103.96 81.84 ;
        RECT 0 86.8 0.48 87.28 ;
        RECT 103.48 86.8 103.96 87.28 ;
    END
  END VSS
  OBS
    LAYER met2 ;
      RECT 58.74 86.735 59.02 87.105 ;
      RECT 29.3 86.735 29.58 87.105 ;
      POLYGON 35.72 26.25 35.72 0.24 35.76 0.24 35.76 0.1 35.58 0.1 35.58 26.25 ;
      POLYGON 9.96 19.96 9.96 0.1 9.78 0.1 9.78 0.24 9.82 0.24 9.82 19.96 ;
      POLYGON 52.28 17.24 52.28 0.24 52.32 0.24 52.32 0.1 52.14 0.1 52.14 17.24 ;
      POLYGON 44.92 15.88 44.92 0.1 44.74 0.1 44.74 0.24 44.78 0.24 44.78 15.88 ;
      POLYGON 80.8 12.14 80.8 11.405 80.87 11.405 80.87 11.035 80.59 11.035 80.59 11.405 80.66 11.405 80.66 12.14 ;
      POLYGON 62.4 10.61 62.4 0.1 62.22 0.1 62.22 0.24 62.26 0.24 62.26 10.61 ;
      RECT 53.92 0.69 54.18 1.01 ;
      RECT 40.12 0.69 40.38 1.01 ;
      RECT 34.6 0.69 34.86 1.01 ;
      RECT 58.74 -0.065 59.02 0.305 ;
      RECT 29.3 -0.065 29.58 0.305 ;
      POLYGON 103.68 86.76 103.68 11.16 99.94 11.16 99.94 11.645 99.24 11.645 99.24 11.16 94.88 11.16 94.88 11.645 94.18 11.645 94.18 11.16 93.96 11.16 93.96 11.645 93.26 11.645 93.26 11.16 91.2 11.16 91.2 11.645 90.5 11.645 90.5 11.16 87.98 11.16 87.98 11.645 87.28 11.645 87.28 11.16 76.48 11.16 76.48 11.645 75.78 11.645 75.78 11.16 73.32 11.16 73.32 0.28 70.96 0.28 70.96 0.765 70.26 0.765 70.26 0.28 70.04 0.28 70.04 0.765 69.34 0.765 69.34 0.28 68.66 0.28 68.66 0.765 67.96 0.765 67.96 0.28 67.74 0.28 67.74 0.765 67.04 0.765 67.04 0.28 66.82 0.28 66.82 0.765 66.12 0.765 66.12 0.28 65.9 0.28 65.9 0.765 65.2 0.765 65.2 0.28 64.98 0.28 64.98 0.765 64.28 0.765 64.28 0.28 64.06 0.28 64.06 0.765 63.36 0.765 63.36 0.28 63.14 0.28 63.14 0.765 62.44 0.765 62.44 0.28 62.22 0.28 62.22 0.765 61.52 0.765 61.52 0.28 61.3 0.28 61.3 0.765 60.6 0.765 60.6 0.28 60.38 0.28 60.38 0.765 59.68 0.765 59.68 0.28 58.54 0.28 58.54 0.765 57.84 0.765 57.84 0.28 57.62 0.28 57.62 0.765 56.92 0.765 56.92 0.28 56.7 0.28 56.7 0.765 56 0.765 56 0.28 55.78 0.28 55.78 0.765 55.08 0.765 55.08 0.28 54.86 0.28 54.86 0.765 54.16 0.765 54.16 0.28 53.94 0.28 53.94 0.765 53.24 0.765 53.24 0.28 53.02 0.28 53.02 0.765 52.32 0.765 52.32 0.28 51.18 0.28 51.18 0.765 50.48 0.765 50.48 0.28 45.66 0.28 45.66 0.765 44.96 0.765 44.96 0.28 44.74 0.28 44.74 0.765 44.04 0.765 44.04 0.28 43.82 0.28 43.82 0.765 43.12 0.765 43.12 0.28 42.9 0.28 42.9 0.765 42.2 0.765 42.2 0.28 41.98 0.28 41.98 0.765 41.28 0.765 41.28 0.28 41.06 0.28 41.06 0.765 40.36 0.765 40.36 0.28 40.14 0.28 40.14 0.765 39.44 0.765 39.44 0.28 39.22 0.28 39.22 0.765 38.52 0.765 38.52 0.28 38.3 0.28 38.3 0.765 37.6 0.765 37.6 0.28 37.38 0.28 37.38 0.765 36.68 0.765 36.68 0.28 36.46 0.28 36.46 0.765 35.76 0.765 35.76 0.28 35.54 0.28 35.54 0.765 34.84 0.765 34.84 0.28 34.62 0.28 34.62 0.765 33.92 0.765 33.92 0.28 30.94 0.28 30.94 0.765 30.24 0.765 30.24 0.28 29.1 0.28 29.1 0.765 28.4 0.765 28.4 0.28 25.42 0.28 25.42 0.765 24.72 0.765 24.72 0.28 24.5 0.28 24.5 0.765 23.8 0.765 23.8 0.28 23.58 0.28 23.58 0.765 22.88 0.765 22.88 0.28 22.66 0.28 22.66 0.765 21.96 0.765 21.96 0.28 21.74 0.28 21.74 0.765 21.04 0.765 21.04 0.28 20.82 0.28 20.82 0.765 20.12 0.765 20.12 0.28 19.9 0.28 19.9 0.765 19.2 0.765 19.2 0.28 18.98 0.28 18.98 0.765 18.28 0.765 18.28 0.28 18.06 0.28 18.06 0.765 17.36 0.765 17.36 0.28 17.14 0.28 17.14 0.765 16.44 0.765 16.44 0.28 16.22 0.28 16.22 0.765 15.52 0.765 15.52 0.28 15.3 0.28 15.3 0.765 14.6 0.765 14.6 0.28 14.38 0.28 14.38 0.765 13.68 0.765 13.68 0.28 13.46 0.28 13.46 0.765 12.76 0.765 12.76 0.28 12.54 0.28 12.54 0.765 11.84 0.765 11.84 0.28 11.62 0.28 11.62 0.765 10.92 0.765 10.92 0.28 10.7 0.28 10.7 0.765 10 0.765 10 0.28 9.78 0.28 9.78 0.765 9.08 0.765 9.08 0.28 8.86 0.28 8.86 0.765 8.16 0.765 8.16 0.28 7.94 0.28 7.94 0.765 7.24 0.765 7.24 0.28 7.02 0.28 7.02 0.765 6.32 0.765 6.32 0.28 6.1 0.28 6.1 0.765 5.4 0.765 5.4 0.28 4.72 0.28 4.72 0.765 4.02 0.765 4.02 0.28 3.8 0.28 3.8 0.765 3.1 0.765 3.1 0.28 2.88 0.28 2.88 0.765 2.18 0.765 2.18 0.28 0.28 0.28 0.28 86.76 51.86 86.76 51.86 86.275 52.56 86.275 52.56 86.76 ;
    LAYER met3 ;
      POLYGON 59.045 87.085 59.045 87.08 59.26 87.08 59.26 86.76 59.045 86.76 59.045 86.755 58.715 86.755 58.715 86.76 58.5 86.76 58.5 87.08 58.715 87.08 58.715 87.085 ;
      POLYGON 29.605 87.085 29.605 87.08 29.82 87.08 29.82 86.76 29.605 86.76 29.605 86.755 29.275 86.755 29.275 86.76 29.06 86.76 29.06 87.08 29.275 87.08 29.275 87.085 ;
      POLYGON 103.31 33.13 103.31 32.85 102.76 32.85 102.76 32.83 101.74 32.83 101.74 33.13 ;
      POLYGON 102.76 30.41 102.76 30.39 103.31 30.39 103.31 30.11 100.36 30.11 100.36 30.41 ;
      POLYGON 80.895 11.385 80.895 11.055 80.565 11.055 80.565 11.07 64.48 11.07 64.48 11.37 80.565 11.37 80.565 11.385 ;
      POLYGON 63.875 0.505 63.875 0.49 72.03 0.49 72.03 0.5 72.41 0.5 72.41 0.18 72.03 0.18 72.03 0.19 63.875 0.19 63.875 0.175 63.545 0.175 63.545 0.505 ;
      POLYGON 59.045 0.285 59.045 0.28 59.26 0.28 59.26 -0.04 59.045 -0.04 59.045 -0.045 58.715 -0.045 58.715 -0.04 58.5 -0.04 58.5 0.28 58.715 0.28 58.715 0.285 ;
      POLYGON 29.605 0.285 29.605 0.28 29.82 0.28 29.82 -0.04 29.605 -0.04 29.605 -0.045 29.275 -0.045 29.275 -0.04 29.06 -0.04 29.06 0.28 29.275 0.28 29.275 0.285 ;
      POLYGON 103.56 86.64 103.56 57.33 102.76 57.33 102.76 56.23 103.56 56.23 103.56 55.97 102.76 55.97 102.76 54.87 103.56 54.87 103.56 54.61 102.76 54.61 102.76 53.51 103.56 53.51 103.56 53.25 102.76 53.25 102.76 52.15 103.56 52.15 103.56 51.89 102.76 51.89 102.76 50.79 103.56 50.79 103.56 50.53 102.76 50.53 102.76 49.43 103.56 49.43 103.56 49.17 102.76 49.17 102.76 48.07 103.56 48.07 103.56 47.81 102.76 47.81 102.76 46.71 103.56 46.71 103.56 46.45 102.76 46.45 102.76 45.35 103.56 45.35 103.56 45.09 102.76 45.09 102.76 43.99 103.56 43.99 103.56 43.73 102.76 43.73 102.76 42.63 103.56 42.63 103.56 42.37 102.76 42.37 102.76 41.27 103.56 41.27 103.56 41.01 102.76 41.01 102.76 39.91 103.56 39.91 103.56 39.65 102.76 39.65 102.76 38.55 103.56 38.55 103.56 38.29 102.76 38.29 102.76 37.19 103.56 37.19 103.56 36.93 102.76 36.93 102.76 35.83 103.56 35.83 103.56 35.57 102.76 35.57 102.76 34.47 103.56 34.47 103.56 34.21 102.76 34.21 102.76 33.11 103.56 33.11 103.56 32.85 102.76 32.85 102.76 31.75 103.56 31.75 103.56 31.49 102.76 31.49 102.76 30.39 103.56 30.39 103.56 30.13 102.76 30.13 102.76 29.03 103.56 29.03 103.56 28.77 102.76 28.77 102.76 27.67 103.56 27.67 103.56 27.41 102.76 27.41 102.76 26.31 103.56 26.31 103.56 26.05 102.76 26.05 102.76 24.95 103.56 24.95 103.56 24.69 102.76 24.69 102.76 23.59 103.56 23.59 103.56 23.33 102.76 23.33 102.76 22.23 103.56 22.23 103.56 21.29 102.76 21.29 102.76 20.19 103.56 20.19 103.56 19.93 102.76 19.93 102.76 18.83 103.56 18.83 103.56 18.57 102.76 18.57 102.76 17.47 103.56 17.47 103.56 17.21 102.76 17.21 102.76 16.11 103.56 16.11 103.56 11.28 73.2 11.28 73.2 0.4 0.4 0.4 0.4 86.64 ;
    LAYER met1 ;
      POLYGON 103.2 87.28 103.2 86.8 59.04 86.8 59.04 86.79 58.72 86.79 58.72 86.8 29.6 86.8 29.6 86.79 29.28 86.79 29.28 86.8 0.76 86.8 0.76 87.28 ;
      POLYGON 103.435 48.52 103.435 48.12 103.295 48.12 103.295 48.38 94.46 48.38 94.46 48.52 ;
      RECT 69.92 10.64 103.2 11.12 ;
      POLYGON 59.04 0.25 59.04 0.24 72.84 0.24 72.84 -0.24 0.76 -0.24 0.76 0.24 29.28 0.24 29.28 0.25 29.6 0.25 29.6 0.24 58.72 0.24 58.72 0.25 ;
      POLYGON 103.2 86.76 103.2 86.52 103.68 86.52 103.68 84.84 103.2 84.84 103.2 83.8 103.68 83.8 103.68 82.12 103.2 82.12 103.2 81.08 103.68 81.08 103.68 79.4 103.2 79.4 103.2 78.36 103.68 78.36 103.68 77.7 103.085 77.7 103.085 77 103.68 77 103.68 76.68 103.2 76.68 103.2 75.64 103.68 75.64 103.68 73.96 103.2 73.96 103.2 72.92 103.68 72.92 103.68 71.92 103.085 71.92 103.085 71.22 103.2 71.22 103.2 70.2 103.68 70.2 103.68 69.88 103.085 69.88 103.085 68.5 103.2 68.5 103.2 67.48 103.68 67.48 103.68 65.8 103.2 65.8 103.2 64.76 103.68 64.76 103.68 63.08 103.2 63.08 103.2 62.04 103.68 62.04 103.68 61.72 103.085 61.72 103.085 60.34 103.2 60.34 103.2 59.32 103.68 59.32 103.68 59 103.085 59 103.085 57.62 103.2 57.62 103.2 56.6 103.68 56.6 103.68 56.28 103.085 56.28 103.085 54.9 103.2 54.9 103.2 53.9 103.085 53.9 103.085 53.2 103.68 53.2 103.68 52.88 103.085 52.88 103.085 52.18 103.2 52.18 103.2 51.16 103.68 51.16 103.68 50.84 103.085 50.84 103.085 49.46 103.2 49.46 103.2 48.44 103.68 48.44 103.68 48.12 103.085 48.12 103.085 47.42 103.68 47.42 103.68 46.76 103.2 46.76 103.2 45.72 103.68 45.72 103.68 45.4 103.085 45.4 103.085 44.02 103.2 44.02 103.2 43 103.68 43 103.68 42.68 103.085 42.68 103.085 41.3 103.2 41.3 103.2 40.3 103.085 40.3 103.085 39.6 103.68 39.6 103.68 39.28 103.085 39.28 103.085 38.58 103.2 38.58 103.2 37.58 103.085 37.58 103.085 36.88 103.68 36.88 103.68 36.56 103.085 36.56 103.085 35.86 103.2 35.86 103.2 34.86 103.085 34.86 103.085 33.48 103.68 33.48 103.68 33.16 103.2 33.16 103.2 32.14 103.085 32.14 103.085 31.44 103.68 31.44 103.68 31.12 103.085 31.12 103.085 30.42 103.2 30.42 103.2 29.42 103.085 29.42 103.085 28.04 103.68 28.04 103.68 27.72 103.2 27.72 103.2 26.68 103.68 26.68 103.68 26.36 103.085 26.36 103.085 24.98 103.2 24.98 103.2 23.98 103.085 23.98 103.085 23.28 103.68 23.28 103.68 22.96 103.085 22.96 103.085 22.26 103.2 22.26 103.2 21.24 103.68 21.24 103.68 19.56 103.2 19.56 103.2 18.54 103.085 18.54 103.085 17.16 103.68 17.16 103.68 16.84 103.2 16.84 103.2 15.8 103.68 15.8 103.68 14.8 103.085 14.8 103.085 14.1 103.2 14.1 103.2 13.1 103.085 13.1 103.085 12.4 103.68 12.4 103.68 11.4 103.2 11.4 103.2 11.16 73.32 11.16 73.32 8.68 72.84 8.68 72.84 7.64 73.32 7.64 73.32 5.96 72.84 5.96 72.84 4.92 73.32 4.92 73.32 3.24 72.84 3.24 72.84 2.22 72.725 2.22 72.725 1.52 73.32 1.52 73.32 0.52 72.84 0.52 72.84 0.28 0.76 0.28 0.76 0.52 0.28 0.52 0.28 2.2 0.76 2.2 0.76 3.24 0.28 3.24 0.28 4.92 0.76 4.92 0.76 5.96 0.28 5.96 0.28 7.64 0.76 7.64 0.76 8.68 0.28 8.68 0.28 10.36 0.76 10.36 0.76 11.4 0.28 11.4 0.28 13.08 0.76 13.08 0.76 14.12 0.28 14.12 0.28 15.8 0.76 15.8 0.76 16.84 0.28 16.84 0.28 18.52 0.76 18.52 0.76 19.56 0.28 19.56 0.28 21.24 0.76 21.24 0.76 22.28 0.28 22.28 0.28 23.96 0.76 23.96 0.76 25 0.28 25 0.28 26.68 0.76 26.68 0.76 27.72 0.28 27.72 0.28 29.4 0.76 29.4 0.76 30.44 0.28 30.44 0.28 32.12 0.76 32.12 0.76 33.16 0.28 33.16 0.28 34.84 0.76 34.84 0.76 35.88 0.28 35.88 0.28 37.56 0.76 37.56 0.76 38.6 0.28 38.6 0.28 40.28 0.76 40.28 0.76 41.32 0.28 41.32 0.28 43 0.76 43 0.76 44.04 0.28 44.04 0.28 45.72 0.76 45.72 0.76 46.76 0.28 46.76 0.28 48.44 0.76 48.44 0.76 49.48 0.28 49.48 0.28 51.16 0.76 51.16 0.76 52.2 0.28 52.2 0.28 53.88 0.76 53.88 0.76 54.92 0.28 54.92 0.28 56.6 0.76 56.6 0.76 57.64 0.28 57.64 0.28 59.32 0.76 59.32 0.76 60.36 0.28 60.36 0.28 62.04 0.76 62.04 0.76 63.08 0.28 63.08 0.28 64.76 0.76 64.76 0.76 65.8 0.28 65.8 0.28 67.48 0.76 67.48 0.76 68.52 0.28 68.52 0.28 70.2 0.76 70.2 0.76 71.24 0.28 71.24 0.28 72.92 0.76 72.92 0.76 73.96 0.28 73.96 0.28 75.64 0.76 75.64 0.76 76.68 0.28 76.68 0.28 78.36 0.76 78.36 0.76 79.4 0.28 79.4 0.28 81.08 0.76 81.08 0.76 82.12 0.28 82.12 0.28 83.8 0.76 83.8 0.76 84.84 0.28 84.84 0.28 86.52 0.76 86.52 0.76 86.76 ;
    LAYER met4 ;
      POLYGON 73.29 58.97 73.29 8.35 72.37 8.35 72.37 0.505 72.385 0.505 72.385 0.175 72.055 0.175 72.055 0.505 72.07 0.505 72.07 8.65 72.99 8.65 72.99 58.97 ;
      POLYGON 103.56 86.64 103.56 11.28 90.86 11.28 90.86 11.88 89.46 11.88 89.46 11.28 73.2 11.28 73.2 0.4 59.58 0.4 59.58 1 58.18 1 58.18 0.4 44.86 0.4 44.86 1 43.46 1 43.46 0.4 30.14 0.4 30.14 1 28.74 1 28.74 0.4 22.17 0.4 22.17 1.2 21.07 1.2 21.07 0.4 20.33 0.4 20.33 1.2 19.23 1.2 19.23 0.4 18.49 0.4 18.49 1.2 17.39 1.2 17.39 0.4 15.42 0.4 15.42 1 14.02 1 14.02 0.4 0.4 0.4 0.4 86.64 14.02 86.64 14.02 86.04 15.42 86.04 15.42 86.64 28.74 86.64 28.74 86.04 30.14 86.04 30.14 86.64 43.46 86.64 43.46 86.04 44.86 86.04 44.86 86.64 58.18 86.64 58.18 86.04 59.58 86.04 59.58 86.64 89.46 86.64 89.46 86.04 90.86 86.04 90.86 86.64 ;
    LAYER met5 ;
      POLYGON 102.36 85.44 102.36 72.56 99.16 72.56 99.16 66.16 102.36 66.16 102.36 52.16 99.16 52.16 99.16 45.76 102.36 45.76 102.36 31.76 99.16 31.76 99.16 25.36 102.36 25.36 102.36 12.48 72 12.48 72 1.6 1.6 1.6 1.6 25.36 4.8 25.36 4.8 31.76 1.6 31.76 1.6 45.76 4.8 45.76 4.8 52.16 1.6 52.16 1.6 66.16 4.8 66.16 4.8 72.56 1.6 72.56 1.6 85.44 ;
    LAYER li1 ;
      POLYGON 103.96 87.125 103.96 86.955 97.435 86.955 97.435 86.23 97.145 86.23 97.145 86.955 82.255 86.955 82.255 86.23 81.965 86.23 81.965 86.955 67.535 86.955 67.535 86.23 67.245 86.23 67.245 86.955 52.355 86.955 52.355 86.23 52.065 86.23 52.065 86.955 37.635 86.955 37.635 86.23 37.345 86.23 37.345 86.955 22.455 86.955 22.455 86.23 22.165 86.23 22.165 86.955 7.735 86.955 7.735 86.23 7.445 86.23 7.445 86.955 0 86.955 0 87.125 ;
      RECT 103.04 84.235 103.96 84.405 ;
      RECT 0 84.235 3.68 84.405 ;
      RECT 103.04 81.515 103.96 81.685 ;
      RECT 0 81.515 3.68 81.685 ;
      RECT 103.04 78.795 103.96 78.965 ;
      RECT 0 78.795 3.68 78.965 ;
      RECT 103.04 76.075 103.96 76.245 ;
      RECT 0 76.075 3.68 76.245 ;
      RECT 103.04 73.355 103.96 73.525 ;
      RECT 0 73.355 3.68 73.525 ;
      RECT 103.04 70.635 103.96 70.805 ;
      RECT 0 70.635 3.68 70.805 ;
      RECT 103.5 67.915 103.96 68.085 ;
      RECT 0 67.915 3.68 68.085 ;
      RECT 103.04 65.195 103.96 65.365 ;
      RECT 0 65.195 3.68 65.365 ;
      RECT 103.04 62.475 103.96 62.645 ;
      RECT 0 62.475 3.68 62.645 ;
      RECT 103.04 59.755 103.96 59.925 ;
      RECT 0 59.755 3.68 59.925 ;
      RECT 103.04 57.035 103.96 57.205 ;
      RECT 0 57.035 3.68 57.205 ;
      RECT 103.04 54.315 103.96 54.485 ;
      RECT 0 54.315 3.68 54.485 ;
      RECT 103.04 51.595 103.96 51.765 ;
      RECT 0 51.595 3.68 51.765 ;
      RECT 103.04 48.875 103.96 49.045 ;
      RECT 0 48.875 3.68 49.045 ;
      RECT 103.04 46.155 103.96 46.325 ;
      RECT 0 46.155 3.68 46.325 ;
      RECT 103.04 43.435 103.96 43.605 ;
      RECT 0 43.435 3.68 43.605 ;
      RECT 103.04 40.715 103.96 40.885 ;
      RECT 0 40.715 3.68 40.885 ;
      RECT 103.04 37.995 103.96 38.165 ;
      RECT 0 37.995 3.68 38.165 ;
      RECT 103.04 35.275 103.96 35.445 ;
      RECT 0 35.275 3.68 35.445 ;
      RECT 103.04 32.555 103.96 32.725 ;
      RECT 0 32.555 3.68 32.725 ;
      RECT 103.04 29.835 103.96 30.005 ;
      RECT 0 29.835 3.68 30.005 ;
      RECT 103.04 27.115 103.96 27.285 ;
      RECT 0 27.115 3.68 27.285 ;
      RECT 103.04 24.395 103.96 24.565 ;
      RECT 0 24.395 3.68 24.565 ;
      RECT 103.04 21.675 103.96 21.845 ;
      RECT 0 21.675 3.68 21.845 ;
      RECT 103.04 18.955 103.96 19.125 ;
      RECT 0 18.955 1.84 19.125 ;
      RECT 103.04 16.235 103.96 16.405 ;
      RECT 0 16.235 1.84 16.405 ;
      RECT 103.04 13.515 103.96 13.685 ;
      RECT 0 13.515 3.68 13.685 ;
      POLYGON 86.57 11.785 86.57 10.965 87.535 10.965 87.535 11.425 87.84 11.425 87.84 10.965 88.51 10.965 88.51 11.425 88.68 11.425 88.68 10.965 89.35 10.965 89.35 11.425 89.52 11.425 89.52 10.965 90.19 10.965 90.19 11.425 90.36 11.425 90.36 10.965 91.03 10.965 91.03 11.425 91.285 11.425 91.285 10.965 91.975 10.965 91.975 11.445 92.145 11.445 92.145 10.965 92.815 10.965 92.815 11.445 92.985 11.445 92.985 10.965 93.575 10.965 93.575 11.445 93.905 11.445 93.905 10.965 94.415 10.965 94.415 11.445 94.745 11.445 94.745 10.965 95.255 10.965 95.255 11.765 95.585 11.765 95.585 10.965 97.145 10.965 97.145 11.69 97.435 11.69 97.435 10.965 103.96 10.965 103.96 10.795 69.92 10.795 69.92 10.965 74.495 10.965 74.495 11.445 74.665 11.445 74.665 10.965 75.335 10.965 75.335 11.445 75.505 11.445 75.505 10.965 76.095 10.965 76.095 11.445 76.425 11.445 76.425 10.965 76.935 10.965 76.935 11.445 77.265 11.445 77.265 10.965 77.775 10.965 77.775 11.765 78.105 11.765 78.105 10.965 80.82 10.965 80.82 11.785 81.05 11.785 81.05 10.965 81.965 10.965 81.965 11.69 82.255 11.69 82.255 10.965 84.5 10.965 84.5 11.785 84.73 11.785 84.73 10.965 86.34 10.965 86.34 11.785 ;
      RECT 0 10.795 3.68 10.965 ;
      RECT 69.92 8.075 73.6 8.245 ;
      RECT 0 8.075 3.68 8.245 ;
      RECT 72.68 5.355 73.6 5.525 ;
      RECT 0 5.355 3.68 5.525 ;
      RECT 72.68 2.635 73.6 2.805 ;
      RECT 0 2.635 3.68 2.805 ;
      POLYGON 14.225 0.885 14.225 0.085 14.735 0.085 14.735 0.565 15.065 0.565 15.065 0.085 15.575 0.085 15.575 0.565 15.905 0.565 15.905 0.085 16.495 0.085 16.495 0.565 16.665 0.565 16.665 0.085 17.335 0.085 17.335 0.565 17.505 0.565 17.505 0.085 22.165 0.085 22.165 0.81 22.455 0.81 22.455 0.085 26.275 0.085 26.275 0.465 26.605 0.465 26.605 0.085 27.305 0.085 27.305 0.445 27.635 0.445 27.635 0.085 30.235 0.085 30.235 0.545 30.565 0.545 30.565 0.085 32.465 0.085 32.465 0.525 32.655 0.525 32.655 0.085 34.14 0.085 34.14 0.545 34.445 0.545 34.445 0.085 37.345 0.085 37.345 0.81 37.635 0.81 37.635 0.085 43.295 0.085 43.295 0.465 43.625 0.465 43.625 0.085 44.325 0.085 44.325 0.445 44.655 0.445 44.655 0.085 47.255 0.085 47.255 0.545 47.585 0.545 47.585 0.085 49.485 0.085 49.485 0.525 49.675 0.525 49.675 0.085 51.16 0.085 51.16 0.545 51.465 0.545 51.465 0.085 52.065 0.085 52.065 0.81 52.355 0.81 52.355 0.085 56.945 0.085 56.945 0.62 57.455 0.62 57.455 0.085 59.415 0.085 59.415 0.485 59.745 0.485 59.745 0.085 61.245 0.085 61.245 0.465 61.575 0.465 61.575 0.085 63.535 0.085 63.535 0.485 63.865 0.485 63.865 0.085 65.825 0.085 65.825 0.62 66.335 0.62 66.335 0.085 67.245 0.085 67.245 0.81 67.535 0.81 67.535 0.085 73.6 0.085 73.6 -0.085 0 -0.085 0 0.085 3.315 0.085 3.315 0.885 3.645 0.885 3.645 0.085 4.155 0.085 4.155 0.565 4.485 0.565 4.485 0.085 4.995 0.085 4.995 0.565 5.325 0.565 5.325 0.085 5.915 0.085 5.915 0.565 6.085 0.565 6.085 0.085 6.755 0.085 6.755 0.565 6.925 0.565 6.925 0.085 7.445 0.085 7.445 0.81 7.735 0.81 7.735 0.085 13.895 0.085 13.895 0.885 ;
      POLYGON 103.79 86.87 103.79 11.05 73.43 11.05 73.43 0.17 0.17 0.17 0.17 86.87 ;
    LAYER via ;
      RECT 58.805 86.845 58.955 86.995 ;
      RECT 29.365 86.845 29.515 86.995 ;
      RECT 36.955 0.435 37.105 0.585 ;
      RECT 58.805 0.045 58.955 0.195 ;
      RECT 29.365 0.045 29.515 0.195 ;
    LAYER via2 ;
      RECT 58.78 86.82 58.98 87.02 ;
      RECT 29.34 86.82 29.54 87.02 ;
      RECT 80.63 11.12 80.83 11.32 ;
      RECT 63.61 0.24 63.81 0.44 ;
      RECT 58.78 0.02 58.98 0.22 ;
      RECT 29.34 0.02 29.54 0.22 ;
    LAYER via3 ;
      RECT 58.78 86.82 58.98 87.02 ;
      RECT 29.34 86.82 29.54 87.02 ;
      RECT 72.12 0.24 72.32 0.44 ;
      RECT 58.78 0.02 58.98 0.22 ;
      RECT 29.34 0.02 29.54 0.22 ;
    LAYER OVERLAP ;
      POLYGON 0 0 0 87.04 103.96 87.04 103.96 10.88 73.6 10.88 73.6 0 ;
  END
END sb_0__2_

END LIBRARY
