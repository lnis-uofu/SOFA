//Generated from netlist by SpyDrNet
//netlist name: FPGA88_SOFA_A
module direct_interc
(
    in,
    out
);

    input in;
    output out;

    wire in;
    wire out;

assign out = in;
endmodule

