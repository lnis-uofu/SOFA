VERSION 5.7 ;
BUSBITCHARS "[]" ;

UNITS
  DATABASE MICRONS 1000 ;
END UNITS

MANUFACTURINGGRID 0.005 ;

LAYER nwell
  TYPE MASTERSLICE ;
END nwell

LAYER pwell
  TYPE MASTERSLICE ;
END pwell

LAYER fieldpoly
  TYPE MASTERSLICE ;
END fieldpoly

LAYER li1
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.46 ;
  WIDTH 0.17 ;
END li1

LAYER mcon
  TYPE CUT ;
END mcon

LAYER met1
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.34 ;
  WIDTH 0.14 ;
END met1

LAYER via
  TYPE CUT ;
END via

LAYER met2
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.46 ;
  WIDTH 0.14 ;
END met2

LAYER via2
  TYPE CUT ;
END via2

LAYER met3
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.68 ;
  WIDTH 0.3 ;
END met3

LAYER via3
  TYPE CUT ;
END via3

LAYER met4
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.92 ;
  WIDTH 0.3 ;
END met4

LAYER via4
  TYPE CUT ;
END via4

LAYER met5
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 3.4 ;
  WIDTH 1.6 ;
END met5

LAYER diff
  TYPE MASTERSLICE ;
END diff

LAYER licon1
  TYPE MASTERSLICE ;
END licon1

LAYER OVERLAP
  TYPE OVERLAP ;
END OVERLAP

VIA L1M1_PR
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.145 -0.115 0.145 0.115 ;
END L1M1_PR

VIA L1M1_PR_R
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.115 -0.145 0.115 0.145 ;
END L1M1_PR_R

VIA L1M1_PR_M
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.115 -0.145 0.115 0.145 ;
END L1M1_PR_M

VIA L1M1_PR_MR
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.145 -0.115 0.145 0.115 ;
END L1M1_PR_MR

VIA L1M1_PR_C
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.145 -0.145 0.145 0.145 ;
END L1M1_PR_C

VIA M1M2_PR
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR

VIA M1M2_PR_Enc
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_Enc

VIA M1M2_PR_R
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_R

VIA M1M2_PR_R_Enc
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR_R_Enc

VIA M1M2_PR_M
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_M

VIA M1M2_PR_M_Enc
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR_M_Enc

VIA M1M2_PR_MR
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR_MR

VIA M1M2_PR_MR_Enc
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_MR_Enc

VIA M1M2_PR_C
  LAYER met1 ;
    RECT -0.16 -0.16 0.16 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.16 0.16 0.16 ;
END M1M2_PR_C

VIA M2M3_PR
  LAYER met2 ;
    RECT -0.14 -0.185 0.14 0.185 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR

VIA M2M3_PR_R
  LAYER met2 ;
    RECT -0.185 -0.14 0.185 0.14 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_R

VIA M2M3_PR_M
  LAYER met2 ;
    RECT -0.14 -0.185 0.14 0.185 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_M

VIA M2M3_PR_MR
  LAYER met2 ;
    RECT -0.185 -0.14 0.185 0.14 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_MR

VIA M2M3_PR_C
  LAYER met2 ;
    RECT -0.185 -0.185 0.185 0.185 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_C

VIA M3M4_PR
  LAYER met3 ;
    RECT -0.19 -0.16 0.19 0.16 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR

VIA M3M4_PR_R
  LAYER met3 ;
    RECT -0.16 -0.19 0.16 0.19 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_R

VIA M3M4_PR_M
  LAYER met3 ;
    RECT -0.19 -0.16 0.19 0.16 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_M

VIA M3M4_PR_MR
  LAYER met3 ;
    RECT -0.16 -0.19 0.16 0.19 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_MR

VIA M3M4_PR_C
  LAYER met3 ;
    RECT -0.19 -0.19 0.19 0.19 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_C

VIA M4M5_PR
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR

VIA M4M5_PR_R
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_R

VIA M4M5_PR_M
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_M

VIA M4M5_PR_MR
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_MR

VIA M4M5_PR_C
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_C

SITE unit
  CLASS CORE ;
  SYMMETRY Y ;
  SIZE 0.46 BY 2.72 ;
END unit

SITE unithddbl
  CLASS CORE ;
  SIZE 0.46 BY 5.44 ;
END unithddbl

MACRO sb_1__0_
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  SIZE 141.68 BY 103.36 ;
  SYMMETRY X Y ;
  PIN prog_clk[0]
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER met2 ;
        RECT 30.75 102 30.89 103.36 ;
    END
  END prog_clk[0]
  PIN chany_top_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.43 102 80.57 103.36 ;
    END
  END chany_top_in[0]
  PIN chany_top_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.43 102 57.57 103.36 ;
    END
  END chany_top_in[1]
  PIN chany_top_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.27 102 82.41 103.36 ;
    END
  END chany_top_in[2]
  PIN chany_top_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.99 102 74.13 103.36 ;
    END
  END chany_top_in[3]
  PIN chany_top_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.91 102 52.05 103.36 ;
    END
  END chany_top_in[4]
  PIN chany_top_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.19 102 60.33 103.36 ;
    END
  END chany_top_in[5]
  PIN chany_top_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.91 102 75.05 103.36 ;
    END
  END chany_top_in[6]
  PIN chany_top_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.63 102 66.77 103.36 ;
    END
  END chany_top_in[7]
  PIN chany_top_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.15 102 72.29 103.36 ;
    END
  END chany_top_in[8]
  PIN chany_top_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.55 102 67.69 103.36 ;
    END
  END chany_top_in[9]
  PIN chany_top_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.07 102 73.21 103.36 ;
    END
  END chany_top_in[10]
  PIN chany_top_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.83 102 75.97 103.36 ;
    END
  END chany_top_in[11]
  PIN chany_top_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.83 102 52.97 103.36 ;
    END
  END chany_top_in[12]
  PIN chany_top_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.41 102 63.55 103.36 ;
    END
  END chany_top_in[13]
  PIN chany_top_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.67 102 54.81 103.36 ;
    END
  END chany_top_in[14]
  PIN chany_top_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.75 102 53.89 103.36 ;
    END
  END chany_top_in[15]
  PIN chany_top_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.39 102 69.53 103.36 ;
    END
  END chany_top_in[16]
  PIN chany_top_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.35 102 81.49 103.36 ;
    END
  END chany_top_in[17]
  PIN chany_top_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.57 102 84.71 103.36 ;
    END
  END chany_top_in[18]
  PIN chany_top_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.27 102 59.41 103.36 ;
    END
  END chany_top_in[19]
  PIN top_left_grid_pin_34_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.05 102 33.19 103.36 ;
    END
  END top_left_grid_pin_34_[0]
  PIN top_left_grid_pin_35_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 32.97 102 33.27 103.36 ;
    END
  END top_left_grid_pin_35_[0]
  PIN top_left_grid_pin_36_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 28.52 99.81 29.9 100.11 ;
    END
  END top_left_grid_pin_36_[0]
  PIN top_left_grid_pin_37_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.13 102 32.27 103.36 ;
    END
  END top_left_grid_pin_37_[0]
  PIN top_left_grid_pin_38_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 28.52 97.77 29.9 98.07 ;
    END
  END top_left_grid_pin_38_[0]
  PIN top_left_grid_pin_39_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 28.52 96.41 29.9 96.71 ;
    END
  END top_left_grid_pin_39_[0]
  PIN top_left_grid_pin_40_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 28.52 95.05 29.9 95.35 ;
    END
  END top_left_grid_pin_40_[0]
  PIN top_left_grid_pin_41_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 28.52 90.29 29.9 90.59 ;
    END
  END top_left_grid_pin_41_[0]
  PIN chanx_right_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 140.3 46.09 141.68 46.39 ;
    END
  END chanx_right_in[0]
  PIN chanx_right_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 140.3 16.17 141.68 16.47 ;
    END
  END chanx_right_in[1]
  PIN chanx_right_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 140.3 12.09 141.68 12.39 ;
    END
  END chanx_right_in[2]
  PIN chanx_right_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 140.3 8.01 141.68 8.31 ;
    END
  END chanx_right_in[3]
  PIN chanx_right_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 140.3 13.45 141.68 13.75 ;
    END
  END chanx_right_in[4]
  PIN chanx_right_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 140.3 9.37 141.68 9.67 ;
    END
  END chanx_right_in[5]
  PIN chanx_right_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 140.3 31.13 141.68 31.43 ;
    END
  END chanx_right_in[6]
  PIN chanx_right_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 140.3 47.45 141.68 47.75 ;
    END
  END chanx_right_in[7]
  PIN chanx_right_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 140.3 14.81 141.68 15.11 ;
    END
  END chanx_right_in[8]
  PIN chanx_right_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 140.3 71.93 141.68 72.23 ;
    END
  END chanx_right_in[9]
  PIN chanx_right_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 140.3 25.69 141.68 25.99 ;
    END
  END chanx_right_in[10]
  PIN chanx_right_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 140.3 29.77 141.68 30.07 ;
    END
  END chanx_right_in[11]
  PIN chanx_right_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 140.3 18.89 141.68 19.19 ;
    END
  END chanx_right_in[12]
  PIN chanx_right_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 140.3 44.73 141.68 45.03 ;
    END
  END chanx_right_in[13]
  PIN chanx_right_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 140.3 17.53 141.68 17.83 ;
    END
  END chanx_right_in[14]
  PIN chanx_right_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 140.3 42.01 141.68 42.31 ;
    END
  END chanx_right_in[15]
  PIN chanx_right_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 140.3 3.93 141.68 4.23 ;
    END
  END chanx_right_in[16]
  PIN chanx_right_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 140.3 63.77 141.68 64.07 ;
    END
  END chanx_right_in[17]
  PIN chanx_right_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 140.3 50.17 141.68 50.47 ;
    END
  END chanx_right_in[18]
  PIN chanx_right_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 140.3 58.33 141.68 58.63 ;
    END
  END chanx_right_in[19]
  PIN right_top_grid_pin_42_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.39 74.8 138.53 76.16 ;
    END
  END right_top_grid_pin_42_[0]
  PIN right_top_grid_pin_43_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.78 99.13 113.16 99.43 ;
    END
  END right_top_grid_pin_43_[0]
  PIN right_top_grid_pin_44_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.31 74.8 139.45 76.16 ;
    END
  END right_top_grid_pin_44_[0]
  PIN right_top_grid_pin_45_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.47 74.8 137.61 76.16 ;
    END
  END right_top_grid_pin_45_[0]
  PIN right_top_grid_pin_46_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.78 91.65 113.16 91.95 ;
    END
  END right_top_grid_pin_46_[0]
  PIN right_top_grid_pin_47_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.78 90.29 113.16 90.59 ;
    END
  END right_top_grid_pin_47_[0]
  PIN right_top_grid_pin_48_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.63 74.8 135.77 76.16 ;
    END
  END right_top_grid_pin_48_[0]
  PIN right_top_grid_pin_49_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 136.55 74.8 136.69 76.16 ;
    END
  END right_top_grid_pin_49_[0]
  PIN right_bottom_grid_pin_1_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.31 0 139.45 1.36 ;
    END
  END right_bottom_grid_pin_1_[0]
  PIN chanx_left_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 67.17 1.38 67.47 ;
    END
  END chanx_left_in[0]
  PIN chanx_left_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 54.25 1.38 54.55 ;
    END
  END chanx_left_in[1]
  PIN chanx_left_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 51.53 1.38 51.83 ;
    END
  END chanx_left_in[2]
  PIN chanx_left_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 52.89 1.38 53.19 ;
    END
  END chanx_left_in[3]
  PIN chanx_left_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 62.41 1.38 62.71 ;
    END
  END chanx_left_in[4]
  PIN chanx_left_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 50.17 1.38 50.47 ;
    END
  END chanx_left_in[5]
  PIN chanx_left_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 47.45 1.38 47.75 ;
    END
  END chanx_left_in[6]
  PIN chanx_left_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 70.57 1.38 70.87 ;
    END
  END chanx_left_in[7]
  PIN chanx_left_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 32.49 1.38 32.79 ;
    END
  END chanx_left_in[8]
  PIN chanx_left_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 71.93 1.38 72.23 ;
    END
  END chanx_left_in[9]
  PIN chanx_left_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 56.97 1.38 57.27 ;
    END
  END chanx_left_in[10]
  PIN chanx_left_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 69.21 1.38 69.51 ;
    END
  END chanx_left_in[11]
  PIN chanx_left_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 36.57 1.38 36.87 ;
    END
  END chanx_left_in[12]
  PIN chanx_left_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 44.73 1.38 45.03 ;
    END
  END chanx_left_in[13]
  PIN chanx_left_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 6.65 1.38 6.95 ;
    END
  END chanx_left_in[14]
  PIN chanx_left_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 42.01 1.38 42.31 ;
    END
  END chanx_left_in[15]
  PIN chanx_left_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 28.41 1.38 28.71 ;
    END
  END chanx_left_in[16]
  PIN chanx_left_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 18.89 1.38 19.19 ;
    END
  END chanx_left_in[17]
  PIN chanx_left_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 5.29 1.38 5.59 ;
    END
  END chanx_left_in[18]
  PIN chanx_left_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 3.93 1.38 4.23 ;
    END
  END chanx_left_in[19]
  PIN left_top_grid_pin_42_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.29 74.8 7.43 76.16 ;
    END
  END left_top_grid_pin_42_[0]
  PIN left_top_grid_pin_43_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 28.52 91.65 29.9 91.95 ;
    END
  END left_top_grid_pin_43_[0]
  PIN left_top_grid_pin_44_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.07 74.8 4.21 76.16 ;
    END
  END left_top_grid_pin_44_[0]
  PIN left_top_grid_pin_45_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.99 74.8 5.13 76.16 ;
    END
  END left_top_grid_pin_45_[0]
  PIN left_top_grid_pin_46_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.23 74.8 2.37 76.16 ;
    END
  END left_top_grid_pin_46_[0]
  PIN left_top_grid_pin_47_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.15 74.8 3.29 76.16 ;
    END
  END left_top_grid_pin_47_[0]
  PIN left_top_grid_pin_48_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.43 74.8 11.57 76.16 ;
    END
  END left_top_grid_pin_48_[0]
  PIN left_top_grid_pin_49_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.51 74.8 10.65 76.16 ;
    END
  END left_top_grid_pin_49_[0]
  PIN left_bottom_grid_pin_1_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.23 0 2.37 1.36 ;
    END
  END left_bottom_grid_pin_1_[0]
  PIN ccff_head[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.39 0 138.53 1.36 ;
    END
  END ccff_head[0]
  PIN chany_top_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.75 102 76.89 103.36 ;
    END
  END chany_top_out[0]
  PIN chany_top_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.11 102 61.25 103.36 ;
    END
  END chany_top_out[1]
  PIN chany_top_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.67 102 77.81 103.36 ;
    END
  END chany_top_out[2]
  PIN chany_top_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.23 102 71.37 103.36 ;
    END
  END chany_top_out[3]
  PIN chany_top_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.83 102 98.97 103.36 ;
    END
  END chany_top_out[4]
  PIN chany_top_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.65 102 83.79 103.36 ;
    END
  END chany_top_out[5]
  PIN chany_top_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.31 102 70.45 103.36 ;
    END
  END chany_top_out[6]
  PIN chany_top_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.07 102 50.21 103.36 ;
    END
  END chany_top_out[7]
  PIN chany_top_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.47 102 68.61 103.36 ;
    END
  END chany_top_out[8]
  PIN chany_top_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.35 102 58.49 103.36 ;
    END
  END chany_top_out[9]
  PIN chany_top_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.53 102 96.67 103.36 ;
    END
  END chany_top_out[10]
  PIN chany_top_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.77 102 93.91 103.36 ;
    END
  END chany_top_out[11]
  PIN chany_top_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.51 102 79.65 103.36 ;
    END
  END chany_top_out[12]
  PIN chany_top_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.33 102 64.47 103.36 ;
    END
  END chany_top_out[13]
  PIN chany_top_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.45 102 97.59 103.36 ;
    END
  END chany_top_out[14]
  PIN chany_top_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.99 102 51.13 103.36 ;
    END
  END chany_top_out[15]
  PIN chany_top_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.87 102 87.01 103.36 ;
    END
  END chany_top_out[16]
  PIN chany_top_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.03 102 62.17 103.36 ;
    END
  END chany_top_out[17]
  PIN chany_top_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.61 102 95.75 103.36 ;
    END
  END chany_top_out[18]
  PIN chany_top_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.59 102 78.73 103.36 ;
    END
  END chany_top_out[19]
  PIN chanx_right_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 140.3 59.69 141.68 59.99 ;
    END
  END chanx_right_out[0]
  PIN chanx_right_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 140.3 66.49 141.68 66.79 ;
    END
  END chanx_right_out[1]
  PIN chanx_right_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 140.3 6.65 141.68 6.95 ;
    END
  END chanx_right_out[2]
  PIN chanx_right_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 140.3 67.85 141.68 68.15 ;
    END
  END chanx_right_out[3]
  PIN chanx_right_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 140.3 35.21 141.68 35.51 ;
    END
  END chanx_right_out[4]
  PIN chanx_right_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 140.3 56.97 141.68 57.27 ;
    END
  END chanx_right_out[5]
  PIN chanx_right_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 140.3 28.41 141.68 28.71 ;
    END
  END chanx_right_out[6]
  PIN chanx_right_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 140.3 51.53 141.68 51.83 ;
    END
  END chanx_right_out[7]
  PIN chanx_right_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 140.3 33.85 141.68 34.15 ;
    END
  END chanx_right_out[8]
  PIN chanx_right_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 140.3 40.65 141.68 40.95 ;
    END
  END chanx_right_out[9]
  PIN chanx_right_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 140.3 24.33 141.68 24.63 ;
    END
  END chanx_right_out[10]
  PIN chanx_right_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 140.3 55.61 141.68 55.91 ;
    END
  END chanx_right_out[11]
  PIN chanx_right_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 140.3 69.21 141.68 69.51 ;
    END
  END chanx_right_out[12]
  PIN chanx_right_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 140.3 61.05 141.68 61.35 ;
    END
  END chanx_right_out[13]
  PIN chanx_right_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 140.3 22.97 141.68 23.27 ;
    END
  END chanx_right_out[14]
  PIN chanx_right_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 140.3 39.29 141.68 39.59 ;
    END
  END chanx_right_out[15]
  PIN chanx_right_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 140.3 36.57 141.68 36.87 ;
    END
  END chanx_right_out[16]
  PIN chanx_right_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 140.3 62.41 141.68 62.71 ;
    END
  END chanx_right_out[17]
  PIN chanx_right_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 140.3 20.25 141.68 20.55 ;
    END
  END chanx_right_out[18]
  PIN chanx_right_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 140.3 52.89 141.68 53.19 ;
    END
  END chanx_right_out[19]
  PIN chanx_left_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 27.05 1.38 27.35 ;
    END
  END chanx_left_out[0]
  PIN chanx_left_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 64.45 1.38 64.75 ;
    END
  END chanx_left_out[1]
  PIN chanx_left_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 15.49 1.38 15.79 ;
    END
  END chanx_left_out[2]
  PIN chanx_left_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 59.69 1.38 59.99 ;
    END
  END chanx_left_out[3]
  PIN chanx_left_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 11.41 1.38 11.71 ;
    END
  END chanx_left_out[4]
  PIN chanx_left_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 61.05 1.38 61.35 ;
    END
  END chanx_left_out[5]
  PIN chanx_left_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 25.69 1.38 25.99 ;
    END
  END chanx_left_out[6]
  PIN chanx_left_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 48.81 1.38 49.11 ;
    END
  END chanx_left_out[7]
  PIN chanx_left_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 21.61 1.38 21.91 ;
    END
  END chanx_left_out[8]
  PIN chanx_left_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 33.85 1.38 34.15 ;
    END
  END chanx_left_out[9]
  PIN chanx_left_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 20.25 1.38 20.55 ;
    END
  END chanx_left_out[10]
  PIN chanx_left_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 37.93 1.38 38.23 ;
    END
  END chanx_left_out[11]
  PIN chanx_left_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 22.97 1.38 23.27 ;
    END
  END chanx_left_out[12]
  PIN chanx_left_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 65.81 1.38 66.11 ;
    END
  END chanx_left_out[13]
  PIN chanx_left_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 17.53 1.38 17.83 ;
    END
  END chanx_left_out[14]
  PIN chanx_left_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 39.29 1.38 39.59 ;
    END
  END chanx_left_out[15]
  PIN chanx_left_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 31.13 1.38 31.43 ;
    END
  END chanx_left_out[16]
  PIN chanx_left_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 43.37 1.38 43.67 ;
    END
  END chanx_left_out[17]
  PIN chanx_left_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 10.05 1.38 10.35 ;
    END
  END chanx_left_out[18]
  PIN chanx_left_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 58.33 1.38 58.63 ;
    END
  END chanx_left_out[19]
  PIN ccff_tail[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 55.61 1.38 55.91 ;
    END
  END ccff_tail[0]
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 0.48 2.96 ;
        RECT 141.2 2.48 141.68 2.96 ;
        RECT 0 7.92 0.48 8.4 ;
        RECT 141.2 7.92 141.68 8.4 ;
        RECT 0 13.36 0.48 13.84 ;
        RECT 141.2 13.36 141.68 13.84 ;
        RECT 0 18.8 0.48 19.28 ;
        RECT 141.2 18.8 141.68 19.28 ;
        RECT 0 24.24 0.48 24.72 ;
        RECT 141.2 24.24 141.68 24.72 ;
        RECT 0 29.68 0.48 30.16 ;
        RECT 141.2 29.68 141.68 30.16 ;
        RECT 0 35.12 0.48 35.6 ;
        RECT 141.2 35.12 141.68 35.6 ;
        RECT 0 40.56 0.48 41.04 ;
        RECT 141.2 40.56 141.68 41.04 ;
        RECT 0 46 0.48 46.48 ;
        RECT 141.2 46 141.68 46.48 ;
        RECT 0 51.44 0.48 51.92 ;
        RECT 141.2 51.44 141.68 51.92 ;
        RECT 0 56.88 0.48 57.36 ;
        RECT 141.2 56.88 141.68 57.36 ;
        RECT 0 62.32 0.48 62.8 ;
        RECT 141.2 62.32 141.68 62.8 ;
        RECT 0 67.76 0.48 68.24 ;
        RECT 141.2 67.76 141.68 68.24 ;
        RECT 0 73.2 0.48 73.68 ;
        RECT 141.2 73.2 141.68 73.68 ;
        RECT 28.52 78.64 29 79.12 ;
        RECT 112.68 78.64 113.16 79.12 ;
        RECT 28.52 84.08 29 84.56 ;
        RECT 112.68 84.08 113.16 84.56 ;
        RECT 28.52 89.52 29 90 ;
        RECT 112.68 89.52 113.16 90 ;
        RECT 28.52 94.96 29 95.44 ;
        RECT 112.68 94.96 113.16 95.44 ;
        RECT 28.52 100.4 29 100.88 ;
        RECT 112.68 100.4 113.16 100.88 ;
      LAYER met4 ;
        RECT 41.1 0 41.7 0.6 ;
        RECT 70.54 0 71.14 0.6 ;
        RECT 99.98 0 100.58 0.6 ;
        RECT 134.94 0 135.54 0.6 ;
        RECT 134.94 75.56 135.54 76.16 ;
        RECT 41.1 102.76 41.7 103.36 ;
        RECT 70.54 102.76 71.14 103.36 ;
        RECT 99.98 102.76 100.58 103.36 ;
      LAYER met5 ;
        RECT 0 16.08 3.2 19.28 ;
        RECT 138.48 16.08 141.68 19.28 ;
        RECT 0 56.88 3.2 60.08 ;
        RECT 138.48 56.88 141.68 60.08 ;
        RECT 28.52 95.64 31.72 98.84 ;
        RECT 109.96 95.64 113.16 98.84 ;
    END
  END VDD
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 0 141.68 0.24 ;
        RECT 0 5.2 0.48 5.68 ;
        RECT 141.2 5.2 141.68 5.68 ;
        RECT 0 10.64 0.48 11.12 ;
        RECT 141.2 10.64 141.68 11.12 ;
        RECT 0 16.08 0.48 16.56 ;
        RECT 141.2 16.08 141.68 16.56 ;
        RECT 0 21.52 0.48 22 ;
        RECT 141.2 21.52 141.68 22 ;
        RECT 0 26.96 0.48 27.44 ;
        RECT 141.2 26.96 141.68 27.44 ;
        RECT 0 32.4 0.48 32.88 ;
        RECT 141.2 32.4 141.68 32.88 ;
        RECT 0 37.84 0.48 38.32 ;
        RECT 141.2 37.84 141.68 38.32 ;
        RECT 0 43.28 0.48 43.76 ;
        RECT 141.2 43.28 141.68 43.76 ;
        RECT 0 48.72 0.48 49.2 ;
        RECT 141.2 48.72 141.68 49.2 ;
        RECT 0 54.16 0.48 54.64 ;
        RECT 141.2 54.16 141.68 54.64 ;
        RECT 0 59.6 0.48 60.08 ;
        RECT 141.2 59.6 141.68 60.08 ;
        RECT 0 65.04 0.48 65.52 ;
        RECT 141.2 65.04 141.68 65.52 ;
        RECT 0 70.48 0.48 70.96 ;
        RECT 141.2 70.48 141.68 70.96 ;
        RECT 0 75.92 141.68 76.4 ;
        RECT 28.52 81.36 29 81.84 ;
        RECT 112.68 81.36 113.16 81.84 ;
        RECT 28.52 86.8 29 87.28 ;
        RECT 112.68 86.8 113.16 87.28 ;
        RECT 28.52 92.24 29 92.72 ;
        RECT 112.68 92.24 113.16 92.72 ;
        RECT 28.52 97.68 29 98.16 ;
        RECT 112.68 97.68 113.16 98.16 ;
        RECT 28.52 103.12 113.16 103.36 ;
      LAYER met4 ;
        RECT 6.14 0 6.74 0.6 ;
        RECT 55.82 0 56.42 0.6 ;
        RECT 85.26 0 85.86 0.6 ;
        RECT 6.14 75.56 6.74 76.16 ;
        RECT 55.82 102.76 56.42 103.36 ;
        RECT 85.26 102.76 85.86 103.36 ;
      LAYER met5 ;
        RECT 0 36.48 3.2 39.68 ;
        RECT 138.48 36.48 141.68 39.68 ;
    END
  END VSS
  OBS
    LAYER li1 ;
      RECT 28.52 103.275 113.16 103.445 ;
      RECT 109.48 100.555 113.16 100.725 ;
      RECT 28.52 100.555 32.2 100.725 ;
      RECT 109.48 97.835 113.16 98.005 ;
      RECT 28.52 97.835 32.2 98.005 ;
      RECT 109.48 95.115 113.16 95.285 ;
      RECT 28.52 95.115 32.2 95.285 ;
      RECT 112.24 92.395 113.16 92.565 ;
      RECT 28.52 92.395 32.2 92.565 ;
      RECT 112.7 89.675 113.16 89.845 ;
      RECT 28.52 89.675 32.2 89.845 ;
      RECT 112.24 86.955 113.16 87.125 ;
      RECT 28.52 86.955 32.2 87.125 ;
      RECT 112.24 84.235 113.16 84.405 ;
      RECT 28.52 84.235 32.2 84.405 ;
      RECT 112.24 81.515 113.16 81.685 ;
      RECT 28.52 81.515 32.2 81.685 ;
      RECT 112.24 78.795 113.16 78.965 ;
      RECT 28.52 78.795 32.2 78.965 ;
      RECT 112.24 76.075 141.68 76.245 ;
      RECT 0 76.075 30.36 76.245 ;
      RECT 138 73.355 141.68 73.525 ;
      RECT 0 73.355 3.68 73.525 ;
      RECT 140.76 70.635 141.68 70.805 ;
      RECT 0 70.635 1.84 70.805 ;
      RECT 140.76 67.915 141.68 68.085 ;
      RECT 0 67.915 1.84 68.085 ;
      RECT 140.76 65.195 141.68 65.365 ;
      RECT 0 65.195 1.84 65.365 ;
      RECT 140.76 62.475 141.68 62.645 ;
      RECT 0 62.475 1.84 62.645 ;
      RECT 140.76 59.755 141.68 59.925 ;
      RECT 0 59.755 1.84 59.925 ;
      RECT 140.76 57.035 141.68 57.205 ;
      RECT 0 57.035 1.84 57.205 ;
      RECT 140.76 54.315 141.68 54.485 ;
      RECT 0 54.315 3.68 54.485 ;
      RECT 140.76 51.595 141.68 51.765 ;
      RECT 0 51.595 3.68 51.765 ;
      RECT 140.76 48.875 141.68 49.045 ;
      RECT 0 48.875 1.84 49.045 ;
      RECT 140.76 46.155 141.68 46.325 ;
      RECT 0 46.155 1.84 46.325 ;
      RECT 140.76 43.435 141.68 43.605 ;
      RECT 0 43.435 1.84 43.605 ;
      RECT 140.76 40.715 141.68 40.885 ;
      RECT 0 40.715 1.84 40.885 ;
      RECT 140.76 37.995 141.68 38.165 ;
      RECT 0 37.995 1.84 38.165 ;
      RECT 140.76 35.275 141.68 35.445 ;
      RECT 0 35.275 1.84 35.445 ;
      RECT 140.76 32.555 141.68 32.725 ;
      RECT 0 32.555 1.84 32.725 ;
      RECT 140.76 29.835 141.68 30.005 ;
      RECT 0 29.835 1.84 30.005 ;
      RECT 140.76 27.115 141.68 27.285 ;
      RECT 0 27.115 1.84 27.285 ;
      RECT 140.76 24.395 141.68 24.565 ;
      RECT 0 24.395 1.84 24.565 ;
      RECT 140.76 21.675 141.68 21.845 ;
      RECT 0 21.675 1.84 21.845 ;
      RECT 139.84 18.955 141.68 19.125 ;
      RECT 0 18.955 1.84 19.125 ;
      RECT 138 16.235 141.68 16.405 ;
      RECT 0 16.235 3.68 16.405 ;
      RECT 138 13.515 141.68 13.685 ;
      RECT 0 13.515 3.68 13.685 ;
      RECT 139.84 10.795 141.68 10.965 ;
      RECT 0 10.795 1.84 10.965 ;
      RECT 139.84 8.075 141.68 8.245 ;
      RECT 0 8.075 3.68 8.245 ;
      RECT 139.84 5.355 141.68 5.525 ;
      RECT 0 5.355 3.68 5.525 ;
      RECT 139.84 2.635 141.68 2.805 ;
      RECT 0 2.635 3.68 2.805 ;
      RECT 0 -0.085 141.68 0.085 ;
    LAYER met2 ;
      RECT 85.42 103.175 85.7 103.545 ;
      RECT 55.98 103.175 56.26 103.545 ;
      RECT 84.05 101.5 84.31 101.82 ;
      RECT 6.3 75.975 6.58 76.345 ;
      RECT 85.42 -0.185 85.7 0.185 ;
      RECT 55.98 -0.185 56.26 0.185 ;
      RECT 6.3 -0.185 6.58 0.185 ;
      POLYGON 112.88 103.08 112.88 75.88 135.35 75.88 135.35 74.52 136.05 74.52 136.05 75.88 136.27 75.88 136.27 74.52 136.97 74.52 136.97 75.88 137.19 75.88 137.19 74.52 137.89 74.52 137.89 75.88 138.11 75.88 138.11 74.52 138.81 74.52 138.81 75.88 139.03 75.88 139.03 74.52 139.73 74.52 139.73 75.88 141.4 75.88 141.4 0.28 139.73 0.28 139.73 1.64 139.03 1.64 139.03 0.28 138.81 0.28 138.81 1.64 138.11 1.64 138.11 0.28 2.65 0.28 2.65 1.64 1.95 1.64 1.95 0.28 0.28 0.28 0.28 75.88 1.95 75.88 1.95 74.52 2.65 74.52 2.65 75.88 2.87 75.88 2.87 74.52 3.57 74.52 3.57 75.88 3.79 75.88 3.79 74.52 4.49 74.52 4.49 75.88 4.71 75.88 4.71 74.52 5.41 74.52 5.41 75.88 7.01 75.88 7.01 74.52 7.71 74.52 7.71 75.88 10.23 75.88 10.23 74.52 10.93 74.52 10.93 75.88 11.15 75.88 11.15 74.52 11.85 74.52 11.85 75.88 28.8 75.88 28.8 103.08 30.47 103.08 30.47 101.72 31.17 101.72 31.17 103.08 31.85 103.08 31.85 101.72 32.55 101.72 32.55 103.08 32.77 103.08 32.77 101.72 33.47 101.72 33.47 103.08 49.79 103.08 49.79 101.72 50.49 101.72 50.49 103.08 50.71 103.08 50.71 101.72 51.41 101.72 51.41 103.08 51.63 103.08 51.63 101.72 52.33 101.72 52.33 103.08 52.55 103.08 52.55 101.72 53.25 101.72 53.25 103.08 53.47 103.08 53.47 101.72 54.17 101.72 54.17 103.08 54.39 103.08 54.39 101.72 55.09 101.72 55.09 103.08 57.15 103.08 57.15 101.72 57.85 101.72 57.85 103.08 58.07 103.08 58.07 101.72 58.77 101.72 58.77 103.08 58.99 103.08 58.99 101.72 59.69 101.72 59.69 103.08 59.91 103.08 59.91 101.72 60.61 101.72 60.61 103.08 60.83 103.08 60.83 101.72 61.53 101.72 61.53 103.08 61.75 103.08 61.75 101.72 62.45 101.72 62.45 103.08 63.13 103.08 63.13 101.72 63.83 101.72 63.83 103.08 64.05 103.08 64.05 101.72 64.75 101.72 64.75 103.08 66.35 103.08 66.35 101.72 67.05 101.72 67.05 103.08 67.27 103.08 67.27 101.72 67.97 101.72 67.97 103.08 68.19 103.08 68.19 101.72 68.89 101.72 68.89 103.08 69.11 103.08 69.11 101.72 69.81 101.72 69.81 103.08 70.03 103.08 70.03 101.72 70.73 101.72 70.73 103.08 70.95 103.08 70.95 101.72 71.65 101.72 71.65 103.08 71.87 103.08 71.87 101.72 72.57 101.72 72.57 103.08 72.79 103.08 72.79 101.72 73.49 101.72 73.49 103.08 73.71 103.08 73.71 101.72 74.41 101.72 74.41 103.08 74.63 103.08 74.63 101.72 75.33 101.72 75.33 103.08 75.55 103.08 75.55 101.72 76.25 101.72 76.25 103.08 76.47 103.08 76.47 101.72 77.17 101.72 77.17 103.08 77.39 103.08 77.39 101.72 78.09 101.72 78.09 103.08 78.31 103.08 78.31 101.72 79.01 101.72 79.01 103.08 79.23 103.08 79.23 101.72 79.93 101.72 79.93 103.08 80.15 103.08 80.15 101.72 80.85 101.72 80.85 103.08 81.07 103.08 81.07 101.72 81.77 101.72 81.77 103.08 81.99 103.08 81.99 101.72 82.69 101.72 82.69 103.08 83.37 103.08 83.37 101.72 84.07 101.72 84.07 103.08 84.29 103.08 84.29 101.72 84.99 101.72 84.99 103.08 86.59 103.08 86.59 101.72 87.29 101.72 87.29 103.08 93.49 103.08 93.49 101.72 94.19 101.72 94.19 103.08 95.33 103.08 95.33 101.72 96.03 101.72 96.03 103.08 96.25 103.08 96.25 101.72 96.95 101.72 96.95 103.08 97.17 103.08 97.17 101.72 97.87 101.72 97.87 103.08 98.55 103.08 98.55 101.72 99.25 101.72 99.25 103.08 ;
    LAYER met4 ;
      POLYGON 112.76 102.96 112.76 75.76 134.54 75.76 134.54 75.16 135.94 75.16 135.94 75.76 141.28 75.76 141.28 0.4 135.94 0.4 135.94 1 134.54 1 134.54 0.4 100.98 0.4 100.98 1 99.58 1 99.58 0.4 86.26 0.4 86.26 1 84.86 1 84.86 0.4 71.54 0.4 71.54 1 70.14 1 70.14 0.4 56.82 0.4 56.82 1 55.42 1 55.42 0.4 42.1 0.4 42.1 1 40.7 1 40.7 0.4 7.14 0.4 7.14 1 5.74 1 5.74 0.4 0.4 0.4 0.4 75.76 5.74 75.76 5.74 75.16 7.14 75.16 7.14 75.76 28.92 75.76 28.92 102.96 32.57 102.96 32.57 101.6 33.67 101.6 33.67 102.96 40.7 102.96 40.7 102.36 42.1 102.36 42.1 102.96 55.42 102.96 55.42 102.36 56.82 102.36 56.82 102.96 70.14 102.96 70.14 102.36 71.54 102.36 71.54 102.96 84.86 102.96 84.86 102.36 86.26 102.36 86.26 102.96 99.58 102.96 99.58 102.36 100.98 102.36 100.98 102.96 ;
    LAYER met3 ;
      POLYGON 85.725 103.525 85.725 103.52 85.94 103.52 85.94 103.2 85.725 103.2 85.725 103.195 85.395 103.195 85.395 103.2 85.18 103.2 85.18 103.52 85.395 103.52 85.395 103.525 ;
      POLYGON 56.285 103.525 56.285 103.52 56.5 103.52 56.5 103.2 56.285 103.2 56.285 103.195 55.955 103.195 55.955 103.2 55.74 103.2 55.74 103.52 55.955 103.52 55.955 103.525 ;
      POLYGON 6.605 76.325 6.605 76.32 6.82 76.32 6.82 76 6.605 76 6.605 75.995 6.275 75.995 6.275 76 6.06 76 6.06 76.32 6.275 76.32 6.275 76.325 ;
      POLYGON 38.79 71.55 38.79 71.25 1.78 71.25 1.78 71.27 1.23 71.27 1.23 71.55 ;
      POLYGON 140.45 57.95 140.45 57.67 139.9 57.67 139.9 57.65 136.93 57.65 136.93 57.95 ;
      POLYGON 24.53 55.23 24.53 54.93 1.78 54.93 1.78 54.95 1.23 54.95 1.23 55.23 ;
      POLYGON 2.03 40.28 2.03 40.27 7.05 40.27 7.05 39.97 2.03 39.97 2.03 39.96 1.65 39.96 1.65 40.28 ;
      POLYGON 6.13 28.03 6.13 27.73 1.78 27.73 1.78 27.75 1.23 27.75 1.23 28.03 ;
      POLYGON 140.03 22.6 140.03 22.28 139.65 22.28 139.65 22.29 58.73 22.29 58.73 22.59 139.65 22.59 139.65 22.6 ;
      POLYGON 85.725 0.165 85.725 0.16 85.94 0.16 85.94 -0.16 85.725 -0.16 85.725 -0.165 85.395 -0.165 85.395 -0.16 85.18 -0.16 85.18 0.16 85.395 0.16 85.395 0.165 ;
      POLYGON 56.285 0.165 56.285 0.16 56.5 0.16 56.5 -0.16 56.285 -0.16 56.285 -0.165 55.955 -0.165 55.955 -0.16 55.74 -0.16 55.74 0.16 55.955 0.16 55.955 0.165 ;
      POLYGON 6.605 0.165 6.605 0.16 6.82 0.16 6.82 -0.16 6.605 -0.16 6.605 -0.165 6.275 -0.165 6.275 -0.16 6.06 -0.16 6.06 0.16 6.275 0.16 6.275 0.165 ;
      POLYGON 112.76 102.96 112.76 99.83 111.38 99.83 111.38 98.73 112.76 98.73 112.76 92.35 111.38 92.35 111.38 91.25 112.76 91.25 112.76 90.99 111.38 90.99 111.38 89.89 112.76 89.89 112.76 75.76 141.28 75.76 141.28 72.63 139.9 72.63 139.9 71.53 141.28 71.53 141.28 69.91 139.9 69.91 139.9 68.81 141.28 68.81 141.28 68.55 139.9 68.55 139.9 67.45 141.28 67.45 141.28 67.19 139.9 67.19 139.9 66.09 141.28 66.09 141.28 64.47 139.9 64.47 139.9 63.37 141.28 63.37 141.28 63.11 139.9 63.11 139.9 62.01 141.28 62.01 141.28 61.75 139.9 61.75 139.9 60.65 141.28 60.65 141.28 60.39 139.9 60.39 139.9 59.29 141.28 59.29 141.28 59.03 139.9 59.03 139.9 57.93 141.28 57.93 141.28 57.67 139.9 57.67 139.9 56.57 141.28 56.57 141.28 56.31 139.9 56.31 139.9 55.21 141.28 55.21 141.28 53.59 139.9 53.59 139.9 52.49 141.28 52.49 141.28 52.23 139.9 52.23 139.9 51.13 141.28 51.13 141.28 50.87 139.9 50.87 139.9 49.77 141.28 49.77 141.28 48.15 139.9 48.15 139.9 47.05 141.28 47.05 141.28 46.79 139.9 46.79 139.9 45.69 141.28 45.69 141.28 45.43 139.9 45.43 139.9 44.33 141.28 44.33 141.28 42.71 139.9 42.71 139.9 41.61 141.28 41.61 141.28 41.35 139.9 41.35 139.9 40.25 141.28 40.25 141.28 39.99 139.9 39.99 139.9 38.89 141.28 38.89 141.28 37.27 139.9 37.27 139.9 36.17 141.28 36.17 141.28 35.91 139.9 35.91 139.9 34.81 141.28 34.81 141.28 34.55 139.9 34.55 139.9 33.45 141.28 33.45 141.28 31.83 139.9 31.83 139.9 30.73 141.28 30.73 141.28 30.47 139.9 30.47 139.9 29.37 141.28 29.37 141.28 29.11 139.9 29.11 139.9 28.01 141.28 28.01 141.28 26.39 139.9 26.39 139.9 25.29 141.28 25.29 141.28 25.03 139.9 25.03 139.9 23.93 141.28 23.93 141.28 23.67 139.9 23.67 139.9 22.57 141.28 22.57 141.28 20.95 139.9 20.95 139.9 19.85 141.28 19.85 141.28 19.59 139.9 19.59 139.9 18.49 141.28 18.49 141.28 18.23 139.9 18.23 139.9 17.13 141.28 17.13 141.28 16.87 139.9 16.87 139.9 15.77 141.28 15.77 141.28 15.51 139.9 15.51 139.9 14.41 141.28 14.41 141.28 14.15 139.9 14.15 139.9 13.05 141.28 13.05 141.28 12.79 139.9 12.79 139.9 11.69 141.28 11.69 141.28 10.07 139.9 10.07 139.9 8.97 141.28 8.97 141.28 8.71 139.9 8.71 139.9 7.61 141.28 7.61 141.28 7.35 139.9 7.35 139.9 6.25 141.28 6.25 141.28 4.63 139.9 4.63 139.9 3.53 141.28 3.53 141.28 0.4 0.4 0.4 0.4 3.53 1.78 3.53 1.78 4.63 0.4 4.63 0.4 4.89 1.78 4.89 1.78 5.99 0.4 5.99 0.4 6.25 1.78 6.25 1.78 7.35 0.4 7.35 0.4 9.65 1.78 9.65 1.78 10.75 0.4 10.75 0.4 11.01 1.78 11.01 1.78 12.11 0.4 12.11 0.4 15.09 1.78 15.09 1.78 16.19 0.4 16.19 0.4 17.13 1.78 17.13 1.78 18.23 0.4 18.23 0.4 18.49 1.78 18.49 1.78 19.59 0.4 19.59 0.4 19.85 1.78 19.85 1.78 20.95 0.4 20.95 0.4 21.21 1.78 21.21 1.78 22.31 0.4 22.31 0.4 22.57 1.78 22.57 1.78 23.67 0.4 23.67 0.4 25.29 1.78 25.29 1.78 26.39 0.4 26.39 0.4 26.65 1.78 26.65 1.78 27.75 0.4 27.75 0.4 28.01 1.78 28.01 1.78 29.11 0.4 29.11 0.4 30.73 1.78 30.73 1.78 31.83 0.4 31.83 0.4 32.09 1.78 32.09 1.78 33.19 0.4 33.19 0.4 33.45 1.78 33.45 1.78 34.55 0.4 34.55 0.4 36.17 1.78 36.17 1.78 37.27 0.4 37.27 0.4 37.53 1.78 37.53 1.78 38.63 0.4 38.63 0.4 38.89 1.78 38.89 1.78 39.99 0.4 39.99 0.4 41.61 1.78 41.61 1.78 42.71 0.4 42.71 0.4 42.97 1.78 42.97 1.78 44.07 0.4 44.07 0.4 44.33 1.78 44.33 1.78 45.43 0.4 45.43 0.4 47.05 1.78 47.05 1.78 48.15 0.4 48.15 0.4 48.41 1.78 48.41 1.78 49.51 0.4 49.51 0.4 49.77 1.78 49.77 1.78 50.87 0.4 50.87 0.4 51.13 1.78 51.13 1.78 52.23 0.4 52.23 0.4 52.49 1.78 52.49 1.78 53.59 0.4 53.59 0.4 53.85 1.78 53.85 1.78 54.95 0.4 54.95 0.4 55.21 1.78 55.21 1.78 56.31 0.4 56.31 0.4 56.57 1.78 56.57 1.78 57.67 0.4 57.67 0.4 57.93 1.78 57.93 1.78 59.03 0.4 59.03 0.4 59.29 1.78 59.29 1.78 60.39 0.4 60.39 0.4 60.65 1.78 60.65 1.78 61.75 0.4 61.75 0.4 62.01 1.78 62.01 1.78 63.11 0.4 63.11 0.4 64.05 1.78 64.05 1.78 65.15 0.4 65.15 0.4 65.41 1.78 65.41 1.78 66.51 0.4 66.51 0.4 66.77 1.78 66.77 1.78 67.87 0.4 67.87 0.4 68.81 1.78 68.81 1.78 69.91 0.4 69.91 0.4 70.17 1.78 70.17 1.78 71.27 0.4 71.27 0.4 71.53 1.78 71.53 1.78 72.63 0.4 72.63 0.4 75.76 28.92 75.76 28.92 89.89 30.3 89.89 30.3 90.99 28.92 90.99 28.92 91.25 30.3 91.25 30.3 92.35 28.92 92.35 28.92 94.65 30.3 94.65 30.3 95.75 28.92 95.75 28.92 96.01 30.3 96.01 30.3 97.11 28.92 97.11 28.92 97.37 30.3 97.37 30.3 98.47 28.92 98.47 28.92 99.41 30.3 99.41 30.3 100.51 28.92 100.51 28.92 102.96 ;
    LAYER met5 ;
      POLYGON 106.76 100.16 106.76 92.44 109.96 92.44 109.96 72.96 138.48 72.96 138.48 63.28 135.28 63.28 135.28 53.68 138.48 53.68 138.48 42.88 135.28 42.88 135.28 33.28 138.48 33.28 138.48 22.48 135.28 22.48 135.28 12.88 138.48 12.88 138.48 3.2 3.2 3.2 3.2 12.88 6.4 12.88 6.4 22.48 3.2 22.48 3.2 33.28 6.4 33.28 6.4 42.88 3.2 42.88 3.2 53.68 6.4 53.68 6.4 63.28 3.2 63.28 3.2 72.96 31.72 72.96 31.72 92.44 34.92 92.44 34.92 100.16 ;
    LAYER met1 ;
      POLYGON 112.88 102.84 112.88 101.16 112.4 101.16 112.4 100.12 112.88 100.12 112.88 98.44 112.4 98.44 112.4 97.4 112.88 97.4 112.88 95.72 112.4 95.72 112.4 94.68 112.88 94.68 112.88 93 112.4 93 112.4 91.96 112.88 91.96 112.88 90.28 112.4 90.28 112.4 89.24 112.88 89.24 112.88 87.56 112.4 87.56 112.4 86.52 112.88 86.52 112.88 84.84 112.4 84.84 112.4 83.8 112.88 83.8 112.88 82.12 112.4 82.12 112.4 81.08 112.88 81.08 112.88 79.4 112.4 79.4 112.4 78.36 112.88 78.36 112.88 76.68 28.8 76.68 28.8 78.36 29.28 78.36 29.28 79.4 28.8 79.4 28.8 81.08 29.28 81.08 29.28 82.12 28.8 82.12 28.8 83.8 29.28 83.8 29.28 84.84 28.8 84.84 28.8 86.52 29.28 86.52 29.28 87.56 28.8 87.56 28.8 89.24 29.28 89.24 29.28 90.28 28.8 90.28 28.8 91.96 29.28 91.96 29.28 93 28.8 93 28.8 94.68 29.28 94.68 29.28 95.72 28.8 95.72 28.8 97.4 29.28 97.4 29.28 98.44 28.8 98.44 28.8 100.12 29.28 100.12 29.28 101.16 28.8 101.16 28.8 102.84 ;
      POLYGON 141.4 75.64 141.4 73.96 140.92 73.96 140.92 72.92 141.4 72.92 141.4 71.24 140.92 71.24 140.92 70.2 141.4 70.2 141.4 68.52 140.92 68.52 140.92 67.48 141.4 67.48 141.4 65.8 140.92 65.8 140.92 64.76 141.4 64.76 141.4 63.08 140.92 63.08 140.92 62.04 141.4 62.04 141.4 60.36 140.92 60.36 140.92 59.32 141.4 59.32 141.4 57.64 140.92 57.64 140.92 56.6 141.4 56.6 141.4 54.92 140.92 54.92 140.92 53.88 141.4 53.88 141.4 52.2 140.92 52.2 140.92 51.16 141.4 51.16 141.4 49.48 140.92 49.48 140.92 48.44 141.4 48.44 141.4 46.76 140.92 46.76 140.92 45.72 141.4 45.72 141.4 44.04 140.92 44.04 140.92 43 141.4 43 141.4 41.32 140.92 41.32 140.92 40.28 141.4 40.28 141.4 38.6 140.92 38.6 140.92 37.56 141.4 37.56 141.4 35.88 140.92 35.88 140.92 34.84 141.4 34.84 141.4 33.16 140.92 33.16 140.92 32.12 141.4 32.12 141.4 30.44 140.92 30.44 140.92 29.4 141.4 29.4 141.4 27.72 140.92 27.72 140.92 26.68 141.4 26.68 141.4 25 140.92 25 140.92 23.96 141.4 23.96 141.4 22.28 140.92 22.28 140.92 21.24 141.4 21.24 141.4 19.56 140.92 19.56 140.92 18.52 141.4 18.52 141.4 16.84 140.92 16.84 140.92 15.8 141.4 15.8 141.4 14.12 140.92 14.12 140.92 13.08 141.4 13.08 141.4 11.4 140.92 11.4 140.92 10.36 141.4 10.36 141.4 8.68 140.92 8.68 140.92 7.64 141.4 7.64 141.4 5.96 140.92 5.96 140.92 4.92 141.4 4.92 141.4 3.24 140.92 3.24 140.92 2.2 141.4 2.2 141.4 0.52 0.28 0.52 0.28 2.2 0.76 2.2 0.76 3.24 0.28 3.24 0.28 4.92 0.76 4.92 0.76 5.96 0.28 5.96 0.28 7.64 0.76 7.64 0.76 8.68 0.28 8.68 0.28 10.36 0.76 10.36 0.76 11.4 0.28 11.4 0.28 13.08 0.76 13.08 0.76 14.12 0.28 14.12 0.28 15.8 0.76 15.8 0.76 16.84 0.28 16.84 0.28 18.52 0.76 18.52 0.76 19.56 0.28 19.56 0.28 21.24 0.76 21.24 0.76 22.28 0.28 22.28 0.28 23.96 0.76 23.96 0.76 25 0.28 25 0.28 26.68 0.76 26.68 0.76 27.72 0.28 27.72 0.28 29.4 0.76 29.4 0.76 30.44 0.28 30.44 0.28 32.12 0.76 32.12 0.76 33.16 0.28 33.16 0.28 34.84 0.76 34.84 0.76 35.88 0.28 35.88 0.28 37.56 0.76 37.56 0.76 38.6 0.28 38.6 0.28 40.28 0.76 40.28 0.76 41.32 0.28 41.32 0.28 43 0.76 43 0.76 44.04 0.28 44.04 0.28 45.72 0.76 45.72 0.76 46.76 0.28 46.76 0.28 48.44 0.76 48.44 0.76 49.48 0.28 49.48 0.28 51.16 0.76 51.16 0.76 52.2 0.28 52.2 0.28 53.88 0.76 53.88 0.76 54.92 0.28 54.92 0.28 56.6 0.76 56.6 0.76 57.64 0.28 57.64 0.28 59.32 0.76 59.32 0.76 60.36 0.28 60.36 0.28 62.04 0.76 62.04 0.76 63.08 0.28 63.08 0.28 64.76 0.76 64.76 0.76 65.8 0.28 65.8 0.28 67.48 0.76 67.48 0.76 68.52 0.28 68.52 0.28 70.2 0.76 70.2 0.76 71.24 0.28 71.24 0.28 72.92 0.76 72.92 0.76 73.96 0.28 73.96 0.28 75.64 ;
    LAYER li1 ;
      POLYGON 112.82 103.02 112.82 75.82 141.34 75.82 141.34 0.34 0.34 0.34 0.34 75.82 28.86 75.82 28.86 103.02 ;
    LAYER mcon ;
      RECT 112.845 103.275 113.015 103.445 ;
      RECT 112.385 103.275 112.555 103.445 ;
      RECT 111.925 103.275 112.095 103.445 ;
      RECT 111.465 103.275 111.635 103.445 ;
      RECT 111.005 103.275 111.175 103.445 ;
      RECT 110.545 103.275 110.715 103.445 ;
      RECT 110.085 103.275 110.255 103.445 ;
      RECT 109.625 103.275 109.795 103.445 ;
      RECT 109.165 103.275 109.335 103.445 ;
      RECT 108.705 103.275 108.875 103.445 ;
      RECT 108.245 103.275 108.415 103.445 ;
      RECT 107.785 103.275 107.955 103.445 ;
      RECT 107.325 103.275 107.495 103.445 ;
      RECT 106.865 103.275 107.035 103.445 ;
      RECT 106.405 103.275 106.575 103.445 ;
      RECT 105.945 103.275 106.115 103.445 ;
      RECT 105.485 103.275 105.655 103.445 ;
      RECT 105.025 103.275 105.195 103.445 ;
      RECT 104.565 103.275 104.735 103.445 ;
      RECT 104.105 103.275 104.275 103.445 ;
      RECT 103.645 103.275 103.815 103.445 ;
      RECT 103.185 103.275 103.355 103.445 ;
      RECT 102.725 103.275 102.895 103.445 ;
      RECT 102.265 103.275 102.435 103.445 ;
      RECT 101.805 103.275 101.975 103.445 ;
      RECT 101.345 103.275 101.515 103.445 ;
      RECT 100.885 103.275 101.055 103.445 ;
      RECT 100.425 103.275 100.595 103.445 ;
      RECT 99.965 103.275 100.135 103.445 ;
      RECT 99.505 103.275 99.675 103.445 ;
      RECT 99.045 103.275 99.215 103.445 ;
      RECT 98.585 103.275 98.755 103.445 ;
      RECT 98.125 103.275 98.295 103.445 ;
      RECT 97.665 103.275 97.835 103.445 ;
      RECT 97.205 103.275 97.375 103.445 ;
      RECT 96.745 103.275 96.915 103.445 ;
      RECT 96.285 103.275 96.455 103.445 ;
      RECT 95.825 103.275 95.995 103.445 ;
      RECT 95.365 103.275 95.535 103.445 ;
      RECT 94.905 103.275 95.075 103.445 ;
      RECT 94.445 103.275 94.615 103.445 ;
      RECT 93.985 103.275 94.155 103.445 ;
      RECT 93.525 103.275 93.695 103.445 ;
      RECT 93.065 103.275 93.235 103.445 ;
      RECT 92.605 103.275 92.775 103.445 ;
      RECT 92.145 103.275 92.315 103.445 ;
      RECT 91.685 103.275 91.855 103.445 ;
      RECT 91.225 103.275 91.395 103.445 ;
      RECT 90.765 103.275 90.935 103.445 ;
      RECT 90.305 103.275 90.475 103.445 ;
      RECT 89.845 103.275 90.015 103.445 ;
      RECT 89.385 103.275 89.555 103.445 ;
      RECT 88.925 103.275 89.095 103.445 ;
      RECT 88.465 103.275 88.635 103.445 ;
      RECT 88.005 103.275 88.175 103.445 ;
      RECT 87.545 103.275 87.715 103.445 ;
      RECT 87.085 103.275 87.255 103.445 ;
      RECT 86.625 103.275 86.795 103.445 ;
      RECT 86.165 103.275 86.335 103.445 ;
      RECT 85.705 103.275 85.875 103.445 ;
      RECT 85.245 103.275 85.415 103.445 ;
      RECT 84.785 103.275 84.955 103.445 ;
      RECT 84.325 103.275 84.495 103.445 ;
      RECT 83.865 103.275 84.035 103.445 ;
      RECT 83.405 103.275 83.575 103.445 ;
      RECT 82.945 103.275 83.115 103.445 ;
      RECT 82.485 103.275 82.655 103.445 ;
      RECT 82.025 103.275 82.195 103.445 ;
      RECT 81.565 103.275 81.735 103.445 ;
      RECT 81.105 103.275 81.275 103.445 ;
      RECT 80.645 103.275 80.815 103.445 ;
      RECT 80.185 103.275 80.355 103.445 ;
      RECT 79.725 103.275 79.895 103.445 ;
      RECT 79.265 103.275 79.435 103.445 ;
      RECT 78.805 103.275 78.975 103.445 ;
      RECT 78.345 103.275 78.515 103.445 ;
      RECT 77.885 103.275 78.055 103.445 ;
      RECT 77.425 103.275 77.595 103.445 ;
      RECT 76.965 103.275 77.135 103.445 ;
      RECT 76.505 103.275 76.675 103.445 ;
      RECT 76.045 103.275 76.215 103.445 ;
      RECT 75.585 103.275 75.755 103.445 ;
      RECT 75.125 103.275 75.295 103.445 ;
      RECT 74.665 103.275 74.835 103.445 ;
      RECT 74.205 103.275 74.375 103.445 ;
      RECT 73.745 103.275 73.915 103.445 ;
      RECT 73.285 103.275 73.455 103.445 ;
      RECT 72.825 103.275 72.995 103.445 ;
      RECT 72.365 103.275 72.535 103.445 ;
      RECT 71.905 103.275 72.075 103.445 ;
      RECT 71.445 103.275 71.615 103.445 ;
      RECT 70.985 103.275 71.155 103.445 ;
      RECT 70.525 103.275 70.695 103.445 ;
      RECT 70.065 103.275 70.235 103.445 ;
      RECT 69.605 103.275 69.775 103.445 ;
      RECT 69.145 103.275 69.315 103.445 ;
      RECT 68.685 103.275 68.855 103.445 ;
      RECT 68.225 103.275 68.395 103.445 ;
      RECT 67.765 103.275 67.935 103.445 ;
      RECT 67.305 103.275 67.475 103.445 ;
      RECT 66.845 103.275 67.015 103.445 ;
      RECT 66.385 103.275 66.555 103.445 ;
      RECT 65.925 103.275 66.095 103.445 ;
      RECT 65.465 103.275 65.635 103.445 ;
      RECT 65.005 103.275 65.175 103.445 ;
      RECT 64.545 103.275 64.715 103.445 ;
      RECT 64.085 103.275 64.255 103.445 ;
      RECT 63.625 103.275 63.795 103.445 ;
      RECT 63.165 103.275 63.335 103.445 ;
      RECT 62.705 103.275 62.875 103.445 ;
      RECT 62.245 103.275 62.415 103.445 ;
      RECT 61.785 103.275 61.955 103.445 ;
      RECT 61.325 103.275 61.495 103.445 ;
      RECT 60.865 103.275 61.035 103.445 ;
      RECT 60.405 103.275 60.575 103.445 ;
      RECT 59.945 103.275 60.115 103.445 ;
      RECT 59.485 103.275 59.655 103.445 ;
      RECT 59.025 103.275 59.195 103.445 ;
      RECT 58.565 103.275 58.735 103.445 ;
      RECT 58.105 103.275 58.275 103.445 ;
      RECT 57.645 103.275 57.815 103.445 ;
      RECT 57.185 103.275 57.355 103.445 ;
      RECT 56.725 103.275 56.895 103.445 ;
      RECT 56.265 103.275 56.435 103.445 ;
      RECT 55.805 103.275 55.975 103.445 ;
      RECT 55.345 103.275 55.515 103.445 ;
      RECT 54.885 103.275 55.055 103.445 ;
      RECT 54.425 103.275 54.595 103.445 ;
      RECT 53.965 103.275 54.135 103.445 ;
      RECT 53.505 103.275 53.675 103.445 ;
      RECT 53.045 103.275 53.215 103.445 ;
      RECT 52.585 103.275 52.755 103.445 ;
      RECT 52.125 103.275 52.295 103.445 ;
      RECT 51.665 103.275 51.835 103.445 ;
      RECT 51.205 103.275 51.375 103.445 ;
      RECT 50.745 103.275 50.915 103.445 ;
      RECT 50.285 103.275 50.455 103.445 ;
      RECT 49.825 103.275 49.995 103.445 ;
      RECT 49.365 103.275 49.535 103.445 ;
      RECT 48.905 103.275 49.075 103.445 ;
      RECT 48.445 103.275 48.615 103.445 ;
      RECT 47.985 103.275 48.155 103.445 ;
      RECT 47.525 103.275 47.695 103.445 ;
      RECT 47.065 103.275 47.235 103.445 ;
      RECT 46.605 103.275 46.775 103.445 ;
      RECT 46.145 103.275 46.315 103.445 ;
      RECT 45.685 103.275 45.855 103.445 ;
      RECT 45.225 103.275 45.395 103.445 ;
      RECT 44.765 103.275 44.935 103.445 ;
      RECT 44.305 103.275 44.475 103.445 ;
      RECT 43.845 103.275 44.015 103.445 ;
      RECT 43.385 103.275 43.555 103.445 ;
      RECT 42.925 103.275 43.095 103.445 ;
      RECT 42.465 103.275 42.635 103.445 ;
      RECT 42.005 103.275 42.175 103.445 ;
      RECT 41.545 103.275 41.715 103.445 ;
      RECT 41.085 103.275 41.255 103.445 ;
      RECT 40.625 103.275 40.795 103.445 ;
      RECT 40.165 103.275 40.335 103.445 ;
      RECT 39.705 103.275 39.875 103.445 ;
      RECT 39.245 103.275 39.415 103.445 ;
      RECT 38.785 103.275 38.955 103.445 ;
      RECT 38.325 103.275 38.495 103.445 ;
      RECT 37.865 103.275 38.035 103.445 ;
      RECT 37.405 103.275 37.575 103.445 ;
      RECT 36.945 103.275 37.115 103.445 ;
      RECT 36.485 103.275 36.655 103.445 ;
      RECT 36.025 103.275 36.195 103.445 ;
      RECT 35.565 103.275 35.735 103.445 ;
      RECT 35.105 103.275 35.275 103.445 ;
      RECT 34.645 103.275 34.815 103.445 ;
      RECT 34.185 103.275 34.355 103.445 ;
      RECT 33.725 103.275 33.895 103.445 ;
      RECT 33.265 103.275 33.435 103.445 ;
      RECT 32.805 103.275 32.975 103.445 ;
      RECT 32.345 103.275 32.515 103.445 ;
      RECT 31.885 103.275 32.055 103.445 ;
      RECT 31.425 103.275 31.595 103.445 ;
      RECT 30.965 103.275 31.135 103.445 ;
      RECT 30.505 103.275 30.675 103.445 ;
      RECT 30.045 103.275 30.215 103.445 ;
      RECT 29.585 103.275 29.755 103.445 ;
      RECT 29.125 103.275 29.295 103.445 ;
      RECT 28.665 103.275 28.835 103.445 ;
      RECT 112.845 100.555 113.015 100.725 ;
      RECT 112.385 100.555 112.555 100.725 ;
      RECT 29.125 100.555 29.295 100.725 ;
      RECT 28.665 100.555 28.835 100.725 ;
      RECT 112.845 97.835 113.015 98.005 ;
      RECT 112.385 97.835 112.555 98.005 ;
      RECT 29.125 97.835 29.295 98.005 ;
      RECT 28.665 97.835 28.835 98.005 ;
      RECT 112.845 95.115 113.015 95.285 ;
      RECT 112.385 95.115 112.555 95.285 ;
      RECT 29.125 95.115 29.295 95.285 ;
      RECT 28.665 95.115 28.835 95.285 ;
      RECT 112.845 92.395 113.015 92.565 ;
      RECT 112.385 92.395 112.555 92.565 ;
      RECT 29.125 92.395 29.295 92.565 ;
      RECT 28.665 92.395 28.835 92.565 ;
      RECT 112.845 89.675 113.015 89.845 ;
      RECT 112.385 89.675 112.555 89.845 ;
      RECT 29.125 89.675 29.295 89.845 ;
      RECT 28.665 89.675 28.835 89.845 ;
      RECT 112.845 86.955 113.015 87.125 ;
      RECT 112.385 86.955 112.555 87.125 ;
      RECT 29.125 86.955 29.295 87.125 ;
      RECT 28.665 86.955 28.835 87.125 ;
      RECT 112.845 84.235 113.015 84.405 ;
      RECT 112.385 84.235 112.555 84.405 ;
      RECT 29.125 84.235 29.295 84.405 ;
      RECT 28.665 84.235 28.835 84.405 ;
      RECT 112.845 81.515 113.015 81.685 ;
      RECT 112.385 81.515 112.555 81.685 ;
      RECT 29.125 81.515 29.295 81.685 ;
      RECT 28.665 81.515 28.835 81.685 ;
      RECT 112.845 78.795 113.015 78.965 ;
      RECT 112.385 78.795 112.555 78.965 ;
      RECT 29.125 78.795 29.295 78.965 ;
      RECT 28.665 78.795 28.835 78.965 ;
      RECT 141.365 76.075 141.535 76.245 ;
      RECT 140.905 76.075 141.075 76.245 ;
      RECT 140.445 76.075 140.615 76.245 ;
      RECT 139.985 76.075 140.155 76.245 ;
      RECT 139.525 76.075 139.695 76.245 ;
      RECT 139.065 76.075 139.235 76.245 ;
      RECT 138.605 76.075 138.775 76.245 ;
      RECT 138.145 76.075 138.315 76.245 ;
      RECT 137.685 76.075 137.855 76.245 ;
      RECT 137.225 76.075 137.395 76.245 ;
      RECT 136.765 76.075 136.935 76.245 ;
      RECT 136.305 76.075 136.475 76.245 ;
      RECT 135.845 76.075 136.015 76.245 ;
      RECT 135.385 76.075 135.555 76.245 ;
      RECT 134.925 76.075 135.095 76.245 ;
      RECT 134.465 76.075 134.635 76.245 ;
      RECT 134.005 76.075 134.175 76.245 ;
      RECT 133.545 76.075 133.715 76.245 ;
      RECT 133.085 76.075 133.255 76.245 ;
      RECT 132.625 76.075 132.795 76.245 ;
      RECT 132.165 76.075 132.335 76.245 ;
      RECT 131.705 76.075 131.875 76.245 ;
      RECT 131.245 76.075 131.415 76.245 ;
      RECT 130.785 76.075 130.955 76.245 ;
      RECT 130.325 76.075 130.495 76.245 ;
      RECT 129.865 76.075 130.035 76.245 ;
      RECT 129.405 76.075 129.575 76.245 ;
      RECT 128.945 76.075 129.115 76.245 ;
      RECT 128.485 76.075 128.655 76.245 ;
      RECT 128.025 76.075 128.195 76.245 ;
      RECT 127.565 76.075 127.735 76.245 ;
      RECT 127.105 76.075 127.275 76.245 ;
      RECT 126.645 76.075 126.815 76.245 ;
      RECT 126.185 76.075 126.355 76.245 ;
      RECT 125.725 76.075 125.895 76.245 ;
      RECT 125.265 76.075 125.435 76.245 ;
      RECT 124.805 76.075 124.975 76.245 ;
      RECT 124.345 76.075 124.515 76.245 ;
      RECT 123.885 76.075 124.055 76.245 ;
      RECT 123.425 76.075 123.595 76.245 ;
      RECT 122.965 76.075 123.135 76.245 ;
      RECT 122.505 76.075 122.675 76.245 ;
      RECT 122.045 76.075 122.215 76.245 ;
      RECT 121.585 76.075 121.755 76.245 ;
      RECT 121.125 76.075 121.295 76.245 ;
      RECT 120.665 76.075 120.835 76.245 ;
      RECT 120.205 76.075 120.375 76.245 ;
      RECT 119.745 76.075 119.915 76.245 ;
      RECT 119.285 76.075 119.455 76.245 ;
      RECT 118.825 76.075 118.995 76.245 ;
      RECT 118.365 76.075 118.535 76.245 ;
      RECT 117.905 76.075 118.075 76.245 ;
      RECT 117.445 76.075 117.615 76.245 ;
      RECT 116.985 76.075 117.155 76.245 ;
      RECT 116.525 76.075 116.695 76.245 ;
      RECT 116.065 76.075 116.235 76.245 ;
      RECT 115.605 76.075 115.775 76.245 ;
      RECT 115.145 76.075 115.315 76.245 ;
      RECT 114.685 76.075 114.855 76.245 ;
      RECT 114.225 76.075 114.395 76.245 ;
      RECT 113.765 76.075 113.935 76.245 ;
      RECT 113.305 76.075 113.475 76.245 ;
      RECT 112.845 76.075 113.015 76.245 ;
      RECT 112.385 76.075 112.555 76.245 ;
      RECT 111.925 76.075 112.095 76.245 ;
      RECT 111.465 76.075 111.635 76.245 ;
      RECT 111.005 76.075 111.175 76.245 ;
      RECT 110.545 76.075 110.715 76.245 ;
      RECT 110.085 76.075 110.255 76.245 ;
      RECT 109.625 76.075 109.795 76.245 ;
      RECT 109.165 76.075 109.335 76.245 ;
      RECT 108.705 76.075 108.875 76.245 ;
      RECT 108.245 76.075 108.415 76.245 ;
      RECT 107.785 76.075 107.955 76.245 ;
      RECT 107.325 76.075 107.495 76.245 ;
      RECT 106.865 76.075 107.035 76.245 ;
      RECT 106.405 76.075 106.575 76.245 ;
      RECT 105.945 76.075 106.115 76.245 ;
      RECT 105.485 76.075 105.655 76.245 ;
      RECT 105.025 76.075 105.195 76.245 ;
      RECT 104.565 76.075 104.735 76.245 ;
      RECT 104.105 76.075 104.275 76.245 ;
      RECT 103.645 76.075 103.815 76.245 ;
      RECT 103.185 76.075 103.355 76.245 ;
      RECT 102.725 76.075 102.895 76.245 ;
      RECT 102.265 76.075 102.435 76.245 ;
      RECT 101.805 76.075 101.975 76.245 ;
      RECT 101.345 76.075 101.515 76.245 ;
      RECT 100.885 76.075 101.055 76.245 ;
      RECT 100.425 76.075 100.595 76.245 ;
      RECT 99.965 76.075 100.135 76.245 ;
      RECT 99.505 76.075 99.675 76.245 ;
      RECT 99.045 76.075 99.215 76.245 ;
      RECT 98.585 76.075 98.755 76.245 ;
      RECT 98.125 76.075 98.295 76.245 ;
      RECT 97.665 76.075 97.835 76.245 ;
      RECT 97.205 76.075 97.375 76.245 ;
      RECT 96.745 76.075 96.915 76.245 ;
      RECT 96.285 76.075 96.455 76.245 ;
      RECT 95.825 76.075 95.995 76.245 ;
      RECT 95.365 76.075 95.535 76.245 ;
      RECT 94.905 76.075 95.075 76.245 ;
      RECT 94.445 76.075 94.615 76.245 ;
      RECT 93.985 76.075 94.155 76.245 ;
      RECT 93.525 76.075 93.695 76.245 ;
      RECT 93.065 76.075 93.235 76.245 ;
      RECT 92.605 76.075 92.775 76.245 ;
      RECT 92.145 76.075 92.315 76.245 ;
      RECT 91.685 76.075 91.855 76.245 ;
      RECT 91.225 76.075 91.395 76.245 ;
      RECT 90.765 76.075 90.935 76.245 ;
      RECT 90.305 76.075 90.475 76.245 ;
      RECT 89.845 76.075 90.015 76.245 ;
      RECT 89.385 76.075 89.555 76.245 ;
      RECT 88.925 76.075 89.095 76.245 ;
      RECT 88.465 76.075 88.635 76.245 ;
      RECT 88.005 76.075 88.175 76.245 ;
      RECT 87.545 76.075 87.715 76.245 ;
      RECT 87.085 76.075 87.255 76.245 ;
      RECT 86.625 76.075 86.795 76.245 ;
      RECT 86.165 76.075 86.335 76.245 ;
      RECT 85.705 76.075 85.875 76.245 ;
      RECT 85.245 76.075 85.415 76.245 ;
      RECT 84.785 76.075 84.955 76.245 ;
      RECT 84.325 76.075 84.495 76.245 ;
      RECT 83.865 76.075 84.035 76.245 ;
      RECT 83.405 76.075 83.575 76.245 ;
      RECT 82.945 76.075 83.115 76.245 ;
      RECT 82.485 76.075 82.655 76.245 ;
      RECT 82.025 76.075 82.195 76.245 ;
      RECT 81.565 76.075 81.735 76.245 ;
      RECT 81.105 76.075 81.275 76.245 ;
      RECT 80.645 76.075 80.815 76.245 ;
      RECT 80.185 76.075 80.355 76.245 ;
      RECT 79.725 76.075 79.895 76.245 ;
      RECT 79.265 76.075 79.435 76.245 ;
      RECT 78.805 76.075 78.975 76.245 ;
      RECT 78.345 76.075 78.515 76.245 ;
      RECT 77.885 76.075 78.055 76.245 ;
      RECT 77.425 76.075 77.595 76.245 ;
      RECT 76.965 76.075 77.135 76.245 ;
      RECT 76.505 76.075 76.675 76.245 ;
      RECT 76.045 76.075 76.215 76.245 ;
      RECT 75.585 76.075 75.755 76.245 ;
      RECT 75.125 76.075 75.295 76.245 ;
      RECT 74.665 76.075 74.835 76.245 ;
      RECT 74.205 76.075 74.375 76.245 ;
      RECT 73.745 76.075 73.915 76.245 ;
      RECT 73.285 76.075 73.455 76.245 ;
      RECT 72.825 76.075 72.995 76.245 ;
      RECT 72.365 76.075 72.535 76.245 ;
      RECT 71.905 76.075 72.075 76.245 ;
      RECT 71.445 76.075 71.615 76.245 ;
      RECT 70.985 76.075 71.155 76.245 ;
      RECT 70.525 76.075 70.695 76.245 ;
      RECT 70.065 76.075 70.235 76.245 ;
      RECT 69.605 76.075 69.775 76.245 ;
      RECT 69.145 76.075 69.315 76.245 ;
      RECT 68.685 76.075 68.855 76.245 ;
      RECT 68.225 76.075 68.395 76.245 ;
      RECT 67.765 76.075 67.935 76.245 ;
      RECT 67.305 76.075 67.475 76.245 ;
      RECT 66.845 76.075 67.015 76.245 ;
      RECT 66.385 76.075 66.555 76.245 ;
      RECT 65.925 76.075 66.095 76.245 ;
      RECT 65.465 76.075 65.635 76.245 ;
      RECT 65.005 76.075 65.175 76.245 ;
      RECT 64.545 76.075 64.715 76.245 ;
      RECT 64.085 76.075 64.255 76.245 ;
      RECT 63.625 76.075 63.795 76.245 ;
      RECT 63.165 76.075 63.335 76.245 ;
      RECT 62.705 76.075 62.875 76.245 ;
      RECT 62.245 76.075 62.415 76.245 ;
      RECT 61.785 76.075 61.955 76.245 ;
      RECT 61.325 76.075 61.495 76.245 ;
      RECT 60.865 76.075 61.035 76.245 ;
      RECT 60.405 76.075 60.575 76.245 ;
      RECT 59.945 76.075 60.115 76.245 ;
      RECT 59.485 76.075 59.655 76.245 ;
      RECT 59.025 76.075 59.195 76.245 ;
      RECT 58.565 76.075 58.735 76.245 ;
      RECT 58.105 76.075 58.275 76.245 ;
      RECT 57.645 76.075 57.815 76.245 ;
      RECT 57.185 76.075 57.355 76.245 ;
      RECT 56.725 76.075 56.895 76.245 ;
      RECT 56.265 76.075 56.435 76.245 ;
      RECT 55.805 76.075 55.975 76.245 ;
      RECT 55.345 76.075 55.515 76.245 ;
      RECT 54.885 76.075 55.055 76.245 ;
      RECT 54.425 76.075 54.595 76.245 ;
      RECT 53.965 76.075 54.135 76.245 ;
      RECT 53.505 76.075 53.675 76.245 ;
      RECT 53.045 76.075 53.215 76.245 ;
      RECT 52.585 76.075 52.755 76.245 ;
      RECT 52.125 76.075 52.295 76.245 ;
      RECT 51.665 76.075 51.835 76.245 ;
      RECT 51.205 76.075 51.375 76.245 ;
      RECT 50.745 76.075 50.915 76.245 ;
      RECT 50.285 76.075 50.455 76.245 ;
      RECT 49.825 76.075 49.995 76.245 ;
      RECT 49.365 76.075 49.535 76.245 ;
      RECT 48.905 76.075 49.075 76.245 ;
      RECT 48.445 76.075 48.615 76.245 ;
      RECT 47.985 76.075 48.155 76.245 ;
      RECT 47.525 76.075 47.695 76.245 ;
      RECT 47.065 76.075 47.235 76.245 ;
      RECT 46.605 76.075 46.775 76.245 ;
      RECT 46.145 76.075 46.315 76.245 ;
      RECT 45.685 76.075 45.855 76.245 ;
      RECT 45.225 76.075 45.395 76.245 ;
      RECT 44.765 76.075 44.935 76.245 ;
      RECT 44.305 76.075 44.475 76.245 ;
      RECT 43.845 76.075 44.015 76.245 ;
      RECT 43.385 76.075 43.555 76.245 ;
      RECT 42.925 76.075 43.095 76.245 ;
      RECT 42.465 76.075 42.635 76.245 ;
      RECT 42.005 76.075 42.175 76.245 ;
      RECT 41.545 76.075 41.715 76.245 ;
      RECT 41.085 76.075 41.255 76.245 ;
      RECT 40.625 76.075 40.795 76.245 ;
      RECT 40.165 76.075 40.335 76.245 ;
      RECT 39.705 76.075 39.875 76.245 ;
      RECT 39.245 76.075 39.415 76.245 ;
      RECT 38.785 76.075 38.955 76.245 ;
      RECT 38.325 76.075 38.495 76.245 ;
      RECT 37.865 76.075 38.035 76.245 ;
      RECT 37.405 76.075 37.575 76.245 ;
      RECT 36.945 76.075 37.115 76.245 ;
      RECT 36.485 76.075 36.655 76.245 ;
      RECT 36.025 76.075 36.195 76.245 ;
      RECT 35.565 76.075 35.735 76.245 ;
      RECT 35.105 76.075 35.275 76.245 ;
      RECT 34.645 76.075 34.815 76.245 ;
      RECT 34.185 76.075 34.355 76.245 ;
      RECT 33.725 76.075 33.895 76.245 ;
      RECT 33.265 76.075 33.435 76.245 ;
      RECT 32.805 76.075 32.975 76.245 ;
      RECT 32.345 76.075 32.515 76.245 ;
      RECT 31.885 76.075 32.055 76.245 ;
      RECT 31.425 76.075 31.595 76.245 ;
      RECT 30.965 76.075 31.135 76.245 ;
      RECT 30.505 76.075 30.675 76.245 ;
      RECT 30.045 76.075 30.215 76.245 ;
      RECT 29.585 76.075 29.755 76.245 ;
      RECT 29.125 76.075 29.295 76.245 ;
      RECT 28.665 76.075 28.835 76.245 ;
      RECT 28.205 76.075 28.375 76.245 ;
      RECT 27.745 76.075 27.915 76.245 ;
      RECT 27.285 76.075 27.455 76.245 ;
      RECT 26.825 76.075 26.995 76.245 ;
      RECT 26.365 76.075 26.535 76.245 ;
      RECT 25.905 76.075 26.075 76.245 ;
      RECT 25.445 76.075 25.615 76.245 ;
      RECT 24.985 76.075 25.155 76.245 ;
      RECT 24.525 76.075 24.695 76.245 ;
      RECT 24.065 76.075 24.235 76.245 ;
      RECT 23.605 76.075 23.775 76.245 ;
      RECT 23.145 76.075 23.315 76.245 ;
      RECT 22.685 76.075 22.855 76.245 ;
      RECT 22.225 76.075 22.395 76.245 ;
      RECT 21.765 76.075 21.935 76.245 ;
      RECT 21.305 76.075 21.475 76.245 ;
      RECT 20.845 76.075 21.015 76.245 ;
      RECT 20.385 76.075 20.555 76.245 ;
      RECT 19.925 76.075 20.095 76.245 ;
      RECT 19.465 76.075 19.635 76.245 ;
      RECT 19.005 76.075 19.175 76.245 ;
      RECT 18.545 76.075 18.715 76.245 ;
      RECT 18.085 76.075 18.255 76.245 ;
      RECT 17.625 76.075 17.795 76.245 ;
      RECT 17.165 76.075 17.335 76.245 ;
      RECT 16.705 76.075 16.875 76.245 ;
      RECT 16.245 76.075 16.415 76.245 ;
      RECT 15.785 76.075 15.955 76.245 ;
      RECT 15.325 76.075 15.495 76.245 ;
      RECT 14.865 76.075 15.035 76.245 ;
      RECT 14.405 76.075 14.575 76.245 ;
      RECT 13.945 76.075 14.115 76.245 ;
      RECT 13.485 76.075 13.655 76.245 ;
      RECT 13.025 76.075 13.195 76.245 ;
      RECT 12.565 76.075 12.735 76.245 ;
      RECT 12.105 76.075 12.275 76.245 ;
      RECT 11.645 76.075 11.815 76.245 ;
      RECT 11.185 76.075 11.355 76.245 ;
      RECT 10.725 76.075 10.895 76.245 ;
      RECT 10.265 76.075 10.435 76.245 ;
      RECT 9.805 76.075 9.975 76.245 ;
      RECT 9.345 76.075 9.515 76.245 ;
      RECT 8.885 76.075 9.055 76.245 ;
      RECT 8.425 76.075 8.595 76.245 ;
      RECT 7.965 76.075 8.135 76.245 ;
      RECT 7.505 76.075 7.675 76.245 ;
      RECT 7.045 76.075 7.215 76.245 ;
      RECT 6.585 76.075 6.755 76.245 ;
      RECT 6.125 76.075 6.295 76.245 ;
      RECT 5.665 76.075 5.835 76.245 ;
      RECT 5.205 76.075 5.375 76.245 ;
      RECT 4.745 76.075 4.915 76.245 ;
      RECT 4.285 76.075 4.455 76.245 ;
      RECT 3.825 76.075 3.995 76.245 ;
      RECT 3.365 76.075 3.535 76.245 ;
      RECT 2.905 76.075 3.075 76.245 ;
      RECT 2.445 76.075 2.615 76.245 ;
      RECT 1.985 76.075 2.155 76.245 ;
      RECT 1.525 76.075 1.695 76.245 ;
      RECT 1.065 76.075 1.235 76.245 ;
      RECT 0.605 76.075 0.775 76.245 ;
      RECT 0.145 76.075 0.315 76.245 ;
      RECT 141.365 73.355 141.535 73.525 ;
      RECT 140.905 73.355 141.075 73.525 ;
      RECT 0.605 73.355 0.775 73.525 ;
      RECT 0.145 73.355 0.315 73.525 ;
      RECT 141.365 70.635 141.535 70.805 ;
      RECT 140.905 70.635 141.075 70.805 ;
      RECT 0.605 70.635 0.775 70.805 ;
      RECT 0.145 70.635 0.315 70.805 ;
      RECT 141.365 67.915 141.535 68.085 ;
      RECT 140.905 67.915 141.075 68.085 ;
      RECT 0.605 67.915 0.775 68.085 ;
      RECT 0.145 67.915 0.315 68.085 ;
      RECT 141.365 65.195 141.535 65.365 ;
      RECT 140.905 65.195 141.075 65.365 ;
      RECT 0.605 65.195 0.775 65.365 ;
      RECT 0.145 65.195 0.315 65.365 ;
      RECT 141.365 62.475 141.535 62.645 ;
      RECT 140.905 62.475 141.075 62.645 ;
      RECT 0.605 62.475 0.775 62.645 ;
      RECT 0.145 62.475 0.315 62.645 ;
      RECT 141.365 59.755 141.535 59.925 ;
      RECT 140.905 59.755 141.075 59.925 ;
      RECT 0.605 59.755 0.775 59.925 ;
      RECT 0.145 59.755 0.315 59.925 ;
      RECT 141.365 57.035 141.535 57.205 ;
      RECT 140.905 57.035 141.075 57.205 ;
      RECT 0.605 57.035 0.775 57.205 ;
      RECT 0.145 57.035 0.315 57.205 ;
      RECT 141.365 54.315 141.535 54.485 ;
      RECT 140.905 54.315 141.075 54.485 ;
      RECT 0.605 54.315 0.775 54.485 ;
      RECT 0.145 54.315 0.315 54.485 ;
      RECT 141.365 51.595 141.535 51.765 ;
      RECT 140.905 51.595 141.075 51.765 ;
      RECT 0.605 51.595 0.775 51.765 ;
      RECT 0.145 51.595 0.315 51.765 ;
      RECT 141.365 48.875 141.535 49.045 ;
      RECT 140.905 48.875 141.075 49.045 ;
      RECT 0.605 48.875 0.775 49.045 ;
      RECT 0.145 48.875 0.315 49.045 ;
      RECT 141.365 46.155 141.535 46.325 ;
      RECT 140.905 46.155 141.075 46.325 ;
      RECT 0.605 46.155 0.775 46.325 ;
      RECT 0.145 46.155 0.315 46.325 ;
      RECT 141.365 43.435 141.535 43.605 ;
      RECT 140.905 43.435 141.075 43.605 ;
      RECT 0.605 43.435 0.775 43.605 ;
      RECT 0.145 43.435 0.315 43.605 ;
      RECT 141.365 40.715 141.535 40.885 ;
      RECT 140.905 40.715 141.075 40.885 ;
      RECT 0.605 40.715 0.775 40.885 ;
      RECT 0.145 40.715 0.315 40.885 ;
      RECT 141.365 37.995 141.535 38.165 ;
      RECT 140.905 37.995 141.075 38.165 ;
      RECT 0.605 37.995 0.775 38.165 ;
      RECT 0.145 37.995 0.315 38.165 ;
      RECT 141.365 35.275 141.535 35.445 ;
      RECT 140.905 35.275 141.075 35.445 ;
      RECT 0.605 35.275 0.775 35.445 ;
      RECT 0.145 35.275 0.315 35.445 ;
      RECT 141.365 32.555 141.535 32.725 ;
      RECT 140.905 32.555 141.075 32.725 ;
      RECT 0.605 32.555 0.775 32.725 ;
      RECT 0.145 32.555 0.315 32.725 ;
      RECT 141.365 29.835 141.535 30.005 ;
      RECT 140.905 29.835 141.075 30.005 ;
      RECT 0.605 29.835 0.775 30.005 ;
      RECT 0.145 29.835 0.315 30.005 ;
      RECT 141.365 27.115 141.535 27.285 ;
      RECT 140.905 27.115 141.075 27.285 ;
      RECT 0.605 27.115 0.775 27.285 ;
      RECT 0.145 27.115 0.315 27.285 ;
      RECT 141.365 24.395 141.535 24.565 ;
      RECT 140.905 24.395 141.075 24.565 ;
      RECT 0.605 24.395 0.775 24.565 ;
      RECT 0.145 24.395 0.315 24.565 ;
      RECT 141.365 21.675 141.535 21.845 ;
      RECT 140.905 21.675 141.075 21.845 ;
      RECT 0.605 21.675 0.775 21.845 ;
      RECT 0.145 21.675 0.315 21.845 ;
      RECT 141.365 18.955 141.535 19.125 ;
      RECT 140.905 18.955 141.075 19.125 ;
      RECT 0.605 18.955 0.775 19.125 ;
      RECT 0.145 18.955 0.315 19.125 ;
      RECT 141.365 16.235 141.535 16.405 ;
      RECT 140.905 16.235 141.075 16.405 ;
      RECT 0.605 16.235 0.775 16.405 ;
      RECT 0.145 16.235 0.315 16.405 ;
      RECT 141.365 13.515 141.535 13.685 ;
      RECT 140.905 13.515 141.075 13.685 ;
      RECT 0.605 13.515 0.775 13.685 ;
      RECT 0.145 13.515 0.315 13.685 ;
      RECT 141.365 10.795 141.535 10.965 ;
      RECT 140.905 10.795 141.075 10.965 ;
      RECT 0.605 10.795 0.775 10.965 ;
      RECT 0.145 10.795 0.315 10.965 ;
      RECT 141.365 8.075 141.535 8.245 ;
      RECT 140.905 8.075 141.075 8.245 ;
      RECT 0.605 8.075 0.775 8.245 ;
      RECT 0.145 8.075 0.315 8.245 ;
      RECT 141.365 5.355 141.535 5.525 ;
      RECT 140.905 5.355 141.075 5.525 ;
      RECT 0.605 5.355 0.775 5.525 ;
      RECT 0.145 5.355 0.315 5.525 ;
      RECT 141.365 2.635 141.535 2.805 ;
      RECT 140.905 2.635 141.075 2.805 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 141.365 -0.085 141.535 0.085 ;
      RECT 140.905 -0.085 141.075 0.085 ;
      RECT 140.445 -0.085 140.615 0.085 ;
      RECT 139.985 -0.085 140.155 0.085 ;
      RECT 139.525 -0.085 139.695 0.085 ;
      RECT 139.065 -0.085 139.235 0.085 ;
      RECT 138.605 -0.085 138.775 0.085 ;
      RECT 138.145 -0.085 138.315 0.085 ;
      RECT 137.685 -0.085 137.855 0.085 ;
      RECT 137.225 -0.085 137.395 0.085 ;
      RECT 136.765 -0.085 136.935 0.085 ;
      RECT 136.305 -0.085 136.475 0.085 ;
      RECT 135.845 -0.085 136.015 0.085 ;
      RECT 135.385 -0.085 135.555 0.085 ;
      RECT 134.925 -0.085 135.095 0.085 ;
      RECT 134.465 -0.085 134.635 0.085 ;
      RECT 134.005 -0.085 134.175 0.085 ;
      RECT 133.545 -0.085 133.715 0.085 ;
      RECT 133.085 -0.085 133.255 0.085 ;
      RECT 132.625 -0.085 132.795 0.085 ;
      RECT 132.165 -0.085 132.335 0.085 ;
      RECT 131.705 -0.085 131.875 0.085 ;
      RECT 131.245 -0.085 131.415 0.085 ;
      RECT 130.785 -0.085 130.955 0.085 ;
      RECT 130.325 -0.085 130.495 0.085 ;
      RECT 129.865 -0.085 130.035 0.085 ;
      RECT 129.405 -0.085 129.575 0.085 ;
      RECT 128.945 -0.085 129.115 0.085 ;
      RECT 128.485 -0.085 128.655 0.085 ;
      RECT 128.025 -0.085 128.195 0.085 ;
      RECT 127.565 -0.085 127.735 0.085 ;
      RECT 127.105 -0.085 127.275 0.085 ;
      RECT 126.645 -0.085 126.815 0.085 ;
      RECT 126.185 -0.085 126.355 0.085 ;
      RECT 125.725 -0.085 125.895 0.085 ;
      RECT 125.265 -0.085 125.435 0.085 ;
      RECT 124.805 -0.085 124.975 0.085 ;
      RECT 124.345 -0.085 124.515 0.085 ;
      RECT 123.885 -0.085 124.055 0.085 ;
      RECT 123.425 -0.085 123.595 0.085 ;
      RECT 122.965 -0.085 123.135 0.085 ;
      RECT 122.505 -0.085 122.675 0.085 ;
      RECT 122.045 -0.085 122.215 0.085 ;
      RECT 121.585 -0.085 121.755 0.085 ;
      RECT 121.125 -0.085 121.295 0.085 ;
      RECT 120.665 -0.085 120.835 0.085 ;
      RECT 120.205 -0.085 120.375 0.085 ;
      RECT 119.745 -0.085 119.915 0.085 ;
      RECT 119.285 -0.085 119.455 0.085 ;
      RECT 118.825 -0.085 118.995 0.085 ;
      RECT 118.365 -0.085 118.535 0.085 ;
      RECT 117.905 -0.085 118.075 0.085 ;
      RECT 117.445 -0.085 117.615 0.085 ;
      RECT 116.985 -0.085 117.155 0.085 ;
      RECT 116.525 -0.085 116.695 0.085 ;
      RECT 116.065 -0.085 116.235 0.085 ;
      RECT 115.605 -0.085 115.775 0.085 ;
      RECT 115.145 -0.085 115.315 0.085 ;
      RECT 114.685 -0.085 114.855 0.085 ;
      RECT 114.225 -0.085 114.395 0.085 ;
      RECT 113.765 -0.085 113.935 0.085 ;
      RECT 113.305 -0.085 113.475 0.085 ;
      RECT 112.845 -0.085 113.015 0.085 ;
      RECT 112.385 -0.085 112.555 0.085 ;
      RECT 111.925 -0.085 112.095 0.085 ;
      RECT 111.465 -0.085 111.635 0.085 ;
      RECT 111.005 -0.085 111.175 0.085 ;
      RECT 110.545 -0.085 110.715 0.085 ;
      RECT 110.085 -0.085 110.255 0.085 ;
      RECT 109.625 -0.085 109.795 0.085 ;
      RECT 109.165 -0.085 109.335 0.085 ;
      RECT 108.705 -0.085 108.875 0.085 ;
      RECT 108.245 -0.085 108.415 0.085 ;
      RECT 107.785 -0.085 107.955 0.085 ;
      RECT 107.325 -0.085 107.495 0.085 ;
      RECT 106.865 -0.085 107.035 0.085 ;
      RECT 106.405 -0.085 106.575 0.085 ;
      RECT 105.945 -0.085 106.115 0.085 ;
      RECT 105.485 -0.085 105.655 0.085 ;
      RECT 105.025 -0.085 105.195 0.085 ;
      RECT 104.565 -0.085 104.735 0.085 ;
      RECT 104.105 -0.085 104.275 0.085 ;
      RECT 103.645 -0.085 103.815 0.085 ;
      RECT 103.185 -0.085 103.355 0.085 ;
      RECT 102.725 -0.085 102.895 0.085 ;
      RECT 102.265 -0.085 102.435 0.085 ;
      RECT 101.805 -0.085 101.975 0.085 ;
      RECT 101.345 -0.085 101.515 0.085 ;
      RECT 100.885 -0.085 101.055 0.085 ;
      RECT 100.425 -0.085 100.595 0.085 ;
      RECT 99.965 -0.085 100.135 0.085 ;
      RECT 99.505 -0.085 99.675 0.085 ;
      RECT 99.045 -0.085 99.215 0.085 ;
      RECT 98.585 -0.085 98.755 0.085 ;
      RECT 98.125 -0.085 98.295 0.085 ;
      RECT 97.665 -0.085 97.835 0.085 ;
      RECT 97.205 -0.085 97.375 0.085 ;
      RECT 96.745 -0.085 96.915 0.085 ;
      RECT 96.285 -0.085 96.455 0.085 ;
      RECT 95.825 -0.085 95.995 0.085 ;
      RECT 95.365 -0.085 95.535 0.085 ;
      RECT 94.905 -0.085 95.075 0.085 ;
      RECT 94.445 -0.085 94.615 0.085 ;
      RECT 93.985 -0.085 94.155 0.085 ;
      RECT 93.525 -0.085 93.695 0.085 ;
      RECT 93.065 -0.085 93.235 0.085 ;
      RECT 92.605 -0.085 92.775 0.085 ;
      RECT 92.145 -0.085 92.315 0.085 ;
      RECT 91.685 -0.085 91.855 0.085 ;
      RECT 91.225 -0.085 91.395 0.085 ;
      RECT 90.765 -0.085 90.935 0.085 ;
      RECT 90.305 -0.085 90.475 0.085 ;
      RECT 89.845 -0.085 90.015 0.085 ;
      RECT 89.385 -0.085 89.555 0.085 ;
      RECT 88.925 -0.085 89.095 0.085 ;
      RECT 88.465 -0.085 88.635 0.085 ;
      RECT 88.005 -0.085 88.175 0.085 ;
      RECT 87.545 -0.085 87.715 0.085 ;
      RECT 87.085 -0.085 87.255 0.085 ;
      RECT 86.625 -0.085 86.795 0.085 ;
      RECT 86.165 -0.085 86.335 0.085 ;
      RECT 85.705 -0.085 85.875 0.085 ;
      RECT 85.245 -0.085 85.415 0.085 ;
      RECT 84.785 -0.085 84.955 0.085 ;
      RECT 84.325 -0.085 84.495 0.085 ;
      RECT 83.865 -0.085 84.035 0.085 ;
      RECT 83.405 -0.085 83.575 0.085 ;
      RECT 82.945 -0.085 83.115 0.085 ;
      RECT 82.485 -0.085 82.655 0.085 ;
      RECT 82.025 -0.085 82.195 0.085 ;
      RECT 81.565 -0.085 81.735 0.085 ;
      RECT 81.105 -0.085 81.275 0.085 ;
      RECT 80.645 -0.085 80.815 0.085 ;
      RECT 80.185 -0.085 80.355 0.085 ;
      RECT 79.725 -0.085 79.895 0.085 ;
      RECT 79.265 -0.085 79.435 0.085 ;
      RECT 78.805 -0.085 78.975 0.085 ;
      RECT 78.345 -0.085 78.515 0.085 ;
      RECT 77.885 -0.085 78.055 0.085 ;
      RECT 77.425 -0.085 77.595 0.085 ;
      RECT 76.965 -0.085 77.135 0.085 ;
      RECT 76.505 -0.085 76.675 0.085 ;
      RECT 76.045 -0.085 76.215 0.085 ;
      RECT 75.585 -0.085 75.755 0.085 ;
      RECT 75.125 -0.085 75.295 0.085 ;
      RECT 74.665 -0.085 74.835 0.085 ;
      RECT 74.205 -0.085 74.375 0.085 ;
      RECT 73.745 -0.085 73.915 0.085 ;
      RECT 73.285 -0.085 73.455 0.085 ;
      RECT 72.825 -0.085 72.995 0.085 ;
      RECT 72.365 -0.085 72.535 0.085 ;
      RECT 71.905 -0.085 72.075 0.085 ;
      RECT 71.445 -0.085 71.615 0.085 ;
      RECT 70.985 -0.085 71.155 0.085 ;
      RECT 70.525 -0.085 70.695 0.085 ;
      RECT 70.065 -0.085 70.235 0.085 ;
      RECT 69.605 -0.085 69.775 0.085 ;
      RECT 69.145 -0.085 69.315 0.085 ;
      RECT 68.685 -0.085 68.855 0.085 ;
      RECT 68.225 -0.085 68.395 0.085 ;
      RECT 67.765 -0.085 67.935 0.085 ;
      RECT 67.305 -0.085 67.475 0.085 ;
      RECT 66.845 -0.085 67.015 0.085 ;
      RECT 66.385 -0.085 66.555 0.085 ;
      RECT 65.925 -0.085 66.095 0.085 ;
      RECT 65.465 -0.085 65.635 0.085 ;
      RECT 65.005 -0.085 65.175 0.085 ;
      RECT 64.545 -0.085 64.715 0.085 ;
      RECT 64.085 -0.085 64.255 0.085 ;
      RECT 63.625 -0.085 63.795 0.085 ;
      RECT 63.165 -0.085 63.335 0.085 ;
      RECT 62.705 -0.085 62.875 0.085 ;
      RECT 62.245 -0.085 62.415 0.085 ;
      RECT 61.785 -0.085 61.955 0.085 ;
      RECT 61.325 -0.085 61.495 0.085 ;
      RECT 60.865 -0.085 61.035 0.085 ;
      RECT 60.405 -0.085 60.575 0.085 ;
      RECT 59.945 -0.085 60.115 0.085 ;
      RECT 59.485 -0.085 59.655 0.085 ;
      RECT 59.025 -0.085 59.195 0.085 ;
      RECT 58.565 -0.085 58.735 0.085 ;
      RECT 58.105 -0.085 58.275 0.085 ;
      RECT 57.645 -0.085 57.815 0.085 ;
      RECT 57.185 -0.085 57.355 0.085 ;
      RECT 56.725 -0.085 56.895 0.085 ;
      RECT 56.265 -0.085 56.435 0.085 ;
      RECT 55.805 -0.085 55.975 0.085 ;
      RECT 55.345 -0.085 55.515 0.085 ;
      RECT 54.885 -0.085 55.055 0.085 ;
      RECT 54.425 -0.085 54.595 0.085 ;
      RECT 53.965 -0.085 54.135 0.085 ;
      RECT 53.505 -0.085 53.675 0.085 ;
      RECT 53.045 -0.085 53.215 0.085 ;
      RECT 52.585 -0.085 52.755 0.085 ;
      RECT 52.125 -0.085 52.295 0.085 ;
      RECT 51.665 -0.085 51.835 0.085 ;
      RECT 51.205 -0.085 51.375 0.085 ;
      RECT 50.745 -0.085 50.915 0.085 ;
      RECT 50.285 -0.085 50.455 0.085 ;
      RECT 49.825 -0.085 49.995 0.085 ;
      RECT 49.365 -0.085 49.535 0.085 ;
      RECT 48.905 -0.085 49.075 0.085 ;
      RECT 48.445 -0.085 48.615 0.085 ;
      RECT 47.985 -0.085 48.155 0.085 ;
      RECT 47.525 -0.085 47.695 0.085 ;
      RECT 47.065 -0.085 47.235 0.085 ;
      RECT 46.605 -0.085 46.775 0.085 ;
      RECT 46.145 -0.085 46.315 0.085 ;
      RECT 45.685 -0.085 45.855 0.085 ;
      RECT 45.225 -0.085 45.395 0.085 ;
      RECT 44.765 -0.085 44.935 0.085 ;
      RECT 44.305 -0.085 44.475 0.085 ;
      RECT 43.845 -0.085 44.015 0.085 ;
      RECT 43.385 -0.085 43.555 0.085 ;
      RECT 42.925 -0.085 43.095 0.085 ;
      RECT 42.465 -0.085 42.635 0.085 ;
      RECT 42.005 -0.085 42.175 0.085 ;
      RECT 41.545 -0.085 41.715 0.085 ;
      RECT 41.085 -0.085 41.255 0.085 ;
      RECT 40.625 -0.085 40.795 0.085 ;
      RECT 40.165 -0.085 40.335 0.085 ;
      RECT 39.705 -0.085 39.875 0.085 ;
      RECT 39.245 -0.085 39.415 0.085 ;
      RECT 38.785 -0.085 38.955 0.085 ;
      RECT 38.325 -0.085 38.495 0.085 ;
      RECT 37.865 -0.085 38.035 0.085 ;
      RECT 37.405 -0.085 37.575 0.085 ;
      RECT 36.945 -0.085 37.115 0.085 ;
      RECT 36.485 -0.085 36.655 0.085 ;
      RECT 36.025 -0.085 36.195 0.085 ;
      RECT 35.565 -0.085 35.735 0.085 ;
      RECT 35.105 -0.085 35.275 0.085 ;
      RECT 34.645 -0.085 34.815 0.085 ;
      RECT 34.185 -0.085 34.355 0.085 ;
      RECT 33.725 -0.085 33.895 0.085 ;
      RECT 33.265 -0.085 33.435 0.085 ;
      RECT 32.805 -0.085 32.975 0.085 ;
      RECT 32.345 -0.085 32.515 0.085 ;
      RECT 31.885 -0.085 32.055 0.085 ;
      RECT 31.425 -0.085 31.595 0.085 ;
      RECT 30.965 -0.085 31.135 0.085 ;
      RECT 30.505 -0.085 30.675 0.085 ;
      RECT 30.045 -0.085 30.215 0.085 ;
      RECT 29.585 -0.085 29.755 0.085 ;
      RECT 29.125 -0.085 29.295 0.085 ;
      RECT 28.665 -0.085 28.835 0.085 ;
      RECT 28.205 -0.085 28.375 0.085 ;
      RECT 27.745 -0.085 27.915 0.085 ;
      RECT 27.285 -0.085 27.455 0.085 ;
      RECT 26.825 -0.085 26.995 0.085 ;
      RECT 26.365 -0.085 26.535 0.085 ;
      RECT 25.905 -0.085 26.075 0.085 ;
      RECT 25.445 -0.085 25.615 0.085 ;
      RECT 24.985 -0.085 25.155 0.085 ;
      RECT 24.525 -0.085 24.695 0.085 ;
      RECT 24.065 -0.085 24.235 0.085 ;
      RECT 23.605 -0.085 23.775 0.085 ;
      RECT 23.145 -0.085 23.315 0.085 ;
      RECT 22.685 -0.085 22.855 0.085 ;
      RECT 22.225 -0.085 22.395 0.085 ;
      RECT 21.765 -0.085 21.935 0.085 ;
      RECT 21.305 -0.085 21.475 0.085 ;
      RECT 20.845 -0.085 21.015 0.085 ;
      RECT 20.385 -0.085 20.555 0.085 ;
      RECT 19.925 -0.085 20.095 0.085 ;
      RECT 19.465 -0.085 19.635 0.085 ;
      RECT 19.005 -0.085 19.175 0.085 ;
      RECT 18.545 -0.085 18.715 0.085 ;
      RECT 18.085 -0.085 18.255 0.085 ;
      RECT 17.625 -0.085 17.795 0.085 ;
      RECT 17.165 -0.085 17.335 0.085 ;
      RECT 16.705 -0.085 16.875 0.085 ;
      RECT 16.245 -0.085 16.415 0.085 ;
      RECT 15.785 -0.085 15.955 0.085 ;
      RECT 15.325 -0.085 15.495 0.085 ;
      RECT 14.865 -0.085 15.035 0.085 ;
      RECT 14.405 -0.085 14.575 0.085 ;
      RECT 13.945 -0.085 14.115 0.085 ;
      RECT 13.485 -0.085 13.655 0.085 ;
      RECT 13.025 -0.085 13.195 0.085 ;
      RECT 12.565 -0.085 12.735 0.085 ;
      RECT 12.105 -0.085 12.275 0.085 ;
      RECT 11.645 -0.085 11.815 0.085 ;
      RECT 11.185 -0.085 11.355 0.085 ;
      RECT 10.725 -0.085 10.895 0.085 ;
      RECT 10.265 -0.085 10.435 0.085 ;
      RECT 9.805 -0.085 9.975 0.085 ;
      RECT 9.345 -0.085 9.515 0.085 ;
      RECT 8.885 -0.085 9.055 0.085 ;
      RECT 8.425 -0.085 8.595 0.085 ;
      RECT 7.965 -0.085 8.135 0.085 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.145 -0.085 0.315 0.085 ;
    LAYER via ;
      RECT 85.485 103.285 85.635 103.435 ;
      RECT 56.045 103.285 56.195 103.435 ;
      RECT 71.225 101.585 71.375 101.735 ;
      RECT 53.745 101.585 53.895 101.735 ;
      RECT 85.485 76.085 85.635 76.235 ;
      RECT 56.045 76.085 56.195 76.235 ;
      RECT 6.365 76.085 6.515 76.235 ;
      RECT 139.305 74.385 139.455 74.535 ;
      RECT 135.625 74.385 135.775 74.535 ;
      RECT 2.225 74.385 2.375 74.535 ;
      RECT 85.485 -0.075 85.635 0.075 ;
      RECT 56.045 -0.075 56.195 0.075 ;
      RECT 6.365 -0.075 6.515 0.075 ;
    LAYER via2 ;
      RECT 85.46 103.26 85.66 103.46 ;
      RECT 56.02 103.26 56.22 103.46 ;
      RECT 29.8 95.1 30 95.3 ;
      RECT 111.22 91.7 111.42 91.9 ;
      RECT 30.26 91.7 30.46 91.9 ;
      RECT 6.34 76.06 6.54 76.26 ;
      RECT 1.28 71.98 1.48 72.18 ;
      RECT 140.2 66.54 140.4 66.74 ;
      RECT 1.74 65.86 1.94 66.06 ;
      RECT 139.74 61.1 139.94 61.3 ;
      RECT 1.28 61.1 1.48 61.3 ;
      RECT 140.2 55.66 140.4 55.86 ;
      RECT 1.28 55.66 1.48 55.86 ;
      RECT 140.2 51.58 140.4 51.78 ;
      RECT 1.28 39.34 1.48 39.54 ;
      RECT 1.28 33.9 1.48 34.1 ;
      RECT 140.2 28.46 140.4 28.66 ;
      RECT 1.28 21.66 1.48 21.86 ;
      RECT 139.74 20.3 139.94 20.5 ;
      RECT 140.2 16.22 140.4 16.42 ;
      RECT 140.2 8.06 140.4 8.26 ;
      RECT 85.46 -0.1 85.66 0.1 ;
      RECT 56.02 -0.1 56.22 0.1 ;
      RECT 6.34 -0.1 6.54 0.1 ;
    LAYER via3 ;
      RECT 85.46 103.26 85.66 103.46 ;
      RECT 56.02 103.26 56.22 103.46 ;
      RECT 6.34 76.06 6.54 76.26 ;
      RECT 1.74 37.98 1.94 38.18 ;
      RECT 139.74 18.94 139.94 19.14 ;
      RECT 85.46 -0.1 85.66 0.1 ;
      RECT 56.02 -0.1 56.22 0.1 ;
      RECT 6.34 -0.1 6.54 0.1 ;
    LAYER via4 ;
      RECT 134.84 58.88 135.64 59.68 ;
      RECT 134.84 57.28 135.64 58.08 ;
      RECT 6.04 38.48 6.84 39.28 ;
      RECT 6.04 36.88 6.84 37.68 ;
      RECT 134.84 18.08 135.64 18.88 ;
      RECT 134.84 16.48 135.64 17.28 ;
    LAYER fieldpoly ;
      POLYGON 113.02 103.22 113.02 76.02 141.54 76.02 141.54 0.14 0.14 0.14 0.14 76.02 28.66 76.02 28.66 103.22 ;
    LAYER diff ;
      POLYGON 113.16 103.36 113.16 76.16 141.68 76.16 141.68 0 0 0 0 76.16 28.52 76.16 28.52 103.36 ;
    LAYER nwell ;
      POLYGON 113.35 102.055 113.35 99.225 111.13 99.225 111.13 100.45 109.29 100.45 109.29 102.055 ;
      POLYGON 32.39 102.055 32.39 100.45 30.55 100.45 30.55 99.225 28.33 99.225 28.33 102.055 ;
      POLYGON 113.35 96.615 113.35 93.785 112.05 93.785 112.05 95.01 109.29 95.01 109.29 96.615 ;
      RECT 28.33 93.785 32.39 96.615 ;
      RECT 112.51 88.345 113.35 91.175 ;
      POLYGON 30.55 91.175 30.55 89.95 32.39 89.95 32.39 88.345 28.33 88.345 28.33 91.175 ;
      RECT 112.05 82.905 113.35 85.735 ;
      RECT 28.33 82.905 32.39 85.735 ;
      POLYGON 113.35 80.295 113.35 77.465 112.51 77.465 112.51 78.69 112.05 78.69 112.05 80.295 ;
      POLYGON 32.39 80.295 32.39 78.69 30.55 78.69 30.55 77.465 28.33 77.465 28.33 80.295 ;
      POLYGON 141.87 74.855 141.87 72.025 140.57 72.025 140.57 73.25 137.81 73.25 137.81 74.855 ;
      POLYGON 3.87 74.855 3.87 73.25 2.03 73.25 2.03 72.025 -0.19 72.025 -0.19 74.855 ;
      RECT 140.57 66.585 141.87 69.415 ;
      RECT -0.19 66.585 2.03 69.415 ;
      RECT 140.57 61.145 141.87 63.975 ;
      RECT -0.19 61.145 2.03 63.975 ;
      RECT 140.57 55.705 141.87 58.535 ;
      RECT -0.19 55.705 2.03 58.535 ;
      RECT 140.57 50.265 141.87 53.095 ;
      POLYGON 3.87 53.095 3.87 51.49 2.03 51.49 2.03 50.265 -0.19 50.265 -0.19 53.095 ;
      RECT 140.57 44.825 141.87 47.655 ;
      RECT -0.19 44.825 2.03 47.655 ;
      RECT 140.57 39.385 141.87 42.215 ;
      RECT -0.19 39.385 2.03 42.215 ;
      RECT 140.57 33.945 141.87 36.775 ;
      RECT -0.19 33.945 2.03 36.775 ;
      RECT 140.57 28.505 141.87 31.335 ;
      RECT -0.19 28.505 2.03 31.335 ;
      RECT 140.57 23.065 141.87 25.895 ;
      RECT -0.19 23.065 2.03 25.895 ;
      POLYGON 141.87 20.455 141.87 17.625 139.65 17.625 139.65 19.23 140.57 19.23 140.57 20.455 ;
      RECT -0.19 17.625 2.03 20.455 ;
      POLYGON 141.87 15.015 141.87 12.185 139.65 12.185 139.65 13.41 137.81 13.41 137.81 15.015 ;
      POLYGON 3.87 15.015 3.87 13.41 2.03 13.41 2.03 12.185 -0.19 12.185 -0.19 15.015 ;
      RECT 139.65 6.745 141.87 9.575 ;
      POLYGON 2.03 9.575 2.03 8.35 3.87 8.35 3.87 6.745 -0.19 6.745 -0.19 9.575 ;
      RECT 139.65 1.305 141.87 4.135 ;
      RECT -0.19 1.305 3.87 4.135 ;
      POLYGON 113.16 103.36 113.16 76.16 141.68 76.16 141.68 0 0 0 0 76.16 28.52 76.16 28.52 103.36 ;
    LAYER pwell ;
      RECT 109.61 103.31 109.83 103.48 ;
      RECT 105.93 103.31 106.15 103.48 ;
      RECT 102.25 103.31 102.47 103.48 ;
      RECT 98.57 103.31 98.79 103.48 ;
      RECT 94.89 103.31 95.11 103.48 ;
      RECT 91.21 103.31 91.43 103.48 ;
      RECT 87.53 103.31 87.75 103.48 ;
      RECT 83.85 103.31 84.07 103.48 ;
      RECT 80.17 103.31 80.39 103.48 ;
      RECT 76.49 103.31 76.71 103.48 ;
      RECT 72.81 103.31 73.03 103.48 ;
      RECT 69.13 103.31 69.35 103.48 ;
      RECT 65.45 103.31 65.67 103.48 ;
      RECT 61.77 103.31 61.99 103.48 ;
      RECT 58.09 103.31 58.31 103.48 ;
      RECT 54.41 103.31 54.63 103.48 ;
      RECT 50.73 103.31 50.95 103.48 ;
      RECT 47.05 103.31 47.27 103.48 ;
      RECT 43.37 103.31 43.59 103.48 ;
      RECT 39.69 103.31 39.91 103.48 ;
      RECT 36.01 103.31 36.23 103.48 ;
      RECT 32.33 103.31 32.55 103.48 ;
      RECT 28.65 103.31 28.87 103.48 ;
      RECT 138.13 76.11 138.35 76.28 ;
      RECT 134.45 76.11 134.67 76.28 ;
      RECT 130.77 76.11 130.99 76.28 ;
      RECT 127.09 76.11 127.31 76.28 ;
      RECT 123.41 76.11 123.63 76.28 ;
      RECT 119.73 76.11 119.95 76.28 ;
      RECT 116.05 76.11 116.27 76.28 ;
      RECT 25.89 76.11 26.11 76.28 ;
      RECT 22.21 76.11 22.43 76.28 ;
      RECT 18.53 76.11 18.75 76.28 ;
      RECT 14.85 76.11 15.07 76.28 ;
      RECT 11.17 76.11 11.39 76.28 ;
      RECT 7.49 76.11 7.71 76.28 ;
      RECT 3.81 76.11 4.03 76.28 ;
      RECT 0.13 76.11 0.35 76.28 ;
      RECT 140.015 -0.06 140.125 0.06 ;
      RECT 136.29 -0.12 136.51 0.05 ;
      RECT 132.61 -0.12 132.83 0.05 ;
      RECT 128.93 -0.12 129.15 0.05 ;
      RECT 125.25 -0.12 125.47 0.05 ;
      RECT 121.57 -0.12 121.79 0.05 ;
      RECT 117.89 -0.12 118.11 0.05 ;
      RECT 114.21 -0.12 114.43 0.05 ;
      RECT 110.53 -0.12 110.75 0.05 ;
      RECT 106.85 -0.12 107.07 0.05 ;
      RECT 103.17 -0.12 103.39 0.05 ;
      RECT 99.49 -0.12 99.71 0.05 ;
      RECT 95.81 -0.12 96.03 0.05 ;
      RECT 92.13 -0.12 92.35 0.05 ;
      RECT 88.45 -0.12 88.67 0.05 ;
      RECT 84.77 -0.12 84.99 0.05 ;
      RECT 81.09 -0.12 81.31 0.05 ;
      RECT 77.41 -0.12 77.63 0.05 ;
      RECT 73.73 -0.12 73.95 0.05 ;
      RECT 70.05 -0.12 70.27 0.05 ;
      RECT 66.37 -0.12 66.59 0.05 ;
      RECT 62.69 -0.12 62.91 0.05 ;
      RECT 59.01 -0.12 59.23 0.05 ;
      RECT 55.33 -0.12 55.55 0.05 ;
      RECT 51.65 -0.12 51.87 0.05 ;
      RECT 47.97 -0.12 48.19 0.05 ;
      RECT 44.29 -0.12 44.51 0.05 ;
      RECT 40.61 -0.12 40.83 0.05 ;
      RECT 36.93 -0.12 37.15 0.05 ;
      RECT 33.25 -0.12 33.47 0.05 ;
      RECT 29.57 -0.12 29.79 0.05 ;
      RECT 25.89 -0.12 26.11 0.05 ;
      RECT 22.21 -0.12 22.43 0.05 ;
      RECT 18.53 -0.12 18.75 0.05 ;
      RECT 14.85 -0.12 15.07 0.05 ;
      RECT 11.17 -0.12 11.39 0.05 ;
      RECT 7.49 -0.12 7.71 0.05 ;
      RECT 3.81 -0.12 4.03 0.05 ;
      RECT 0.13 -0.12 0.35 0.05 ;
      POLYGON 113.16 103.36 113.16 76.16 141.68 76.16 141.68 0 0 0 0 76.16 28.52 76.16 28.52 103.36 ;
    LAYER OVERLAP ;
      POLYGON 0 0 0 76.16 28.52 76.16 28.52 103.36 113.16 103.36 113.16 76.16 141.68 76.16 141.68 0 ;
  END
END sb_1__0_

END LIBRARY
