//Generated from netlist by SpyDrNet
//netlist name: FPGA88_SOFA_A
module sky130_fd_sc_hd__sdfrtp_1
(
    CLK,
    D,
    RESET_B,
    SCD,
    SCE,
    Q
);

    input CLK;
    input D;
    input RESET_B;
    input SCD;
    input SCE;
    output Q;

    wire CLK;
    wire D;
    wire Q;
    wire RESET_B;
    wire SCD;
    wire SCE;

endmodule

