VERSION 5.7 ;
BUSBITCHARS "[]" ;

UNITS
  DATABASE MICRONS 1000 ;
END UNITS

MANUFACTURINGGRID 0.005 ;

LAYER li1
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.46 ;
  WIDTH 0.17 ;
END li1

LAYER mcon
  TYPE CUT ;
END mcon

LAYER met1
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.34 ;
  WIDTH 0.14 ;
END met1

LAYER via
  TYPE CUT ;
END via

LAYER met2
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.46 ;
  WIDTH 0.14 ;
END met2

LAYER via2
  TYPE CUT ;
END via2

LAYER met3
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.68 ;
  WIDTH 0.3 ;
END met3

LAYER via3
  TYPE CUT ;
END via3

LAYER met4
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.92 ;
  WIDTH 0.3 ;
END met4

LAYER via4
  TYPE CUT ;
END via4

LAYER met5
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 3.4 ;
  WIDTH 1.6 ;
END met5

LAYER nwell
  TYPE MASTERSLICE ;
END nwell

LAYER pwell
  TYPE MASTERSLICE ;
END pwell

LAYER OVERLAP
  TYPE OVERLAP ;
END OVERLAP

VIA L1M1_PR
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.145 -0.115 0.145 0.115 ;
END L1M1_PR

VIA L1M1_PR_R
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.115 -0.145 0.115 0.145 ;
END L1M1_PR_R

VIA L1M1_PR_M
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.115 -0.145 0.115 0.145 ;
END L1M1_PR_M

VIA L1M1_PR_MR
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.145 -0.115 0.145 0.115 ;
END L1M1_PR_MR

VIA L1M1_PR_C
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.145 -0.145 0.145 0.145 ;
END L1M1_PR_C

VIA M1M2_PR
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR

VIA M1M2_PR_Enc
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_Enc

VIA M1M2_PR_R
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_R

VIA M1M2_PR_R_Enc
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR_R_Enc

VIA M1M2_PR_M
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_M

VIA M1M2_PR_M_Enc
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR_M_Enc

VIA M1M2_PR_MR
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR_MR

VIA M1M2_PR_MR_Enc
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_MR_Enc

VIA M1M2_PR_C
  LAYER met1 ;
    RECT -0.16 -0.16 0.16 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.16 0.16 0.16 ;
END M1M2_PR_C

VIA M2M3_PR
  LAYER met2 ;
    RECT -0.14 -0.185 0.14 0.185 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR

VIA M2M3_PR_R
  LAYER met2 ;
    RECT -0.185 -0.14 0.185 0.14 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_R

VIA M2M3_PR_M
  LAYER met2 ;
    RECT -0.14 -0.185 0.14 0.185 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_M

VIA M2M3_PR_MR
  LAYER met2 ;
    RECT -0.185 -0.14 0.185 0.14 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_MR

VIA M2M3_PR_C
  LAYER met2 ;
    RECT -0.185 -0.185 0.185 0.185 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_C

VIA M3M4_PR
  LAYER met3 ;
    RECT -0.19 -0.16 0.19 0.16 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR

VIA M3M4_PR_R
  LAYER met3 ;
    RECT -0.16 -0.19 0.16 0.19 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_R

VIA M3M4_PR_M
  LAYER met3 ;
    RECT -0.19 -0.16 0.19 0.16 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_M

VIA M3M4_PR_MR
  LAYER met3 ;
    RECT -0.16 -0.19 0.16 0.19 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_MR

VIA M3M4_PR_C
  LAYER met3 ;
    RECT -0.19 -0.19 0.19 0.19 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_C

VIA M4M5_PR
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR

VIA M4M5_PR_R
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_R

VIA M4M5_PR_M
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_M

VIA M4M5_PR_MR
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_MR

VIA M4M5_PR_C
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_C

SITE unit
  CLASS CORE ;
  SYMMETRY Y ;
  SIZE 0.46 BY 2.72 ;
END unit

SITE unithddbl
  CLASS CORE ;
  SIZE 0.46 BY 5.44 ;
END unithddbl

MACRO sb_1__0_
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  SIZE 117.76 BY 97.92 ;
  SYMMETRY X Y ;
  PIN prog_clk[0]
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER met2 ;
        RECT 55.59 0 55.73 1.36 ;
    END
  END prog_clk[0]
  PIN chany_top_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.87 96.56 64.01 97.92 ;
    END
  END chany_top_in[0]
  PIN chany_top_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.27 96.56 59.41 97.92 ;
    END
  END chany_top_in[1]
  PIN chany_top_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 67.93 96.56 68.23 97.92 ;
    END
  END chany_top_in[2]
  PIN chany_top_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.13 96.56 78.27 97.92 ;
    END
  END chany_top_in[3]
  PIN chany_top_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.35 96.56 58.49 97.92 ;
    END
  END chany_top_in[4]
  PIN chany_top_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.93 96.56 69.07 97.92 ;
    END
  END chany_top_in[5]
  PIN chany_top_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.39 96.56 46.53 97.92 ;
    END
  END chany_top_in[6]
  PIN chany_top_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.53 96.56 73.67 97.92 ;
    END
  END chany_top_in[7]
  PIN chany_top_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.51 96.56 56.65 97.92 ;
    END
  END chany_top_in[8]
  PIN chany_top_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.21 96.56 77.35 97.92 ;
    END
  END chany_top_in[9]
  PIN chany_top_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.17 96.56 66.31 97.92 ;
    END
  END chany_top_in[10]
  PIN chany_top_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.63 96.56 43.77 97.92 ;
    END
  END chany_top_in[11]
  PIN chany_top_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 63.33 96.56 63.63 97.92 ;
    END
  END chany_top_in[12]
  PIN chany_top_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.61 96.56 49.75 97.92 ;
    END
  END chany_top_in[13]
  PIN chany_top_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.19 96.56 83.33 97.92 ;
    END
  END chany_top_in[14]
  PIN chany_top_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.47 96.56 45.61 97.92 ;
    END
  END chany_top_in[15]
  PIN chany_top_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.05 96.56 79.19 97.92 ;
    END
  END chany_top_in[16]
  PIN chany_top_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.09 96.56 67.23 97.92 ;
    END
  END chany_top_in[17]
  PIN chany_top_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.55 96.56 44.69 97.92 ;
    END
  END chany_top_in[18]
  PIN chany_top_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.65 96.56 60.79 97.92 ;
    END
  END chany_top_in[19]
  PIN top_left_grid_pin_42_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.13 85.68 9.27 87.04 ;
    END
  END top_left_grid_pin_42_[0]
  PIN top_left_grid_pin_43_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.83 85.68 6.97 87.04 ;
    END
  END top_left_grid_pin_43_[0]
  PIN top_left_grid_pin_44_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.81 85.68 12.95 87.04 ;
    END
  END top_left_grid_pin_44_[0]
  PIN top_left_grid_pin_45_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.99 96.56 28.13 97.92 ;
    END
  END top_left_grid_pin_45_[0]
  PIN top_left_grid_pin_46_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.19 85.68 14.33 87.04 ;
    END
  END top_left_grid_pin_46_[0]
  PIN top_left_grid_pin_47_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.75 85.68 7.89 87.04 ;
    END
  END top_left_grid_pin_47_[0]
  PIN top_left_grid_pin_48_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.03 85.68 16.17 87.04 ;
    END
  END top_left_grid_pin_48_[0]
  PIN top_left_grid_pin_49_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.91 96.56 29.05 97.92 ;
    END
  END top_left_grid_pin_49_[0]
  PIN chanx_right_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.38 73.29 117.76 73.59 ;
    END
  END chanx_right_in[0]
  PIN chanx_right_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.38 71.93 117.76 72.23 ;
    END
  END chanx_right_in[1]
  PIN chanx_right_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.38 9.37 117.76 9.67 ;
    END
  END chanx_right_in[2]
  PIN chanx_right_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.38 21.61 117.76 21.91 ;
    END
  END chanx_right_in[3]
  PIN chanx_right_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.38 76.01 117.76 76.31 ;
    END
  END chanx_right_in[4]
  PIN chanx_right_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.38 22.97 117.76 23.27 ;
    END
  END chanx_right_in[5]
  PIN chanx_right_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.38 42.01 117.76 42.31 ;
    END
  END chanx_right_in[6]
  PIN chanx_right_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.38 36.57 117.76 36.87 ;
    END
  END chanx_right_in[7]
  PIN chanx_right_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.38 24.33 117.76 24.63 ;
    END
  END chanx_right_in[8]
  PIN chanx_right_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.38 44.73 117.76 45.03 ;
    END
  END chanx_right_in[9]
  PIN chanx_right_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.38 54.93 117.76 55.23 ;
    END
  END chanx_right_in[10]
  PIN chanx_right_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.38 31.13 117.76 31.43 ;
    END
  END chanx_right_in[11]
  PIN chanx_right_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.38 12.09 117.76 12.39 ;
    END
  END chanx_right_in[12]
  PIN chanx_right_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.38 83.49 117.76 83.79 ;
    END
  END chanx_right_in[13]
  PIN chanx_right_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.38 77.37 117.76 77.67 ;
    END
  END chanx_right_in[14]
  PIN chanx_right_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.38 26.37 117.76 26.67 ;
    END
  END chanx_right_in[15]
  PIN chanx_right_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.38 32.49 117.76 32.79 ;
    END
  END chanx_right_in[16]
  PIN chanx_right_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.38 10.73 117.76 11.03 ;
    END
  END chanx_right_in[17]
  PIN chanx_right_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.38 35.21 117.76 35.51 ;
    END
  END chanx_right_in[18]
  PIN chanx_right_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.38 28.41 117.76 28.71 ;
    END
  END chanx_right_in[19]
  PIN right_bottom_grid_pin_1_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.38 74.65 117.76 74.95 ;
    END
  END right_bottom_grid_pin_1_[0]
  PIN right_bottom_grid_pin_3_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.38 59.69 117.76 59.99 ;
    END
  END right_bottom_grid_pin_3_[0]
  PIN right_bottom_grid_pin_5_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.38 66.49 117.76 66.79 ;
    END
  END right_bottom_grid_pin_5_[0]
  PIN right_bottom_grid_pin_7_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.38 50.17 117.76 50.47 ;
    END
  END right_bottom_grid_pin_7_[0]
  PIN right_bottom_grid_pin_9_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.38 61.73 117.76 62.03 ;
    END
  END right_bottom_grid_pin_9_[0]
  PIN right_bottom_grid_pin_11_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.38 48.81 117.76 49.11 ;
    END
  END right_bottom_grid_pin_11_[0]
  PIN chanx_left_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 11.41 1.38 11.71 ;
    END
  END chanx_left_in[0]
  PIN chanx_left_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 66.49 1.38 66.79 ;
    END
  END chanx_left_in[1]
  PIN chanx_left_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 10.05 1.38 10.35 ;
    END
  END chanx_left_in[2]
  PIN chanx_left_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 21.61 1.38 21.91 ;
    END
  END chanx_left_in[3]
  PIN chanx_left_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 78.73 1.38 79.03 ;
    END
  END chanx_left_in[4]
  PIN chanx_left_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 15.49 1.38 15.79 ;
    END
  END chanx_left_in[5]
  PIN chanx_left_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 33.17 1.38 33.47 ;
    END
  END chanx_left_in[6]
  PIN chanx_left_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 83.49 1.38 83.79 ;
    END
  END chanx_left_in[7]
  PIN chanx_left_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 25.69 1.38 25.99 ;
    END
  END chanx_left_in[8]
  PIN chanx_left_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 34.53 1.38 34.83 ;
    END
  END chanx_left_in[9]
  PIN chanx_left_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 39.29 1.38 39.59 ;
    END
  END chanx_left_in[10]
  PIN chanx_left_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 18.21 1.38 18.51 ;
    END
  END chanx_left_in[11]
  PIN chanx_left_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 76.01 1.38 76.31 ;
    END
  END chanx_left_in[12]
  PIN chanx_left_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 69.21 1.38 69.51 ;
    END
  END chanx_left_in[13]
  PIN chanx_left_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 42.01 1.38 42.31 ;
    END
  END chanx_left_in[14]
  PIN chanx_left_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 46.09 1.38 46.39 ;
    END
  END chanx_left_in[15]
  PIN chanx_left_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 29.77 1.38 30.07 ;
    END
  END chanx_left_in[16]
  PIN chanx_left_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 24.33 1.38 24.63 ;
    END
  END chanx_left_in[17]
  PIN chanx_left_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 22.97 1.38 23.27 ;
    END
  END chanx_left_in[18]
  PIN chanx_left_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 67.85 1.38 68.15 ;
    END
  END chanx_left_in[19]
  PIN left_bottom_grid_pin_1_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 63.77 1.38 64.07 ;
    END
  END left_bottom_grid_pin_1_[0]
  PIN left_bottom_grid_pin_3_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 31.13 1.38 31.43 ;
    END
  END left_bottom_grid_pin_3_[0]
  PIN left_bottom_grid_pin_5_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 43.37 1.38 43.67 ;
    END
  END left_bottom_grid_pin_5_[0]
  PIN left_bottom_grid_pin_7_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 54.25 1.38 54.55 ;
    END
  END left_bottom_grid_pin_7_[0]
  PIN left_bottom_grid_pin_9_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 61.73 1.38 62.03 ;
    END
  END left_bottom_grid_pin_9_[0]
  PIN left_bottom_grid_pin_11_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 37.25 1.38 37.55 ;
    END
  END left_bottom_grid_pin_11_[0]
  PIN ccff_head[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.38 13.45 117.76 13.75 ;
    END
  END ccff_head[0]
  PIN chany_top_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.97 96.56 80.11 97.92 ;
    END
  END chany_top_out[0]
  PIN chany_top_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.49 96.56 62.63 97.92 ;
    END
  END chany_top_out[1]
  PIN chany_top_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.31 96.56 47.45 97.92 ;
    END
  END chany_top_out[2]
  PIN chany_top_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.37 96.56 75.51 97.92 ;
    END
  END chany_top_out[3]
  PIN chany_top_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.37 96.56 52.51 97.92 ;
    END
  END chany_top_out[4]
  PIN chany_top_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.29 96.56 76.43 97.92 ;
    END
  END chany_top_out[5]
  PIN chany_top_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.43 96.56 57.57 97.92 ;
    END
  END chany_top_out[6]
  PIN chany_top_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.85 96.56 69.99 97.92 ;
    END
  END chany_top_out[7]
  PIN chany_top_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.23 96.56 48.37 97.92 ;
    END
  END chany_top_out[8]
  PIN chany_top_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.23 96.56 71.37 97.92 ;
    END
  END chany_top_out[9]
  PIN chany_top_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.57 96.56 61.71 97.92 ;
    END
  END chany_top_out[10]
  PIN chany_top_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.79 96.56 64.93 97.92 ;
    END
  END chany_top_out[11]
  PIN chany_top_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.11 96.56 84.25 97.92 ;
    END
  END chany_top_out[12]
  PIN chany_top_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.01 96.56 68.15 97.92 ;
    END
  END chany_top_out[13]
  PIN chany_top_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.43 96.56 34.57 97.92 ;
    END
  END chany_top_out[14]
  PIN chany_top_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.61 96.56 72.75 97.92 ;
    END
  END chany_top_out[15]
  PIN chany_top_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.53 96.56 50.67 97.92 ;
    END
  END chany_top_out[16]
  PIN chany_top_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.45 96.56 74.59 97.92 ;
    END
  END chany_top_out[17]
  PIN chany_top_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.29 96.56 53.43 97.92 ;
    END
  END chany_top_out[18]
  PIN chany_top_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.27 96.56 82.41 97.92 ;
    END
  END chany_top_out[19]
  PIN chanx_right_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.38 56.97 117.76 57.27 ;
    END
  END chanx_right_out[0]
  PIN chanx_right_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.38 67.85 117.76 68.15 ;
    END
  END chanx_right_out[1]
  PIN chanx_right_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.38 43.37 117.76 43.67 ;
    END
  END chanx_right_out[2]
  PIN chanx_right_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.38 80.09 117.76 80.39 ;
    END
  END chanx_right_out[3]
  PIN chanx_right_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.38 33.85 117.76 34.15 ;
    END
  END chanx_right_out[4]
  PIN chanx_right_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.38 82.13 117.76 82.43 ;
    END
  END chanx_right_out[5]
  PIN chanx_right_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.38 39.29 117.76 39.59 ;
    END
  END chanx_right_out[6]
  PIN chanx_right_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.38 53.57 117.76 53.87 ;
    END
  END chanx_right_out[7]
  PIN chanx_right_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.38 47.45 117.76 47.75 ;
    END
  END chanx_right_out[8]
  PIN chanx_right_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.38 78.73 117.76 79.03 ;
    END
  END chanx_right_out[9]
  PIN chanx_right_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.38 46.09 117.76 46.39 ;
    END
  END chanx_right_out[10]
  PIN chanx_right_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.38 69.21 117.76 69.51 ;
    END
  END chanx_right_out[11]
  PIN chanx_right_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.38 40.65 117.76 40.95 ;
    END
  END chanx_right_out[12]
  PIN chanx_right_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.38 37.93 117.76 38.23 ;
    END
  END chanx_right_out[13]
  PIN chanx_right_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.38 29.77 117.76 30.07 ;
    END
  END chanx_right_out[14]
  PIN chanx_right_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.38 52.21 117.76 52.51 ;
    END
  END chanx_right_out[15]
  PIN chanx_right_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.38 58.33 117.76 58.63 ;
    END
  END chanx_right_out[16]
  PIN chanx_right_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.38 63.09 117.76 63.39 ;
    END
  END chanx_right_out[17]
  PIN chanx_right_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.38 70.57 117.76 70.87 ;
    END
  END chanx_right_out[18]
  PIN chanx_right_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.38 65.13 117.76 65.43 ;
    END
  END chanx_right_out[19]
  PIN chanx_left_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 59.69 1.38 59.99 ;
    END
  END chanx_left_out[0]
  PIN chanx_left_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 56.29 1.38 56.59 ;
    END
  END chanx_left_out[1]
  PIN chanx_left_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 77.37 1.38 77.67 ;
    END
  END chanx_left_out[2]
  PIN chanx_left_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 80.09 1.38 80.39 ;
    END
  END chanx_left_out[3]
  PIN chanx_left_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 48.13 1.38 48.43 ;
    END
  END chanx_left_out[4]
  PIN chanx_left_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 82.13 1.38 82.43 ;
    END
  END chanx_left_out[5]
  PIN chanx_left_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 73.29 1.38 73.59 ;
    END
  END chanx_left_out[6]
  PIN chanx_left_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 58.33 1.38 58.63 ;
    END
  END chanx_left_out[7]
  PIN chanx_left_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 19.57 1.38 19.87 ;
    END
  END chanx_left_out[8]
  PIN chanx_left_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 44.73 1.38 45.03 ;
    END
  END chanx_left_out[9]
  PIN chanx_left_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 71.93 1.38 72.23 ;
    END
  END chanx_left_out[10]
  PIN chanx_left_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 70.57 1.38 70.87 ;
    END
  END chanx_left_out[11]
  PIN chanx_left_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 74.65 1.38 74.95 ;
    END
  END chanx_left_out[12]
  PIN chanx_left_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 65.13 1.38 65.43 ;
    END
  END chanx_left_out[13]
  PIN chanx_left_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 27.73 1.38 28.03 ;
    END
  END chanx_left_out[14]
  PIN chanx_left_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 49.49 1.38 49.79 ;
    END
  END chanx_left_out[15]
  PIN chanx_left_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 40.65 1.38 40.95 ;
    END
  END chanx_left_out[16]
  PIN chanx_left_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 8.69 1.38 8.99 ;
    END
  END chanx_left_out[17]
  PIN chanx_left_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 50.85 1.38 51.15 ;
    END
  END chanx_left_out[18]
  PIN chanx_left_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 52.21 1.38 52.51 ;
    END
  END chanx_left_out[19]
  PIN ccff_tail[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 16.85 1.38 17.15 ;
    END
  END ccff_tail[0]
  PIN SC_IN_TOP
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 35.89 1.38 36.19 ;
    END
  END SC_IN_TOP
  PIN SC_IN_BOT
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 58.73 96.56 59.03 97.92 ;
    END
  END SC_IN_BOT
  PIN SC_OUT_TOP
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.21 96.56 54.35 97.92 ;
    END
  END SC_OUT_TOP
  PIN SC_OUT_BOT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.39 85.68 115.53 87.04 ;
    END
  END SC_OUT_BOT
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 0.48 2.96 ;
        RECT 117.28 2.48 117.76 2.96 ;
        RECT 0 7.92 0.48 8.4 ;
        RECT 117.28 7.92 117.76 8.4 ;
        RECT 0 13.36 0.48 13.84 ;
        RECT 117.28 13.36 117.76 13.84 ;
        RECT 0 18.8 0.48 19.28 ;
        RECT 117.28 18.8 117.76 19.28 ;
        RECT 0 24.24 0.48 24.72 ;
        RECT 117.28 24.24 117.76 24.72 ;
        RECT 0 29.68 0.48 30.16 ;
        RECT 117.28 29.68 117.76 30.16 ;
        RECT 0 35.12 0.48 35.6 ;
        RECT 117.28 35.12 117.76 35.6 ;
        RECT 0 40.56 0.48 41.04 ;
        RECT 117.28 40.56 117.76 41.04 ;
        RECT 0 46 0.48 46.48 ;
        RECT 117.28 46 117.76 46.48 ;
        RECT 0 51.44 0.48 51.92 ;
        RECT 117.28 51.44 117.76 51.92 ;
        RECT 0 56.88 0.48 57.36 ;
        RECT 117.28 56.88 117.76 57.36 ;
        RECT 0 62.32 0.48 62.8 ;
        RECT 117.28 62.32 117.76 62.8 ;
        RECT 0 67.76 0.48 68.24 ;
        RECT 117.28 67.76 117.76 68.24 ;
        RECT 0 73.2 0.48 73.68 ;
        RECT 117.28 73.2 117.76 73.68 ;
        RECT 0 78.64 0.48 79.12 ;
        RECT 117.28 78.64 117.76 79.12 ;
        RECT 0 84.08 0.48 84.56 ;
        RECT 117.28 84.08 117.76 84.56 ;
        RECT 25.76 89.52 26.24 90 ;
        RECT 91.52 89.52 92 90 ;
        RECT 25.76 94.96 26.24 95.44 ;
        RECT 91.52 94.96 92 95.44 ;
      LAYER met4 ;
        RECT 36.5 0 37.1 0.6 ;
        RECT 65.94 0 66.54 0.6 ;
        RECT 106.42 0 107.02 0.6 ;
        RECT 106.42 86.44 107.02 87.04 ;
        RECT 36.5 97.32 37.1 97.92 ;
        RECT 65.94 97.32 66.54 97.92 ;
      LAYER met5 ;
        RECT 0 11.32 3.2 14.52 ;
        RECT 114.56 11.32 117.76 14.52 ;
        RECT 0 52.12 3.2 55.32 ;
        RECT 114.56 52.12 117.76 55.32 ;
    END
  END VDD
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 0 117.76 0.24 ;
        RECT 0 5.2 0.48 5.68 ;
        RECT 117.28 5.2 117.76 5.68 ;
        RECT 0 10.64 0.48 11.12 ;
        RECT 117.28 10.64 117.76 11.12 ;
        RECT 0 16.08 0.48 16.56 ;
        RECT 117.28 16.08 117.76 16.56 ;
        RECT 0 21.52 0.48 22 ;
        RECT 117.28 21.52 117.76 22 ;
        RECT 0 26.96 0.48 27.44 ;
        RECT 117.28 26.96 117.76 27.44 ;
        RECT 0 32.4 0.48 32.88 ;
        RECT 117.28 32.4 117.76 32.88 ;
        RECT 0 37.84 0.48 38.32 ;
        RECT 117.28 37.84 117.76 38.32 ;
        RECT 0 43.28 0.48 43.76 ;
        RECT 117.28 43.28 117.76 43.76 ;
        RECT 0 48.72 0.48 49.2 ;
        RECT 117.28 48.72 117.76 49.2 ;
        RECT 0 54.16 0.48 54.64 ;
        RECT 117.28 54.16 117.76 54.64 ;
        RECT 0 59.6 0.48 60.08 ;
        RECT 117.28 59.6 117.76 60.08 ;
        RECT 0 65.04 0.48 65.52 ;
        RECT 117.28 65.04 117.76 65.52 ;
        RECT 0 70.48 0.48 70.96 ;
        RECT 117.28 70.48 117.76 70.96 ;
        RECT 0 75.92 0.48 76.4 ;
        RECT 117.28 75.92 117.76 76.4 ;
        RECT 0 81.36 0.48 81.84 ;
        RECT 117.28 81.36 117.76 81.84 ;
        RECT 0 86.8 117.76 87.28 ;
        RECT 25.76 92.24 26.24 92.72 ;
        RECT 91.52 92.24 92 92.72 ;
        RECT 25.76 97.68 92 97.92 ;
      LAYER met4 ;
        RECT 10.74 0 11.34 0.6 ;
        RECT 51.22 0 51.82 0.6 ;
        RECT 80.66 0 81.26 0.6 ;
        RECT 10.74 86.44 11.34 87.04 ;
        RECT 51.22 97.32 51.82 97.92 ;
        RECT 80.66 97.32 81.26 97.92 ;
      LAYER met5 ;
        RECT 0 31.72 3.2 34.92 ;
        RECT 114.56 31.72 117.76 34.92 ;
        RECT 0 72.52 3.2 75.72 ;
        RECT 114.56 72.52 117.76 75.72 ;
    END
  END VSS
  PIN prog_clk__FEEDTHRU_1[0]
    DIRECTION OUTPUT ;
    USE CLOCK ;
    PORT
      LAYER met3 ;
        RECT 0 13.45 1.38 13.75 ;
    END
  END prog_clk__FEEDTHRU_1[0]
  PIN prog_clk__FEEDTHRU_2[0]
    DIRECTION OUTPUT ;
    USE CLOCK ;
    PORT
      LAYER met2 ;
        RECT 55.13 96.56 55.27 97.92 ;
    END
  END prog_clk__FEEDTHRU_2[0]
  OBS
    LAYER li1 ;
      RECT 25.76 97.835 92 98.005 ;
      RECT 91.54 95.115 92 95.285 ;
      RECT 25.76 95.115 29.44 95.285 ;
      RECT 91.08 92.395 92 92.565 ;
      RECT 25.76 92.395 29.44 92.565 ;
      RECT 91.08 89.675 92 89.845 ;
      RECT 25.76 89.675 29.44 89.845 ;
      RECT 89.24 86.955 117.76 87.125 ;
      RECT 0 86.955 29.44 87.125 ;
      RECT 116.84 84.235 117.76 84.405 ;
      RECT 0 84.235 3.68 84.405 ;
      RECT 116.84 81.515 117.76 81.685 ;
      RECT 0 81.515 1.84 81.685 ;
      RECT 116.84 78.795 117.76 78.965 ;
      RECT 0 78.795 1.84 78.965 ;
      RECT 116.84 76.075 117.76 76.245 ;
      RECT 0 76.075 1.84 76.245 ;
      RECT 116.84 73.355 117.76 73.525 ;
      RECT 0 73.355 1.84 73.525 ;
      RECT 116.84 70.635 117.76 70.805 ;
      RECT 0 70.635 1.84 70.805 ;
      RECT 116.84 67.915 117.76 68.085 ;
      RECT 0 67.915 1.84 68.085 ;
      RECT 116.84 65.195 117.76 65.365 ;
      RECT 0 65.195 1.84 65.365 ;
      RECT 116.84 62.475 117.76 62.645 ;
      RECT 0 62.475 1.84 62.645 ;
      RECT 116.84 59.755 117.76 59.925 ;
      RECT 0 59.755 1.84 59.925 ;
      RECT 116.84 57.035 117.76 57.205 ;
      RECT 0 57.035 1.84 57.205 ;
      RECT 116.84 54.315 117.76 54.485 ;
      RECT 0 54.315 1.84 54.485 ;
      RECT 116.84 51.595 117.76 51.765 ;
      RECT 0 51.595 1.84 51.765 ;
      RECT 116.84 48.875 117.76 49.045 ;
      RECT 0 48.875 1.84 49.045 ;
      RECT 116.84 46.155 117.76 46.325 ;
      RECT 0 46.155 1.84 46.325 ;
      RECT 116.84 43.435 117.76 43.605 ;
      RECT 0 43.435 1.84 43.605 ;
      RECT 116.84 40.715 117.76 40.885 ;
      RECT 0 40.715 3.68 40.885 ;
      RECT 114.08 37.995 117.76 38.165 ;
      RECT 0 37.995 3.68 38.165 ;
      RECT 114.08 35.275 117.76 35.445 ;
      RECT 0 35.275 3.68 35.445 ;
      RECT 116.84 32.555 117.76 32.725 ;
      RECT 0 32.555 3.68 32.725 ;
      RECT 115.92 29.835 117.76 30.005 ;
      RECT 0 29.835 3.68 30.005 ;
      RECT 115.92 27.115 117.76 27.285 ;
      RECT 0 27.115 1.84 27.285 ;
      RECT 116.84 24.395 117.76 24.565 ;
      RECT 0 24.395 3.68 24.565 ;
      RECT 117.3 21.675 117.76 21.845 ;
      RECT 0 21.675 3.68 21.845 ;
      RECT 117.3 18.955 117.76 19.125 ;
      RECT 0 18.955 1.84 19.125 ;
      RECT 117.3 16.235 117.76 16.405 ;
      RECT 0 16.235 3.68 16.405 ;
      RECT 117.3 13.515 117.76 13.685 ;
      RECT 0 13.515 3.68 13.685 ;
      RECT 117.3 10.795 117.76 10.965 ;
      RECT 0 10.795 1.84 10.965 ;
      RECT 117.3 8.075 117.76 8.245 ;
      RECT 0 8.075 3.68 8.245 ;
      RECT 115.92 5.355 117.76 5.525 ;
      RECT 0 5.355 3.68 5.525 ;
      RECT 115.92 2.635 117.76 2.805 ;
      RECT 0 2.635 3.68 2.805 ;
      RECT 0 -0.085 117.76 0.085 ;
    LAYER met2 ;
      RECT 80.82 97.735 81.1 98.105 ;
      RECT 51.38 97.735 51.66 98.105 ;
      POLYGON 74.13 96.63 74.13 96.38 74.19 96.38 74.19 96.06 73.93 96.06 73.93 96.28 73.95 96.28 73.95 96.63 ;
      RECT 78.53 96.06 78.79 96.38 ;
      RECT 64.27 96.06 64.53 96.38 ;
      RECT 55.53 96.06 55.79 96.38 ;
      RECT 10.9 86.855 11.18 87.225 ;
      RECT 80.82 -0.185 81.1 0.185 ;
      RECT 51.38 -0.185 51.66 0.185 ;
      RECT 10.9 -0.185 11.18 0.185 ;
      POLYGON 91.72 97.64 91.72 86.76 115.11 86.76 115.11 85.4 115.81 85.4 115.81 86.76 117.48 86.76 117.48 0.28 56.01 0.28 56.01 1.64 55.31 1.64 55.31 0.28 0.28 0.28 0.28 86.76 6.55 86.76 6.55 85.4 7.25 85.4 7.25 86.76 7.47 86.76 7.47 85.4 8.17 85.4 8.17 86.76 8.85 86.76 8.85 85.4 9.55 85.4 9.55 86.76 12.53 86.76 12.53 85.4 13.23 85.4 13.23 86.76 13.91 86.76 13.91 85.4 14.61 85.4 14.61 86.76 15.75 86.76 15.75 85.4 16.45 85.4 16.45 86.76 26.04 86.76 26.04 97.64 27.71 97.64 27.71 96.28 28.41 96.28 28.41 97.64 28.63 97.64 28.63 96.28 29.33 96.28 29.33 97.64 34.15 97.64 34.15 96.28 34.85 96.28 34.85 97.64 43.35 97.64 43.35 96.28 44.05 96.28 44.05 97.64 44.27 97.64 44.27 96.28 44.97 96.28 44.97 97.64 45.19 97.64 45.19 96.28 45.89 96.28 45.89 97.64 46.11 97.64 46.11 96.28 46.81 96.28 46.81 97.64 47.03 97.64 47.03 96.28 47.73 96.28 47.73 97.64 47.95 97.64 47.95 96.28 48.65 96.28 48.65 97.64 49.33 97.64 49.33 96.28 50.03 96.28 50.03 97.64 50.25 97.64 50.25 96.28 50.95 96.28 50.95 97.64 52.09 97.64 52.09 96.28 52.79 96.28 52.79 97.64 53.01 97.64 53.01 96.28 53.71 96.28 53.71 97.64 53.93 97.64 53.93 96.28 54.63 96.28 54.63 97.64 54.85 97.64 54.85 96.28 55.55 96.28 55.55 97.64 56.23 97.64 56.23 96.28 56.93 96.28 56.93 97.64 57.15 97.64 57.15 96.28 57.85 96.28 57.85 97.64 58.07 97.64 58.07 96.28 58.77 96.28 58.77 97.64 58.99 97.64 58.99 96.28 59.69 96.28 59.69 97.64 60.37 97.64 60.37 96.28 61.07 96.28 61.07 97.64 61.29 97.64 61.29 96.28 61.99 96.28 61.99 97.64 62.21 97.64 62.21 96.28 62.91 96.28 62.91 97.64 63.59 97.64 63.59 96.28 64.29 96.28 64.29 97.64 64.51 97.64 64.51 96.28 65.21 96.28 65.21 97.64 65.89 97.64 65.89 96.28 66.59 96.28 66.59 97.64 66.81 97.64 66.81 96.28 67.51 96.28 67.51 97.64 67.73 97.64 67.73 96.28 68.43 96.28 68.43 97.64 68.65 97.64 68.65 96.28 69.35 96.28 69.35 97.64 69.57 97.64 69.57 96.28 70.27 96.28 70.27 97.64 70.95 97.64 70.95 96.28 71.65 96.28 71.65 97.64 72.33 97.64 72.33 96.28 73.03 96.28 73.03 97.64 73.25 97.64 73.25 96.28 73.95 96.28 73.95 97.64 74.17 97.64 74.17 96.28 74.87 96.28 74.87 97.64 75.09 97.64 75.09 96.28 75.79 96.28 75.79 97.64 76.01 97.64 76.01 96.28 76.71 96.28 76.71 97.64 76.93 97.64 76.93 96.28 77.63 96.28 77.63 97.64 77.85 97.64 77.85 96.28 78.55 96.28 78.55 97.64 78.77 97.64 78.77 96.28 79.47 96.28 79.47 97.64 79.69 97.64 79.69 96.28 80.39 96.28 80.39 97.64 81.99 97.64 81.99 96.28 82.69 96.28 82.69 97.64 82.91 97.64 82.91 96.28 83.61 96.28 83.61 97.64 83.83 97.64 83.83 96.28 84.53 96.28 84.53 97.64 ;
    LAYER met4 ;
      POLYGON 91.6 97.52 91.6 86.64 106.02 86.64 106.02 86.04 107.42 86.04 107.42 86.64 117.36 86.64 117.36 0.4 107.42 0.4 107.42 1 106.02 1 106.02 0.4 81.66 0.4 81.66 1 80.26 1 80.26 0.4 66.94 0.4 66.94 1 65.54 1 65.54 0.4 52.22 0.4 52.22 1 50.82 1 50.82 0.4 37.5 0.4 37.5 1 36.1 1 36.1 0.4 11.74 0.4 11.74 1 10.34 1 10.34 0.4 0.4 0.4 0.4 86.64 10.34 86.64 10.34 86.04 11.74 86.04 11.74 86.64 26.16 86.64 26.16 97.52 36.1 97.52 36.1 96.92 37.5 96.92 37.5 97.52 50.82 97.52 50.82 96.92 52.22 96.92 52.22 97.52 58.33 97.52 58.33 96.16 59.43 96.16 59.43 97.52 62.93 97.52 62.93 96.16 64.03 96.16 64.03 97.52 65.54 97.52 65.54 96.92 66.94 96.92 66.94 97.52 67.53 97.52 67.53 96.16 68.63 96.16 68.63 97.52 80.26 97.52 80.26 96.92 81.66 96.92 81.66 97.52 ;
    LAYER met3 ;
      POLYGON 81.125 98.085 81.125 98.08 81.34 98.08 81.34 97.76 81.125 97.76 81.125 97.755 80.795 97.755 80.795 97.76 80.58 97.76 80.58 98.08 80.795 98.08 80.795 98.085 ;
      POLYGON 51.685 98.085 51.685 98.08 51.9 98.08 51.9 97.76 51.685 97.76 51.685 97.755 51.355 97.755 51.355 97.76 51.14 97.76 51.14 98.08 51.355 98.08 51.355 98.085 ;
      POLYGON 11.205 87.205 11.205 87.2 11.42 87.2 11.42 86.88 11.205 86.88 11.205 86.875 10.875 86.875 10.875 86.88 10.66 86.88 10.66 87.2 10.875 87.2 10.875 87.205 ;
      POLYGON 2.03 78.36 2.03 78.35 5.21 78.35 5.21 78.05 2.03 78.05 2.03 78.04 1.65 78.04 1.65 78.36 ;
      POLYGON 2.005 77.005 2.005 77 2.03 77 2.03 76.68 2.005 76.68 2.005 76.675 1.275 76.675 1.275 77.005 ;
      RECT 1.69 73.97 2.45 74.27 ;
      POLYGON 87.55 23.95 87.55 23.65 1.78 23.65 1.78 23.67 1.23 23.67 1.23 23.95 ;
      POLYGON 81.125 0.165 81.125 0.16 81.34 0.16 81.34 -0.16 81.125 -0.16 81.125 -0.165 80.795 -0.165 80.795 -0.16 80.58 -0.16 80.58 0.16 80.795 0.16 80.795 0.165 ;
      POLYGON 51.685 0.165 51.685 0.16 51.9 0.16 51.9 -0.16 51.685 -0.16 51.685 -0.165 51.355 -0.165 51.355 -0.16 51.14 -0.16 51.14 0.16 51.355 0.16 51.355 0.165 ;
      POLYGON 11.205 0.165 11.205 0.16 11.42 0.16 11.42 -0.16 11.205 -0.16 11.205 -0.165 10.875 -0.165 10.875 -0.16 10.66 -0.16 10.66 0.16 10.875 0.16 10.875 0.165 ;
      POLYGON 91.6 97.52 91.6 86.64 117.36 86.64 117.36 84.19 115.98 84.19 115.98 83.09 117.36 83.09 117.36 82.83 115.98 82.83 115.98 81.73 117.36 81.73 117.36 80.79 115.98 80.79 115.98 79.69 117.36 79.69 117.36 79.43 115.98 79.43 115.98 78.33 117.36 78.33 117.36 78.07 115.98 78.07 115.98 76.97 117.36 76.97 117.36 76.71 115.98 76.71 115.98 75.61 117.36 75.61 117.36 75.35 115.98 75.35 115.98 74.25 117.36 74.25 117.36 73.99 115.98 73.99 115.98 72.89 117.36 72.89 117.36 72.63 115.98 72.63 115.98 71.53 117.36 71.53 117.36 71.27 115.98 71.27 115.98 70.17 117.36 70.17 117.36 69.91 115.98 69.91 115.98 68.81 117.36 68.81 117.36 68.55 115.98 68.55 115.98 67.45 117.36 67.45 117.36 67.19 115.98 67.19 115.98 66.09 117.36 66.09 117.36 65.83 115.98 65.83 115.98 64.73 117.36 64.73 117.36 63.79 115.98 63.79 115.98 62.69 117.36 62.69 117.36 62.43 115.98 62.43 115.98 61.33 117.36 61.33 117.36 60.39 115.98 60.39 115.98 59.29 117.36 59.29 117.36 59.03 115.98 59.03 115.98 57.93 117.36 57.93 117.36 57.67 115.98 57.67 115.98 56.57 117.36 56.57 117.36 55.63 115.98 55.63 115.98 54.53 117.36 54.53 117.36 54.27 115.98 54.27 115.98 53.17 117.36 53.17 117.36 52.91 115.98 52.91 115.98 51.81 117.36 51.81 117.36 50.87 115.98 50.87 115.98 49.77 117.36 49.77 117.36 49.51 115.98 49.51 115.98 48.41 117.36 48.41 117.36 48.15 115.98 48.15 115.98 47.05 117.36 47.05 117.36 46.79 115.98 46.79 115.98 45.69 117.36 45.69 117.36 45.43 115.98 45.43 115.98 44.33 117.36 44.33 117.36 44.07 115.98 44.07 115.98 42.97 117.36 42.97 117.36 42.71 115.98 42.71 115.98 41.61 117.36 41.61 117.36 41.35 115.98 41.35 115.98 40.25 117.36 40.25 117.36 39.99 115.98 39.99 115.98 38.89 117.36 38.89 117.36 38.63 115.98 38.63 115.98 37.53 117.36 37.53 117.36 37.27 115.98 37.27 115.98 36.17 117.36 36.17 117.36 35.91 115.98 35.91 115.98 34.81 117.36 34.81 117.36 34.55 115.98 34.55 115.98 33.45 117.36 33.45 117.36 33.19 115.98 33.19 115.98 32.09 117.36 32.09 117.36 31.83 115.98 31.83 115.98 30.73 117.36 30.73 117.36 30.47 115.98 30.47 115.98 29.37 117.36 29.37 117.36 29.11 115.98 29.11 115.98 28.01 117.36 28.01 117.36 27.07 115.98 27.07 115.98 25.97 117.36 25.97 117.36 25.03 115.98 25.03 115.98 23.93 117.36 23.93 117.36 23.67 115.98 23.67 115.98 22.57 117.36 22.57 117.36 22.31 115.98 22.31 115.98 21.21 117.36 21.21 117.36 14.15 115.98 14.15 115.98 13.05 117.36 13.05 117.36 12.79 115.98 12.79 115.98 11.69 117.36 11.69 117.36 11.43 115.98 11.43 115.98 10.33 117.36 10.33 117.36 10.07 115.98 10.07 115.98 8.97 117.36 8.97 117.36 0.4 0.4 0.4 0.4 8.29 1.78 8.29 1.78 9.39 0.4 9.39 0.4 9.65 1.78 9.65 1.78 10.75 0.4 10.75 0.4 11.01 1.78 11.01 1.78 12.11 0.4 12.11 0.4 13.05 1.78 13.05 1.78 14.15 0.4 14.15 0.4 15.09 1.78 15.09 1.78 16.19 0.4 16.19 0.4 16.45 1.78 16.45 1.78 17.55 0.4 17.55 0.4 17.81 1.78 17.81 1.78 18.91 0.4 18.91 0.4 19.17 1.78 19.17 1.78 20.27 0.4 20.27 0.4 21.21 1.78 21.21 1.78 22.31 0.4 22.31 0.4 22.57 1.78 22.57 1.78 23.67 0.4 23.67 0.4 23.93 1.78 23.93 1.78 25.03 0.4 25.03 0.4 25.29 1.78 25.29 1.78 26.39 0.4 26.39 0.4 27.33 1.78 27.33 1.78 28.43 0.4 28.43 0.4 29.37 1.78 29.37 1.78 30.47 0.4 30.47 0.4 30.73 1.78 30.73 1.78 31.83 0.4 31.83 0.4 32.77 1.78 32.77 1.78 33.87 0.4 33.87 0.4 34.13 1.78 34.13 1.78 35.23 0.4 35.23 0.4 35.49 1.78 35.49 1.78 36.59 0.4 36.59 0.4 36.85 1.78 36.85 1.78 37.95 0.4 37.95 0.4 38.89 1.78 38.89 1.78 39.99 0.4 39.99 0.4 40.25 1.78 40.25 1.78 41.35 0.4 41.35 0.4 41.61 1.78 41.61 1.78 42.71 0.4 42.71 0.4 42.97 1.78 42.97 1.78 44.07 0.4 44.07 0.4 44.33 1.78 44.33 1.78 45.43 0.4 45.43 0.4 45.69 1.78 45.69 1.78 46.79 0.4 46.79 0.4 47.73 1.78 47.73 1.78 48.83 0.4 48.83 0.4 49.09 1.78 49.09 1.78 50.19 0.4 50.19 0.4 50.45 1.78 50.45 1.78 51.55 0.4 51.55 0.4 51.81 1.78 51.81 1.78 52.91 0.4 52.91 0.4 53.85 1.78 53.85 1.78 54.95 0.4 54.95 0.4 55.89 1.78 55.89 1.78 56.99 0.4 56.99 0.4 57.93 1.78 57.93 1.78 59.03 0.4 59.03 0.4 59.29 1.78 59.29 1.78 60.39 0.4 60.39 0.4 61.33 1.78 61.33 1.78 62.43 0.4 62.43 0.4 63.37 1.78 63.37 1.78 64.47 0.4 64.47 0.4 64.73 1.78 64.73 1.78 65.83 0.4 65.83 0.4 66.09 1.78 66.09 1.78 67.19 0.4 67.19 0.4 67.45 1.78 67.45 1.78 68.55 0.4 68.55 0.4 68.81 1.78 68.81 1.78 69.91 0.4 69.91 0.4 70.17 1.78 70.17 1.78 71.27 0.4 71.27 0.4 71.53 1.78 71.53 1.78 72.63 0.4 72.63 0.4 72.89 1.78 72.89 1.78 73.99 0.4 73.99 0.4 74.25 1.78 74.25 1.78 75.35 0.4 75.35 0.4 75.61 1.78 75.61 1.78 76.71 0.4 76.71 0.4 76.97 1.78 76.97 1.78 78.07 0.4 78.07 0.4 78.33 1.78 78.33 1.78 79.43 0.4 79.43 0.4 79.69 1.78 79.69 1.78 80.79 0.4 80.79 0.4 81.73 1.78 81.73 1.78 82.83 0.4 82.83 0.4 83.09 1.78 83.09 1.78 84.19 0.4 84.19 0.4 86.64 26.16 86.64 26.16 97.52 ;
    LAYER met5 ;
      POLYGON 90.4 96.32 90.4 85.44 116.16 85.44 116.16 77.32 112.96 77.32 112.96 70.92 116.16 70.92 116.16 56.92 112.96 56.92 112.96 50.52 116.16 50.52 116.16 36.52 112.96 36.52 112.96 30.12 116.16 30.12 116.16 16.12 112.96 16.12 112.96 9.72 116.16 9.72 116.16 1.6 1.6 1.6 1.6 9.72 4.8 9.72 4.8 16.12 1.6 16.12 1.6 30.12 4.8 30.12 4.8 36.52 1.6 36.52 1.6 50.52 4.8 50.52 4.8 56.92 1.6 56.92 1.6 70.92 4.8 70.92 4.8 77.32 1.6 77.32 1.6 85.44 27.36 85.44 27.36 96.32 ;
    LAYER met1 ;
      POLYGON 91.72 97.4 91.72 95.72 91.24 95.72 91.24 94.68 91.72 94.68 91.72 93 91.24 93 91.24 91.96 91.72 91.96 91.72 90.28 91.24 90.28 91.24 89.24 91.72 89.24 91.72 87.56 26.04 87.56 26.04 89.24 26.52 89.24 26.52 90.28 26.04 90.28 26.04 91.96 26.52 91.96 26.52 93 26.04 93 26.04 94.68 26.52 94.68 26.52 95.72 26.04 95.72 26.04 97.4 ;
      POLYGON 117.48 86.52 117.48 84.84 117 84.84 117 83.8 117.48 83.8 117.48 82.12 117 82.12 117 81.08 117.48 81.08 117.48 79.4 117 79.4 117 78.36 117.48 78.36 117.48 76.68 117 76.68 117 75.64 117.48 75.64 117.48 73.96 117 73.96 117 72.92 117.48 72.92 117.48 71.24 117 71.24 117 70.2 117.48 70.2 117.48 68.52 117 68.52 117 67.48 117.48 67.48 117.48 65.8 117 65.8 117 64.76 117.48 64.76 117.48 63.08 117 63.08 117 62.04 117.48 62.04 117.48 60.36 117 60.36 117 59.32 117.48 59.32 117.48 57.64 117 57.64 117 56.6 117.48 56.6 117.48 54.92 117 54.92 117 53.88 117.48 53.88 117.48 52.2 117 52.2 117 51.16 117.48 51.16 117.48 49.48 117 49.48 117 48.44 117.48 48.44 117.48 46.76 117 46.76 117 45.72 117.48 45.72 117.48 44.04 117 44.04 117 43 117.48 43 117.48 41.32 117 41.32 117 40.28 117.48 40.28 117.48 38.6 117 38.6 117 37.56 117.48 37.56 117.48 35.88 117 35.88 117 34.84 117.48 34.84 117.48 33.16 117 33.16 117 32.12 117.48 32.12 117.48 30.44 117 30.44 117 29.4 117.48 29.4 117.48 27.72 117 27.72 117 26.68 117.48 26.68 117.48 25 117 25 117 23.96 117.48 23.96 117.48 22.28 117 22.28 117 21.24 117.48 21.24 117.48 19.56 117 19.56 117 18.52 117.48 18.52 117.48 16.84 117 16.84 117 15.8 117.48 15.8 117.48 14.12 117 14.12 117 13.08 117.48 13.08 117.48 11.4 117 11.4 117 10.36 117.48 10.36 117.48 8.68 117 8.68 117 7.64 117.48 7.64 117.48 5.96 117 5.96 117 4.92 117.48 4.92 117.48 3.24 117 3.24 117 2.2 117.48 2.2 117.48 0.52 0.28 0.52 0.28 2.2 0.76 2.2 0.76 3.24 0.28 3.24 0.28 4.92 0.76 4.92 0.76 5.96 0.28 5.96 0.28 7.64 0.76 7.64 0.76 8.68 0.28 8.68 0.28 10.36 0.76 10.36 0.76 11.4 0.28 11.4 0.28 13.08 0.76 13.08 0.76 14.12 0.28 14.12 0.28 15.8 0.76 15.8 0.76 16.84 0.28 16.84 0.28 18.52 0.76 18.52 0.76 19.56 0.28 19.56 0.28 21.24 0.76 21.24 0.76 22.28 0.28 22.28 0.28 23.96 0.76 23.96 0.76 25 0.28 25 0.28 26.68 0.76 26.68 0.76 27.72 0.28 27.72 0.28 29.4 0.76 29.4 0.76 30.44 0.28 30.44 0.28 32.12 0.76 32.12 0.76 33.16 0.28 33.16 0.28 34.84 0.76 34.84 0.76 35.88 0.28 35.88 0.28 37.56 0.76 37.56 0.76 38.6 0.28 38.6 0.28 40.28 0.76 40.28 0.76 41.32 0.28 41.32 0.28 43 0.76 43 0.76 44.04 0.28 44.04 0.28 45.72 0.76 45.72 0.76 46.76 0.28 46.76 0.28 48.44 0.76 48.44 0.76 49.48 0.28 49.48 0.28 51.16 0.76 51.16 0.76 52.2 0.28 52.2 0.28 53.88 0.76 53.88 0.76 54.92 0.28 54.92 0.28 56.6 0.76 56.6 0.76 57.64 0.28 57.64 0.28 59.32 0.76 59.32 0.76 60.36 0.28 60.36 0.28 62.04 0.76 62.04 0.76 63.08 0.28 63.08 0.28 64.76 0.76 64.76 0.76 65.8 0.28 65.8 0.28 67.48 0.76 67.48 0.76 68.52 0.28 68.52 0.28 70.2 0.76 70.2 0.76 71.24 0.28 71.24 0.28 72.92 0.76 72.92 0.76 73.96 0.28 73.96 0.28 75.64 0.76 75.64 0.76 76.68 0.28 76.68 0.28 78.36 0.76 78.36 0.76 79.4 0.28 79.4 0.28 81.08 0.76 81.08 0.76 82.12 0.28 82.12 0.28 83.8 0.76 83.8 0.76 84.84 0.28 84.84 0.28 86.52 ;
    LAYER li1 ;
      POLYGON 91.83 97.75 91.83 86.87 117.59 86.87 117.59 0.17 0.17 0.17 0.17 86.87 25.93 86.87 25.93 97.75 ;
    LAYER mcon ;
      RECT 91.685 97.835 91.855 98.005 ;
      RECT 91.225 97.835 91.395 98.005 ;
      RECT 90.765 97.835 90.935 98.005 ;
      RECT 90.305 97.835 90.475 98.005 ;
      RECT 89.845 97.835 90.015 98.005 ;
      RECT 89.385 97.835 89.555 98.005 ;
      RECT 88.925 97.835 89.095 98.005 ;
      RECT 88.465 97.835 88.635 98.005 ;
      RECT 88.005 97.835 88.175 98.005 ;
      RECT 87.545 97.835 87.715 98.005 ;
      RECT 87.085 97.835 87.255 98.005 ;
      RECT 86.625 97.835 86.795 98.005 ;
      RECT 86.165 97.835 86.335 98.005 ;
      RECT 85.705 97.835 85.875 98.005 ;
      RECT 85.245 97.835 85.415 98.005 ;
      RECT 84.785 97.835 84.955 98.005 ;
      RECT 84.325 97.835 84.495 98.005 ;
      RECT 83.865 97.835 84.035 98.005 ;
      RECT 83.405 97.835 83.575 98.005 ;
      RECT 82.945 97.835 83.115 98.005 ;
      RECT 82.485 97.835 82.655 98.005 ;
      RECT 82.025 97.835 82.195 98.005 ;
      RECT 81.565 97.835 81.735 98.005 ;
      RECT 81.105 97.835 81.275 98.005 ;
      RECT 80.645 97.835 80.815 98.005 ;
      RECT 80.185 97.835 80.355 98.005 ;
      RECT 79.725 97.835 79.895 98.005 ;
      RECT 79.265 97.835 79.435 98.005 ;
      RECT 78.805 97.835 78.975 98.005 ;
      RECT 78.345 97.835 78.515 98.005 ;
      RECT 77.885 97.835 78.055 98.005 ;
      RECT 77.425 97.835 77.595 98.005 ;
      RECT 76.965 97.835 77.135 98.005 ;
      RECT 76.505 97.835 76.675 98.005 ;
      RECT 76.045 97.835 76.215 98.005 ;
      RECT 75.585 97.835 75.755 98.005 ;
      RECT 75.125 97.835 75.295 98.005 ;
      RECT 74.665 97.835 74.835 98.005 ;
      RECT 74.205 97.835 74.375 98.005 ;
      RECT 73.745 97.835 73.915 98.005 ;
      RECT 73.285 97.835 73.455 98.005 ;
      RECT 72.825 97.835 72.995 98.005 ;
      RECT 72.365 97.835 72.535 98.005 ;
      RECT 71.905 97.835 72.075 98.005 ;
      RECT 71.445 97.835 71.615 98.005 ;
      RECT 70.985 97.835 71.155 98.005 ;
      RECT 70.525 97.835 70.695 98.005 ;
      RECT 70.065 97.835 70.235 98.005 ;
      RECT 69.605 97.835 69.775 98.005 ;
      RECT 69.145 97.835 69.315 98.005 ;
      RECT 68.685 97.835 68.855 98.005 ;
      RECT 68.225 97.835 68.395 98.005 ;
      RECT 67.765 97.835 67.935 98.005 ;
      RECT 67.305 97.835 67.475 98.005 ;
      RECT 66.845 97.835 67.015 98.005 ;
      RECT 66.385 97.835 66.555 98.005 ;
      RECT 65.925 97.835 66.095 98.005 ;
      RECT 65.465 97.835 65.635 98.005 ;
      RECT 65.005 97.835 65.175 98.005 ;
      RECT 64.545 97.835 64.715 98.005 ;
      RECT 64.085 97.835 64.255 98.005 ;
      RECT 63.625 97.835 63.795 98.005 ;
      RECT 63.165 97.835 63.335 98.005 ;
      RECT 62.705 97.835 62.875 98.005 ;
      RECT 62.245 97.835 62.415 98.005 ;
      RECT 61.785 97.835 61.955 98.005 ;
      RECT 61.325 97.835 61.495 98.005 ;
      RECT 60.865 97.835 61.035 98.005 ;
      RECT 60.405 97.835 60.575 98.005 ;
      RECT 59.945 97.835 60.115 98.005 ;
      RECT 59.485 97.835 59.655 98.005 ;
      RECT 59.025 97.835 59.195 98.005 ;
      RECT 58.565 97.835 58.735 98.005 ;
      RECT 58.105 97.835 58.275 98.005 ;
      RECT 57.645 97.835 57.815 98.005 ;
      RECT 57.185 97.835 57.355 98.005 ;
      RECT 56.725 97.835 56.895 98.005 ;
      RECT 56.265 97.835 56.435 98.005 ;
      RECT 55.805 97.835 55.975 98.005 ;
      RECT 55.345 97.835 55.515 98.005 ;
      RECT 54.885 97.835 55.055 98.005 ;
      RECT 54.425 97.835 54.595 98.005 ;
      RECT 53.965 97.835 54.135 98.005 ;
      RECT 53.505 97.835 53.675 98.005 ;
      RECT 53.045 97.835 53.215 98.005 ;
      RECT 52.585 97.835 52.755 98.005 ;
      RECT 52.125 97.835 52.295 98.005 ;
      RECT 51.665 97.835 51.835 98.005 ;
      RECT 51.205 97.835 51.375 98.005 ;
      RECT 50.745 97.835 50.915 98.005 ;
      RECT 50.285 97.835 50.455 98.005 ;
      RECT 49.825 97.835 49.995 98.005 ;
      RECT 49.365 97.835 49.535 98.005 ;
      RECT 48.905 97.835 49.075 98.005 ;
      RECT 48.445 97.835 48.615 98.005 ;
      RECT 47.985 97.835 48.155 98.005 ;
      RECT 47.525 97.835 47.695 98.005 ;
      RECT 47.065 97.835 47.235 98.005 ;
      RECT 46.605 97.835 46.775 98.005 ;
      RECT 46.145 97.835 46.315 98.005 ;
      RECT 45.685 97.835 45.855 98.005 ;
      RECT 45.225 97.835 45.395 98.005 ;
      RECT 44.765 97.835 44.935 98.005 ;
      RECT 44.305 97.835 44.475 98.005 ;
      RECT 43.845 97.835 44.015 98.005 ;
      RECT 43.385 97.835 43.555 98.005 ;
      RECT 42.925 97.835 43.095 98.005 ;
      RECT 42.465 97.835 42.635 98.005 ;
      RECT 42.005 97.835 42.175 98.005 ;
      RECT 41.545 97.835 41.715 98.005 ;
      RECT 41.085 97.835 41.255 98.005 ;
      RECT 40.625 97.835 40.795 98.005 ;
      RECT 40.165 97.835 40.335 98.005 ;
      RECT 39.705 97.835 39.875 98.005 ;
      RECT 39.245 97.835 39.415 98.005 ;
      RECT 38.785 97.835 38.955 98.005 ;
      RECT 38.325 97.835 38.495 98.005 ;
      RECT 37.865 97.835 38.035 98.005 ;
      RECT 37.405 97.835 37.575 98.005 ;
      RECT 36.945 97.835 37.115 98.005 ;
      RECT 36.485 97.835 36.655 98.005 ;
      RECT 36.025 97.835 36.195 98.005 ;
      RECT 35.565 97.835 35.735 98.005 ;
      RECT 35.105 97.835 35.275 98.005 ;
      RECT 34.645 97.835 34.815 98.005 ;
      RECT 34.185 97.835 34.355 98.005 ;
      RECT 33.725 97.835 33.895 98.005 ;
      RECT 33.265 97.835 33.435 98.005 ;
      RECT 32.805 97.835 32.975 98.005 ;
      RECT 32.345 97.835 32.515 98.005 ;
      RECT 31.885 97.835 32.055 98.005 ;
      RECT 31.425 97.835 31.595 98.005 ;
      RECT 30.965 97.835 31.135 98.005 ;
      RECT 30.505 97.835 30.675 98.005 ;
      RECT 30.045 97.835 30.215 98.005 ;
      RECT 29.585 97.835 29.755 98.005 ;
      RECT 29.125 97.835 29.295 98.005 ;
      RECT 28.665 97.835 28.835 98.005 ;
      RECT 28.205 97.835 28.375 98.005 ;
      RECT 27.745 97.835 27.915 98.005 ;
      RECT 27.285 97.835 27.455 98.005 ;
      RECT 26.825 97.835 26.995 98.005 ;
      RECT 26.365 97.835 26.535 98.005 ;
      RECT 25.905 97.835 26.075 98.005 ;
      RECT 91.685 95.115 91.855 95.285 ;
      RECT 91.225 95.115 91.395 95.285 ;
      RECT 26.365 95.115 26.535 95.285 ;
      RECT 25.905 95.115 26.075 95.285 ;
      RECT 91.685 92.395 91.855 92.565 ;
      RECT 91.225 92.395 91.395 92.565 ;
      RECT 26.365 92.395 26.535 92.565 ;
      RECT 25.905 92.395 26.075 92.565 ;
      RECT 91.685 89.675 91.855 89.845 ;
      RECT 91.225 89.675 91.395 89.845 ;
      RECT 26.365 89.675 26.535 89.845 ;
      RECT 25.905 89.675 26.075 89.845 ;
      RECT 117.445 86.955 117.615 87.125 ;
      RECT 116.985 86.955 117.155 87.125 ;
      RECT 116.525 86.955 116.695 87.125 ;
      RECT 116.065 86.955 116.235 87.125 ;
      RECT 115.605 86.955 115.775 87.125 ;
      RECT 115.145 86.955 115.315 87.125 ;
      RECT 114.685 86.955 114.855 87.125 ;
      RECT 114.225 86.955 114.395 87.125 ;
      RECT 113.765 86.955 113.935 87.125 ;
      RECT 113.305 86.955 113.475 87.125 ;
      RECT 112.845 86.955 113.015 87.125 ;
      RECT 112.385 86.955 112.555 87.125 ;
      RECT 111.925 86.955 112.095 87.125 ;
      RECT 111.465 86.955 111.635 87.125 ;
      RECT 111.005 86.955 111.175 87.125 ;
      RECT 110.545 86.955 110.715 87.125 ;
      RECT 110.085 86.955 110.255 87.125 ;
      RECT 109.625 86.955 109.795 87.125 ;
      RECT 109.165 86.955 109.335 87.125 ;
      RECT 108.705 86.955 108.875 87.125 ;
      RECT 108.245 86.955 108.415 87.125 ;
      RECT 107.785 86.955 107.955 87.125 ;
      RECT 107.325 86.955 107.495 87.125 ;
      RECT 106.865 86.955 107.035 87.125 ;
      RECT 106.405 86.955 106.575 87.125 ;
      RECT 105.945 86.955 106.115 87.125 ;
      RECT 105.485 86.955 105.655 87.125 ;
      RECT 105.025 86.955 105.195 87.125 ;
      RECT 104.565 86.955 104.735 87.125 ;
      RECT 104.105 86.955 104.275 87.125 ;
      RECT 103.645 86.955 103.815 87.125 ;
      RECT 103.185 86.955 103.355 87.125 ;
      RECT 102.725 86.955 102.895 87.125 ;
      RECT 102.265 86.955 102.435 87.125 ;
      RECT 101.805 86.955 101.975 87.125 ;
      RECT 101.345 86.955 101.515 87.125 ;
      RECT 100.885 86.955 101.055 87.125 ;
      RECT 100.425 86.955 100.595 87.125 ;
      RECT 99.965 86.955 100.135 87.125 ;
      RECT 99.505 86.955 99.675 87.125 ;
      RECT 99.045 86.955 99.215 87.125 ;
      RECT 98.585 86.955 98.755 87.125 ;
      RECT 98.125 86.955 98.295 87.125 ;
      RECT 97.665 86.955 97.835 87.125 ;
      RECT 97.205 86.955 97.375 87.125 ;
      RECT 96.745 86.955 96.915 87.125 ;
      RECT 96.285 86.955 96.455 87.125 ;
      RECT 95.825 86.955 95.995 87.125 ;
      RECT 95.365 86.955 95.535 87.125 ;
      RECT 94.905 86.955 95.075 87.125 ;
      RECT 94.445 86.955 94.615 87.125 ;
      RECT 93.985 86.955 94.155 87.125 ;
      RECT 93.525 86.955 93.695 87.125 ;
      RECT 93.065 86.955 93.235 87.125 ;
      RECT 92.605 86.955 92.775 87.125 ;
      RECT 92.145 86.955 92.315 87.125 ;
      RECT 91.685 86.955 91.855 87.125 ;
      RECT 91.225 86.955 91.395 87.125 ;
      RECT 90.765 86.955 90.935 87.125 ;
      RECT 90.305 86.955 90.475 87.125 ;
      RECT 89.845 86.955 90.015 87.125 ;
      RECT 89.385 86.955 89.555 87.125 ;
      RECT 88.925 86.955 89.095 87.125 ;
      RECT 88.465 86.955 88.635 87.125 ;
      RECT 88.005 86.955 88.175 87.125 ;
      RECT 87.545 86.955 87.715 87.125 ;
      RECT 87.085 86.955 87.255 87.125 ;
      RECT 86.625 86.955 86.795 87.125 ;
      RECT 86.165 86.955 86.335 87.125 ;
      RECT 85.705 86.955 85.875 87.125 ;
      RECT 85.245 86.955 85.415 87.125 ;
      RECT 84.785 86.955 84.955 87.125 ;
      RECT 84.325 86.955 84.495 87.125 ;
      RECT 83.865 86.955 84.035 87.125 ;
      RECT 83.405 86.955 83.575 87.125 ;
      RECT 82.945 86.955 83.115 87.125 ;
      RECT 82.485 86.955 82.655 87.125 ;
      RECT 82.025 86.955 82.195 87.125 ;
      RECT 81.565 86.955 81.735 87.125 ;
      RECT 81.105 86.955 81.275 87.125 ;
      RECT 80.645 86.955 80.815 87.125 ;
      RECT 80.185 86.955 80.355 87.125 ;
      RECT 79.725 86.955 79.895 87.125 ;
      RECT 79.265 86.955 79.435 87.125 ;
      RECT 78.805 86.955 78.975 87.125 ;
      RECT 78.345 86.955 78.515 87.125 ;
      RECT 77.885 86.955 78.055 87.125 ;
      RECT 77.425 86.955 77.595 87.125 ;
      RECT 76.965 86.955 77.135 87.125 ;
      RECT 76.505 86.955 76.675 87.125 ;
      RECT 76.045 86.955 76.215 87.125 ;
      RECT 75.585 86.955 75.755 87.125 ;
      RECT 75.125 86.955 75.295 87.125 ;
      RECT 74.665 86.955 74.835 87.125 ;
      RECT 74.205 86.955 74.375 87.125 ;
      RECT 73.745 86.955 73.915 87.125 ;
      RECT 73.285 86.955 73.455 87.125 ;
      RECT 72.825 86.955 72.995 87.125 ;
      RECT 72.365 86.955 72.535 87.125 ;
      RECT 71.905 86.955 72.075 87.125 ;
      RECT 71.445 86.955 71.615 87.125 ;
      RECT 70.985 86.955 71.155 87.125 ;
      RECT 70.525 86.955 70.695 87.125 ;
      RECT 70.065 86.955 70.235 87.125 ;
      RECT 69.605 86.955 69.775 87.125 ;
      RECT 69.145 86.955 69.315 87.125 ;
      RECT 68.685 86.955 68.855 87.125 ;
      RECT 68.225 86.955 68.395 87.125 ;
      RECT 67.765 86.955 67.935 87.125 ;
      RECT 67.305 86.955 67.475 87.125 ;
      RECT 66.845 86.955 67.015 87.125 ;
      RECT 66.385 86.955 66.555 87.125 ;
      RECT 65.925 86.955 66.095 87.125 ;
      RECT 65.465 86.955 65.635 87.125 ;
      RECT 65.005 86.955 65.175 87.125 ;
      RECT 64.545 86.955 64.715 87.125 ;
      RECT 64.085 86.955 64.255 87.125 ;
      RECT 63.625 86.955 63.795 87.125 ;
      RECT 63.165 86.955 63.335 87.125 ;
      RECT 62.705 86.955 62.875 87.125 ;
      RECT 62.245 86.955 62.415 87.125 ;
      RECT 61.785 86.955 61.955 87.125 ;
      RECT 61.325 86.955 61.495 87.125 ;
      RECT 60.865 86.955 61.035 87.125 ;
      RECT 60.405 86.955 60.575 87.125 ;
      RECT 59.945 86.955 60.115 87.125 ;
      RECT 59.485 86.955 59.655 87.125 ;
      RECT 59.025 86.955 59.195 87.125 ;
      RECT 58.565 86.955 58.735 87.125 ;
      RECT 58.105 86.955 58.275 87.125 ;
      RECT 57.645 86.955 57.815 87.125 ;
      RECT 57.185 86.955 57.355 87.125 ;
      RECT 56.725 86.955 56.895 87.125 ;
      RECT 56.265 86.955 56.435 87.125 ;
      RECT 55.805 86.955 55.975 87.125 ;
      RECT 55.345 86.955 55.515 87.125 ;
      RECT 54.885 86.955 55.055 87.125 ;
      RECT 54.425 86.955 54.595 87.125 ;
      RECT 53.965 86.955 54.135 87.125 ;
      RECT 53.505 86.955 53.675 87.125 ;
      RECT 53.045 86.955 53.215 87.125 ;
      RECT 52.585 86.955 52.755 87.125 ;
      RECT 52.125 86.955 52.295 87.125 ;
      RECT 51.665 86.955 51.835 87.125 ;
      RECT 51.205 86.955 51.375 87.125 ;
      RECT 50.745 86.955 50.915 87.125 ;
      RECT 50.285 86.955 50.455 87.125 ;
      RECT 49.825 86.955 49.995 87.125 ;
      RECT 49.365 86.955 49.535 87.125 ;
      RECT 48.905 86.955 49.075 87.125 ;
      RECT 48.445 86.955 48.615 87.125 ;
      RECT 47.985 86.955 48.155 87.125 ;
      RECT 47.525 86.955 47.695 87.125 ;
      RECT 47.065 86.955 47.235 87.125 ;
      RECT 46.605 86.955 46.775 87.125 ;
      RECT 46.145 86.955 46.315 87.125 ;
      RECT 45.685 86.955 45.855 87.125 ;
      RECT 45.225 86.955 45.395 87.125 ;
      RECT 44.765 86.955 44.935 87.125 ;
      RECT 44.305 86.955 44.475 87.125 ;
      RECT 43.845 86.955 44.015 87.125 ;
      RECT 43.385 86.955 43.555 87.125 ;
      RECT 42.925 86.955 43.095 87.125 ;
      RECT 42.465 86.955 42.635 87.125 ;
      RECT 42.005 86.955 42.175 87.125 ;
      RECT 41.545 86.955 41.715 87.125 ;
      RECT 41.085 86.955 41.255 87.125 ;
      RECT 40.625 86.955 40.795 87.125 ;
      RECT 40.165 86.955 40.335 87.125 ;
      RECT 39.705 86.955 39.875 87.125 ;
      RECT 39.245 86.955 39.415 87.125 ;
      RECT 38.785 86.955 38.955 87.125 ;
      RECT 38.325 86.955 38.495 87.125 ;
      RECT 37.865 86.955 38.035 87.125 ;
      RECT 37.405 86.955 37.575 87.125 ;
      RECT 36.945 86.955 37.115 87.125 ;
      RECT 36.485 86.955 36.655 87.125 ;
      RECT 36.025 86.955 36.195 87.125 ;
      RECT 35.565 86.955 35.735 87.125 ;
      RECT 35.105 86.955 35.275 87.125 ;
      RECT 34.645 86.955 34.815 87.125 ;
      RECT 34.185 86.955 34.355 87.125 ;
      RECT 33.725 86.955 33.895 87.125 ;
      RECT 33.265 86.955 33.435 87.125 ;
      RECT 32.805 86.955 32.975 87.125 ;
      RECT 32.345 86.955 32.515 87.125 ;
      RECT 31.885 86.955 32.055 87.125 ;
      RECT 31.425 86.955 31.595 87.125 ;
      RECT 30.965 86.955 31.135 87.125 ;
      RECT 30.505 86.955 30.675 87.125 ;
      RECT 30.045 86.955 30.215 87.125 ;
      RECT 29.585 86.955 29.755 87.125 ;
      RECT 29.125 86.955 29.295 87.125 ;
      RECT 28.665 86.955 28.835 87.125 ;
      RECT 28.205 86.955 28.375 87.125 ;
      RECT 27.745 86.955 27.915 87.125 ;
      RECT 27.285 86.955 27.455 87.125 ;
      RECT 26.825 86.955 26.995 87.125 ;
      RECT 26.365 86.955 26.535 87.125 ;
      RECT 25.905 86.955 26.075 87.125 ;
      RECT 25.445 86.955 25.615 87.125 ;
      RECT 24.985 86.955 25.155 87.125 ;
      RECT 24.525 86.955 24.695 87.125 ;
      RECT 24.065 86.955 24.235 87.125 ;
      RECT 23.605 86.955 23.775 87.125 ;
      RECT 23.145 86.955 23.315 87.125 ;
      RECT 22.685 86.955 22.855 87.125 ;
      RECT 22.225 86.955 22.395 87.125 ;
      RECT 21.765 86.955 21.935 87.125 ;
      RECT 21.305 86.955 21.475 87.125 ;
      RECT 20.845 86.955 21.015 87.125 ;
      RECT 20.385 86.955 20.555 87.125 ;
      RECT 19.925 86.955 20.095 87.125 ;
      RECT 19.465 86.955 19.635 87.125 ;
      RECT 19.005 86.955 19.175 87.125 ;
      RECT 18.545 86.955 18.715 87.125 ;
      RECT 18.085 86.955 18.255 87.125 ;
      RECT 17.625 86.955 17.795 87.125 ;
      RECT 17.165 86.955 17.335 87.125 ;
      RECT 16.705 86.955 16.875 87.125 ;
      RECT 16.245 86.955 16.415 87.125 ;
      RECT 15.785 86.955 15.955 87.125 ;
      RECT 15.325 86.955 15.495 87.125 ;
      RECT 14.865 86.955 15.035 87.125 ;
      RECT 14.405 86.955 14.575 87.125 ;
      RECT 13.945 86.955 14.115 87.125 ;
      RECT 13.485 86.955 13.655 87.125 ;
      RECT 13.025 86.955 13.195 87.125 ;
      RECT 12.565 86.955 12.735 87.125 ;
      RECT 12.105 86.955 12.275 87.125 ;
      RECT 11.645 86.955 11.815 87.125 ;
      RECT 11.185 86.955 11.355 87.125 ;
      RECT 10.725 86.955 10.895 87.125 ;
      RECT 10.265 86.955 10.435 87.125 ;
      RECT 9.805 86.955 9.975 87.125 ;
      RECT 9.345 86.955 9.515 87.125 ;
      RECT 8.885 86.955 9.055 87.125 ;
      RECT 8.425 86.955 8.595 87.125 ;
      RECT 7.965 86.955 8.135 87.125 ;
      RECT 7.505 86.955 7.675 87.125 ;
      RECT 7.045 86.955 7.215 87.125 ;
      RECT 6.585 86.955 6.755 87.125 ;
      RECT 6.125 86.955 6.295 87.125 ;
      RECT 5.665 86.955 5.835 87.125 ;
      RECT 5.205 86.955 5.375 87.125 ;
      RECT 4.745 86.955 4.915 87.125 ;
      RECT 4.285 86.955 4.455 87.125 ;
      RECT 3.825 86.955 3.995 87.125 ;
      RECT 3.365 86.955 3.535 87.125 ;
      RECT 2.905 86.955 3.075 87.125 ;
      RECT 2.445 86.955 2.615 87.125 ;
      RECT 1.985 86.955 2.155 87.125 ;
      RECT 1.525 86.955 1.695 87.125 ;
      RECT 1.065 86.955 1.235 87.125 ;
      RECT 0.605 86.955 0.775 87.125 ;
      RECT 0.145 86.955 0.315 87.125 ;
      RECT 117.445 84.235 117.615 84.405 ;
      RECT 116.985 84.235 117.155 84.405 ;
      RECT 0.605 84.235 0.775 84.405 ;
      RECT 0.145 84.235 0.315 84.405 ;
      RECT 117.445 81.515 117.615 81.685 ;
      RECT 116.985 81.515 117.155 81.685 ;
      RECT 0.605 81.515 0.775 81.685 ;
      RECT 0.145 81.515 0.315 81.685 ;
      RECT 117.445 78.795 117.615 78.965 ;
      RECT 116.985 78.795 117.155 78.965 ;
      RECT 0.605 78.795 0.775 78.965 ;
      RECT 0.145 78.795 0.315 78.965 ;
      RECT 117.445 76.075 117.615 76.245 ;
      RECT 116.985 76.075 117.155 76.245 ;
      RECT 0.605 76.075 0.775 76.245 ;
      RECT 0.145 76.075 0.315 76.245 ;
      RECT 117.445 73.355 117.615 73.525 ;
      RECT 116.985 73.355 117.155 73.525 ;
      RECT 0.605 73.355 0.775 73.525 ;
      RECT 0.145 73.355 0.315 73.525 ;
      RECT 117.445 70.635 117.615 70.805 ;
      RECT 116.985 70.635 117.155 70.805 ;
      RECT 0.605 70.635 0.775 70.805 ;
      RECT 0.145 70.635 0.315 70.805 ;
      RECT 117.445 67.915 117.615 68.085 ;
      RECT 116.985 67.915 117.155 68.085 ;
      RECT 0.605 67.915 0.775 68.085 ;
      RECT 0.145 67.915 0.315 68.085 ;
      RECT 117.445 65.195 117.615 65.365 ;
      RECT 116.985 65.195 117.155 65.365 ;
      RECT 0.605 65.195 0.775 65.365 ;
      RECT 0.145 65.195 0.315 65.365 ;
      RECT 117.445 62.475 117.615 62.645 ;
      RECT 116.985 62.475 117.155 62.645 ;
      RECT 0.605 62.475 0.775 62.645 ;
      RECT 0.145 62.475 0.315 62.645 ;
      RECT 117.445 59.755 117.615 59.925 ;
      RECT 116.985 59.755 117.155 59.925 ;
      RECT 0.605 59.755 0.775 59.925 ;
      RECT 0.145 59.755 0.315 59.925 ;
      RECT 117.445 57.035 117.615 57.205 ;
      RECT 116.985 57.035 117.155 57.205 ;
      RECT 0.605 57.035 0.775 57.205 ;
      RECT 0.145 57.035 0.315 57.205 ;
      RECT 117.445 54.315 117.615 54.485 ;
      RECT 116.985 54.315 117.155 54.485 ;
      RECT 0.605 54.315 0.775 54.485 ;
      RECT 0.145 54.315 0.315 54.485 ;
      RECT 117.445 51.595 117.615 51.765 ;
      RECT 116.985 51.595 117.155 51.765 ;
      RECT 0.605 51.595 0.775 51.765 ;
      RECT 0.145 51.595 0.315 51.765 ;
      RECT 117.445 48.875 117.615 49.045 ;
      RECT 116.985 48.875 117.155 49.045 ;
      RECT 0.605 48.875 0.775 49.045 ;
      RECT 0.145 48.875 0.315 49.045 ;
      RECT 117.445 46.155 117.615 46.325 ;
      RECT 116.985 46.155 117.155 46.325 ;
      RECT 0.605 46.155 0.775 46.325 ;
      RECT 0.145 46.155 0.315 46.325 ;
      RECT 117.445 43.435 117.615 43.605 ;
      RECT 116.985 43.435 117.155 43.605 ;
      RECT 0.605 43.435 0.775 43.605 ;
      RECT 0.145 43.435 0.315 43.605 ;
      RECT 117.445 40.715 117.615 40.885 ;
      RECT 116.985 40.715 117.155 40.885 ;
      RECT 0.605 40.715 0.775 40.885 ;
      RECT 0.145 40.715 0.315 40.885 ;
      RECT 117.445 37.995 117.615 38.165 ;
      RECT 116.985 37.995 117.155 38.165 ;
      RECT 0.605 37.995 0.775 38.165 ;
      RECT 0.145 37.995 0.315 38.165 ;
      RECT 117.445 35.275 117.615 35.445 ;
      RECT 116.985 35.275 117.155 35.445 ;
      RECT 0.605 35.275 0.775 35.445 ;
      RECT 0.145 35.275 0.315 35.445 ;
      RECT 117.445 32.555 117.615 32.725 ;
      RECT 116.985 32.555 117.155 32.725 ;
      RECT 0.605 32.555 0.775 32.725 ;
      RECT 0.145 32.555 0.315 32.725 ;
      RECT 117.445 29.835 117.615 30.005 ;
      RECT 116.985 29.835 117.155 30.005 ;
      RECT 0.605 29.835 0.775 30.005 ;
      RECT 0.145 29.835 0.315 30.005 ;
      RECT 117.445 27.115 117.615 27.285 ;
      RECT 116.985 27.115 117.155 27.285 ;
      RECT 0.605 27.115 0.775 27.285 ;
      RECT 0.145 27.115 0.315 27.285 ;
      RECT 117.445 24.395 117.615 24.565 ;
      RECT 116.985 24.395 117.155 24.565 ;
      RECT 0.605 24.395 0.775 24.565 ;
      RECT 0.145 24.395 0.315 24.565 ;
      RECT 117.445 21.675 117.615 21.845 ;
      RECT 116.985 21.675 117.155 21.845 ;
      RECT 0.605 21.675 0.775 21.845 ;
      RECT 0.145 21.675 0.315 21.845 ;
      RECT 117.445 18.955 117.615 19.125 ;
      RECT 116.985 18.955 117.155 19.125 ;
      RECT 0.605 18.955 0.775 19.125 ;
      RECT 0.145 18.955 0.315 19.125 ;
      RECT 117.445 16.235 117.615 16.405 ;
      RECT 116.985 16.235 117.155 16.405 ;
      RECT 0.605 16.235 0.775 16.405 ;
      RECT 0.145 16.235 0.315 16.405 ;
      RECT 117.445 13.515 117.615 13.685 ;
      RECT 116.985 13.515 117.155 13.685 ;
      RECT 0.605 13.515 0.775 13.685 ;
      RECT 0.145 13.515 0.315 13.685 ;
      RECT 117.445 10.795 117.615 10.965 ;
      RECT 116.985 10.795 117.155 10.965 ;
      RECT 0.605 10.795 0.775 10.965 ;
      RECT 0.145 10.795 0.315 10.965 ;
      RECT 117.445 8.075 117.615 8.245 ;
      RECT 116.985 8.075 117.155 8.245 ;
      RECT 0.605 8.075 0.775 8.245 ;
      RECT 0.145 8.075 0.315 8.245 ;
      RECT 117.445 5.355 117.615 5.525 ;
      RECT 116.985 5.355 117.155 5.525 ;
      RECT 0.605 5.355 0.775 5.525 ;
      RECT 0.145 5.355 0.315 5.525 ;
      RECT 117.445 2.635 117.615 2.805 ;
      RECT 116.985 2.635 117.155 2.805 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 117.445 -0.085 117.615 0.085 ;
      RECT 116.985 -0.085 117.155 0.085 ;
      RECT 116.525 -0.085 116.695 0.085 ;
      RECT 116.065 -0.085 116.235 0.085 ;
      RECT 115.605 -0.085 115.775 0.085 ;
      RECT 115.145 -0.085 115.315 0.085 ;
      RECT 114.685 -0.085 114.855 0.085 ;
      RECT 114.225 -0.085 114.395 0.085 ;
      RECT 113.765 -0.085 113.935 0.085 ;
      RECT 113.305 -0.085 113.475 0.085 ;
      RECT 112.845 -0.085 113.015 0.085 ;
      RECT 112.385 -0.085 112.555 0.085 ;
      RECT 111.925 -0.085 112.095 0.085 ;
      RECT 111.465 -0.085 111.635 0.085 ;
      RECT 111.005 -0.085 111.175 0.085 ;
      RECT 110.545 -0.085 110.715 0.085 ;
      RECT 110.085 -0.085 110.255 0.085 ;
      RECT 109.625 -0.085 109.795 0.085 ;
      RECT 109.165 -0.085 109.335 0.085 ;
      RECT 108.705 -0.085 108.875 0.085 ;
      RECT 108.245 -0.085 108.415 0.085 ;
      RECT 107.785 -0.085 107.955 0.085 ;
      RECT 107.325 -0.085 107.495 0.085 ;
      RECT 106.865 -0.085 107.035 0.085 ;
      RECT 106.405 -0.085 106.575 0.085 ;
      RECT 105.945 -0.085 106.115 0.085 ;
      RECT 105.485 -0.085 105.655 0.085 ;
      RECT 105.025 -0.085 105.195 0.085 ;
      RECT 104.565 -0.085 104.735 0.085 ;
      RECT 104.105 -0.085 104.275 0.085 ;
      RECT 103.645 -0.085 103.815 0.085 ;
      RECT 103.185 -0.085 103.355 0.085 ;
      RECT 102.725 -0.085 102.895 0.085 ;
      RECT 102.265 -0.085 102.435 0.085 ;
      RECT 101.805 -0.085 101.975 0.085 ;
      RECT 101.345 -0.085 101.515 0.085 ;
      RECT 100.885 -0.085 101.055 0.085 ;
      RECT 100.425 -0.085 100.595 0.085 ;
      RECT 99.965 -0.085 100.135 0.085 ;
      RECT 99.505 -0.085 99.675 0.085 ;
      RECT 99.045 -0.085 99.215 0.085 ;
      RECT 98.585 -0.085 98.755 0.085 ;
      RECT 98.125 -0.085 98.295 0.085 ;
      RECT 97.665 -0.085 97.835 0.085 ;
      RECT 97.205 -0.085 97.375 0.085 ;
      RECT 96.745 -0.085 96.915 0.085 ;
      RECT 96.285 -0.085 96.455 0.085 ;
      RECT 95.825 -0.085 95.995 0.085 ;
      RECT 95.365 -0.085 95.535 0.085 ;
      RECT 94.905 -0.085 95.075 0.085 ;
      RECT 94.445 -0.085 94.615 0.085 ;
      RECT 93.985 -0.085 94.155 0.085 ;
      RECT 93.525 -0.085 93.695 0.085 ;
      RECT 93.065 -0.085 93.235 0.085 ;
      RECT 92.605 -0.085 92.775 0.085 ;
      RECT 92.145 -0.085 92.315 0.085 ;
      RECT 91.685 -0.085 91.855 0.085 ;
      RECT 91.225 -0.085 91.395 0.085 ;
      RECT 90.765 -0.085 90.935 0.085 ;
      RECT 90.305 -0.085 90.475 0.085 ;
      RECT 89.845 -0.085 90.015 0.085 ;
      RECT 89.385 -0.085 89.555 0.085 ;
      RECT 88.925 -0.085 89.095 0.085 ;
      RECT 88.465 -0.085 88.635 0.085 ;
      RECT 88.005 -0.085 88.175 0.085 ;
      RECT 87.545 -0.085 87.715 0.085 ;
      RECT 87.085 -0.085 87.255 0.085 ;
      RECT 86.625 -0.085 86.795 0.085 ;
      RECT 86.165 -0.085 86.335 0.085 ;
      RECT 85.705 -0.085 85.875 0.085 ;
      RECT 85.245 -0.085 85.415 0.085 ;
      RECT 84.785 -0.085 84.955 0.085 ;
      RECT 84.325 -0.085 84.495 0.085 ;
      RECT 83.865 -0.085 84.035 0.085 ;
      RECT 83.405 -0.085 83.575 0.085 ;
      RECT 82.945 -0.085 83.115 0.085 ;
      RECT 82.485 -0.085 82.655 0.085 ;
      RECT 82.025 -0.085 82.195 0.085 ;
      RECT 81.565 -0.085 81.735 0.085 ;
      RECT 81.105 -0.085 81.275 0.085 ;
      RECT 80.645 -0.085 80.815 0.085 ;
      RECT 80.185 -0.085 80.355 0.085 ;
      RECT 79.725 -0.085 79.895 0.085 ;
      RECT 79.265 -0.085 79.435 0.085 ;
      RECT 78.805 -0.085 78.975 0.085 ;
      RECT 78.345 -0.085 78.515 0.085 ;
      RECT 77.885 -0.085 78.055 0.085 ;
      RECT 77.425 -0.085 77.595 0.085 ;
      RECT 76.965 -0.085 77.135 0.085 ;
      RECT 76.505 -0.085 76.675 0.085 ;
      RECT 76.045 -0.085 76.215 0.085 ;
      RECT 75.585 -0.085 75.755 0.085 ;
      RECT 75.125 -0.085 75.295 0.085 ;
      RECT 74.665 -0.085 74.835 0.085 ;
      RECT 74.205 -0.085 74.375 0.085 ;
      RECT 73.745 -0.085 73.915 0.085 ;
      RECT 73.285 -0.085 73.455 0.085 ;
      RECT 72.825 -0.085 72.995 0.085 ;
      RECT 72.365 -0.085 72.535 0.085 ;
      RECT 71.905 -0.085 72.075 0.085 ;
      RECT 71.445 -0.085 71.615 0.085 ;
      RECT 70.985 -0.085 71.155 0.085 ;
      RECT 70.525 -0.085 70.695 0.085 ;
      RECT 70.065 -0.085 70.235 0.085 ;
      RECT 69.605 -0.085 69.775 0.085 ;
      RECT 69.145 -0.085 69.315 0.085 ;
      RECT 68.685 -0.085 68.855 0.085 ;
      RECT 68.225 -0.085 68.395 0.085 ;
      RECT 67.765 -0.085 67.935 0.085 ;
      RECT 67.305 -0.085 67.475 0.085 ;
      RECT 66.845 -0.085 67.015 0.085 ;
      RECT 66.385 -0.085 66.555 0.085 ;
      RECT 65.925 -0.085 66.095 0.085 ;
      RECT 65.465 -0.085 65.635 0.085 ;
      RECT 65.005 -0.085 65.175 0.085 ;
      RECT 64.545 -0.085 64.715 0.085 ;
      RECT 64.085 -0.085 64.255 0.085 ;
      RECT 63.625 -0.085 63.795 0.085 ;
      RECT 63.165 -0.085 63.335 0.085 ;
      RECT 62.705 -0.085 62.875 0.085 ;
      RECT 62.245 -0.085 62.415 0.085 ;
      RECT 61.785 -0.085 61.955 0.085 ;
      RECT 61.325 -0.085 61.495 0.085 ;
      RECT 60.865 -0.085 61.035 0.085 ;
      RECT 60.405 -0.085 60.575 0.085 ;
      RECT 59.945 -0.085 60.115 0.085 ;
      RECT 59.485 -0.085 59.655 0.085 ;
      RECT 59.025 -0.085 59.195 0.085 ;
      RECT 58.565 -0.085 58.735 0.085 ;
      RECT 58.105 -0.085 58.275 0.085 ;
      RECT 57.645 -0.085 57.815 0.085 ;
      RECT 57.185 -0.085 57.355 0.085 ;
      RECT 56.725 -0.085 56.895 0.085 ;
      RECT 56.265 -0.085 56.435 0.085 ;
      RECT 55.805 -0.085 55.975 0.085 ;
      RECT 55.345 -0.085 55.515 0.085 ;
      RECT 54.885 -0.085 55.055 0.085 ;
      RECT 54.425 -0.085 54.595 0.085 ;
      RECT 53.965 -0.085 54.135 0.085 ;
      RECT 53.505 -0.085 53.675 0.085 ;
      RECT 53.045 -0.085 53.215 0.085 ;
      RECT 52.585 -0.085 52.755 0.085 ;
      RECT 52.125 -0.085 52.295 0.085 ;
      RECT 51.665 -0.085 51.835 0.085 ;
      RECT 51.205 -0.085 51.375 0.085 ;
      RECT 50.745 -0.085 50.915 0.085 ;
      RECT 50.285 -0.085 50.455 0.085 ;
      RECT 49.825 -0.085 49.995 0.085 ;
      RECT 49.365 -0.085 49.535 0.085 ;
      RECT 48.905 -0.085 49.075 0.085 ;
      RECT 48.445 -0.085 48.615 0.085 ;
      RECT 47.985 -0.085 48.155 0.085 ;
      RECT 47.525 -0.085 47.695 0.085 ;
      RECT 47.065 -0.085 47.235 0.085 ;
      RECT 46.605 -0.085 46.775 0.085 ;
      RECT 46.145 -0.085 46.315 0.085 ;
      RECT 45.685 -0.085 45.855 0.085 ;
      RECT 45.225 -0.085 45.395 0.085 ;
      RECT 44.765 -0.085 44.935 0.085 ;
      RECT 44.305 -0.085 44.475 0.085 ;
      RECT 43.845 -0.085 44.015 0.085 ;
      RECT 43.385 -0.085 43.555 0.085 ;
      RECT 42.925 -0.085 43.095 0.085 ;
      RECT 42.465 -0.085 42.635 0.085 ;
      RECT 42.005 -0.085 42.175 0.085 ;
      RECT 41.545 -0.085 41.715 0.085 ;
      RECT 41.085 -0.085 41.255 0.085 ;
      RECT 40.625 -0.085 40.795 0.085 ;
      RECT 40.165 -0.085 40.335 0.085 ;
      RECT 39.705 -0.085 39.875 0.085 ;
      RECT 39.245 -0.085 39.415 0.085 ;
      RECT 38.785 -0.085 38.955 0.085 ;
      RECT 38.325 -0.085 38.495 0.085 ;
      RECT 37.865 -0.085 38.035 0.085 ;
      RECT 37.405 -0.085 37.575 0.085 ;
      RECT 36.945 -0.085 37.115 0.085 ;
      RECT 36.485 -0.085 36.655 0.085 ;
      RECT 36.025 -0.085 36.195 0.085 ;
      RECT 35.565 -0.085 35.735 0.085 ;
      RECT 35.105 -0.085 35.275 0.085 ;
      RECT 34.645 -0.085 34.815 0.085 ;
      RECT 34.185 -0.085 34.355 0.085 ;
      RECT 33.725 -0.085 33.895 0.085 ;
      RECT 33.265 -0.085 33.435 0.085 ;
      RECT 32.805 -0.085 32.975 0.085 ;
      RECT 32.345 -0.085 32.515 0.085 ;
      RECT 31.885 -0.085 32.055 0.085 ;
      RECT 31.425 -0.085 31.595 0.085 ;
      RECT 30.965 -0.085 31.135 0.085 ;
      RECT 30.505 -0.085 30.675 0.085 ;
      RECT 30.045 -0.085 30.215 0.085 ;
      RECT 29.585 -0.085 29.755 0.085 ;
      RECT 29.125 -0.085 29.295 0.085 ;
      RECT 28.665 -0.085 28.835 0.085 ;
      RECT 28.205 -0.085 28.375 0.085 ;
      RECT 27.745 -0.085 27.915 0.085 ;
      RECT 27.285 -0.085 27.455 0.085 ;
      RECT 26.825 -0.085 26.995 0.085 ;
      RECT 26.365 -0.085 26.535 0.085 ;
      RECT 25.905 -0.085 26.075 0.085 ;
      RECT 25.445 -0.085 25.615 0.085 ;
      RECT 24.985 -0.085 25.155 0.085 ;
      RECT 24.525 -0.085 24.695 0.085 ;
      RECT 24.065 -0.085 24.235 0.085 ;
      RECT 23.605 -0.085 23.775 0.085 ;
      RECT 23.145 -0.085 23.315 0.085 ;
      RECT 22.685 -0.085 22.855 0.085 ;
      RECT 22.225 -0.085 22.395 0.085 ;
      RECT 21.765 -0.085 21.935 0.085 ;
      RECT 21.305 -0.085 21.475 0.085 ;
      RECT 20.845 -0.085 21.015 0.085 ;
      RECT 20.385 -0.085 20.555 0.085 ;
      RECT 19.925 -0.085 20.095 0.085 ;
      RECT 19.465 -0.085 19.635 0.085 ;
      RECT 19.005 -0.085 19.175 0.085 ;
      RECT 18.545 -0.085 18.715 0.085 ;
      RECT 18.085 -0.085 18.255 0.085 ;
      RECT 17.625 -0.085 17.795 0.085 ;
      RECT 17.165 -0.085 17.335 0.085 ;
      RECT 16.705 -0.085 16.875 0.085 ;
      RECT 16.245 -0.085 16.415 0.085 ;
      RECT 15.785 -0.085 15.955 0.085 ;
      RECT 15.325 -0.085 15.495 0.085 ;
      RECT 14.865 -0.085 15.035 0.085 ;
      RECT 14.405 -0.085 14.575 0.085 ;
      RECT 13.945 -0.085 14.115 0.085 ;
      RECT 13.485 -0.085 13.655 0.085 ;
      RECT 13.025 -0.085 13.195 0.085 ;
      RECT 12.565 -0.085 12.735 0.085 ;
      RECT 12.105 -0.085 12.275 0.085 ;
      RECT 11.645 -0.085 11.815 0.085 ;
      RECT 11.185 -0.085 11.355 0.085 ;
      RECT 10.725 -0.085 10.895 0.085 ;
      RECT 10.265 -0.085 10.435 0.085 ;
      RECT 9.805 -0.085 9.975 0.085 ;
      RECT 9.345 -0.085 9.515 0.085 ;
      RECT 8.885 -0.085 9.055 0.085 ;
      RECT 8.425 -0.085 8.595 0.085 ;
      RECT 7.965 -0.085 8.135 0.085 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.145 -0.085 0.315 0.085 ;
    LAYER via ;
      RECT 80.885 97.845 81.035 97.995 ;
      RECT 51.445 97.845 51.595 97.995 ;
      RECT 53.285 96.145 53.435 96.295 ;
      RECT 47.305 96.145 47.455 96.295 ;
      RECT 27.985 96.145 28.135 96.295 ;
      RECT 80.885 86.965 81.035 87.115 ;
      RECT 51.445 86.965 51.595 87.115 ;
      RECT 10.965 86.965 11.115 87.115 ;
      RECT 14.185 85.265 14.335 85.415 ;
      RECT 80.885 -0.075 81.035 0.075 ;
      RECT 51.445 -0.075 51.595 0.075 ;
      RECT 10.965 -0.075 11.115 0.075 ;
    LAYER via2 ;
      RECT 80.86 97.82 81.06 98.02 ;
      RECT 51.42 97.82 51.62 98.02 ;
      RECT 10.94 86.94 11.14 87.14 ;
      RECT 1.74 82.18 1.94 82.38 ;
      RECT 1.28 65.18 1.48 65.38 ;
      RECT 1.74 58.38 1.94 58.58 ;
      RECT 1.28 52.26 1.48 52.46 ;
      RECT 1.74 49.54 1.94 49.74 ;
      RECT 116.28 48.86 116.48 49.06 ;
      RECT 116.28 39.34 116.48 39.54 ;
      RECT 116.28 29.82 116.48 30.02 ;
      RECT 116.28 23.02 116.48 23.22 ;
      RECT 1.28 19.62 1.48 19.82 ;
      RECT 1.28 16.9 1.48 17.1 ;
      RECT 1.28 15.54 1.48 15.74 ;
      RECT 80.86 -0.1 81.06 0.1 ;
      RECT 51.42 -0.1 51.62 0.1 ;
      RECT 10.94 -0.1 11.14 0.1 ;
    LAYER via3 ;
      RECT 80.86 97.82 81.06 98.02 ;
      RECT 51.42 97.82 51.62 98.02 ;
      RECT 10.94 86.94 11.14 87.14 ;
      RECT 80.86 -0.1 81.06 0.1 ;
      RECT 51.42 -0.1 51.62 0.1 ;
      RECT 10.94 -0.1 11.14 0.1 ;
    LAYER OVERLAP ;
      POLYGON 0 0 0 87.04 25.76 87.04 25.76 97.92 92 97.92 92 87.04 117.76 87.04 117.76 0 ;
  END
END sb_1__0_

END LIBRARY
