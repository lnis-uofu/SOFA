VERSION 5.7 ;
BUSBITCHARS "[]" ;

UNITS
  DATABASE MICRONS 1000 ;
END UNITS

MANUFACTURINGGRID 0.005 ;

LAYER li1
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.46 ;
  WIDTH 0.17 ;
END li1

LAYER mcon
  TYPE CUT ;
END mcon

LAYER met1
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.34 ;
  WIDTH 0.14 ;
END met1

LAYER via
  TYPE CUT ;
END via

LAYER met2
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.46 ;
  WIDTH 0.14 ;
END met2

LAYER via2
  TYPE CUT ;
END via2

LAYER met3
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.68 ;
  WIDTH 0.3 ;
END met3

LAYER via3
  TYPE CUT ;
END via3

LAYER met4
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.92 ;
  WIDTH 0.3 ;
END met4

LAYER via4
  TYPE CUT ;
END via4

LAYER met5
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 3.4 ;
  WIDTH 1.6 ;
END met5

LAYER nwell
  TYPE MASTERSLICE ;
END nwell

LAYER pwell
  TYPE MASTERSLICE ;
END pwell

LAYER OVERLAP
  TYPE OVERLAP ;
END OVERLAP

VIA L1M1_PR
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.145 -0.115 0.145 0.115 ;
END L1M1_PR

VIA L1M1_PR_R
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.115 -0.145 0.115 0.145 ;
END L1M1_PR_R

VIA L1M1_PR_M
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.115 -0.145 0.115 0.145 ;
END L1M1_PR_M

VIA L1M1_PR_MR
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.145 -0.115 0.145 0.115 ;
END L1M1_PR_MR

VIA L1M1_PR_C
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.145 -0.145 0.145 0.145 ;
END L1M1_PR_C

VIA M1M2_PR
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR

VIA M1M2_PR_Enc
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_Enc

VIA M1M2_PR_R
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_R

VIA M1M2_PR_R_Enc
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR_R_Enc

VIA M1M2_PR_M
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_M

VIA M1M2_PR_M_Enc
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR_M_Enc

VIA M1M2_PR_MR
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR_MR

VIA M1M2_PR_MR_Enc
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_MR_Enc

VIA M1M2_PR_C
  LAYER met1 ;
    RECT -0.16 -0.16 0.16 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.16 0.16 0.16 ;
END M1M2_PR_C

VIA M2M3_PR
  LAYER met2 ;
    RECT -0.14 -0.185 0.14 0.185 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR

VIA M2M3_PR_R
  LAYER met2 ;
    RECT -0.185 -0.14 0.185 0.14 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_R

VIA M2M3_PR_M
  LAYER met2 ;
    RECT -0.14 -0.185 0.14 0.185 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_M

VIA M2M3_PR_MR
  LAYER met2 ;
    RECT -0.185 -0.14 0.185 0.14 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_MR

VIA M2M3_PR_C
  LAYER met2 ;
    RECT -0.185 -0.185 0.185 0.185 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_C

VIA M3M4_PR
  LAYER met3 ;
    RECT -0.19 -0.16 0.19 0.16 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR

VIA M3M4_PR_R
  LAYER met3 ;
    RECT -0.16 -0.19 0.16 0.19 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_R

VIA M3M4_PR_M
  LAYER met3 ;
    RECT -0.19 -0.16 0.19 0.16 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_M

VIA M3M4_PR_MR
  LAYER met3 ;
    RECT -0.16 -0.19 0.16 0.19 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_MR

VIA M3M4_PR_C
  LAYER met3 ;
    RECT -0.19 -0.19 0.19 0.19 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_C

VIA M4M5_PR
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR

VIA M4M5_PR_R
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_R

VIA M4M5_PR_M
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_M

VIA M4M5_PR_MR
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_MR

VIA M4M5_PR_C
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_C

SITE unit
  CLASS CORE ;
  SYMMETRY Y ;
  SIZE 0.46 BY 2.72 ;
END unit

SITE unithddbl
  CLASS CORE ;
  SIZE 0.46 BY 5.44 ;
END unithddbl

MACRO sb_0__2_
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  SIZE 84.64 BY 81.6 ;
  SYMMETRY X Y ;
  PIN prog_clk[0]
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER met2 ;
        RECT 14.19 0 14.33 1.36 ;
    END
  END prog_clk[0]
  PIN chanx_right_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 83.26 54.25 84.64 54.55 ;
    END
  END chanx_right_in[0]
  PIN chanx_right_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 83.26 42.01 84.64 42.31 ;
    END
  END chanx_right_in[1]
  PIN chanx_right_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 83.26 56.29 84.64 56.59 ;
    END
  END chanx_right_in[2]
  PIN chanx_right_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 83.26 26.37 84.64 26.67 ;
    END
  END chanx_right_in[3]
  PIN chanx_right_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 83.26 35.89 84.64 36.19 ;
    END
  END chanx_right_in[4]
  PIN chanx_right_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 83.26 69.21 84.64 69.51 ;
    END
  END chanx_right_in[5]
  PIN chanx_right_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 83.26 33.17 84.64 33.47 ;
    END
  END chanx_right_in[6]
  PIN chanx_right_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 83.26 63.77 84.64 64.07 ;
    END
  END chanx_right_in[7]
  PIN chanx_right_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 83.26 43.37 84.64 43.67 ;
    END
  END chanx_right_in[8]
  PIN chanx_right_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 83.26 76.01 84.64 76.31 ;
    END
  END chanx_right_in[9]
  PIN chanx_right_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.27 16.32 82.41 17.68 ;
    END
  END chanx_right_in[10]
  PIN chanx_right_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 83.26 77.37 84.64 77.67 ;
    END
  END chanx_right_in[11]
  PIN chanx_right_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 83.26 59.01 84.64 59.31 ;
    END
  END chanx_right_in[12]
  PIN chanx_right_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 83.26 22.97 84.64 23.27 ;
    END
  END chanx_right_in[13]
  PIN chanx_right_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.35 16.32 81.49 17.68 ;
    END
  END chanx_right_in[14]
  PIN chanx_right_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 83.26 67.85 84.64 68.15 ;
    END
  END chanx_right_in[15]
  PIN chanx_right_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 83.26 44.73 84.64 45.03 ;
    END
  END chanx_right_in[16]
  PIN chanx_right_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 83.26 21.61 84.64 21.91 ;
    END
  END chanx_right_in[17]
  PIN chanx_right_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 83.26 61.05 84.64 61.35 ;
    END
  END chanx_right_in[18]
  PIN chanx_right_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 83.26 65.13 84.64 65.43 ;
    END
  END chanx_right_in[19]
  PIN right_top_grid_pin_1_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 83.26 37.25 84.64 37.55 ;
    END
  END right_top_grid_pin_1_[0]
  PIN right_bottom_grid_pin_34_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 64.86 5.29 66.24 5.59 ;
    END
  END right_bottom_grid_pin_34_[0]
  PIN right_bottom_grid_pin_35_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 64.86 8.01 66.24 8.31 ;
    END
  END right_bottom_grid_pin_35_[0]
  PIN right_bottom_grid_pin_36_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 64.86 6.65 66.24 6.95 ;
    END
  END right_bottom_grid_pin_36_[0]
  PIN right_bottom_grid_pin_37_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.83 16.32 75.97 17.68 ;
    END
  END right_bottom_grid_pin_37_[0]
  PIN right_bottom_grid_pin_38_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.75 16.32 76.89 17.68 ;
    END
  END right_bottom_grid_pin_38_[0]
  PIN right_bottom_grid_pin_39_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.43 16.32 80.57 17.68 ;
    END
  END right_bottom_grid_pin_39_[0]
  PIN right_bottom_grid_pin_40_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.13 16.32 78.27 17.68 ;
    END
  END right_bottom_grid_pin_40_[0]
  PIN right_bottom_grid_pin_41_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.95 0 63.09 1.36 ;
    END
  END right_bottom_grid_pin_41_[0]
  PIN chany_bottom_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.91 0 52.05 1.36 ;
    END
  END chany_bottom_in[0]
  PIN chany_bottom_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.47 0 45.61 1.36 ;
    END
  END chany_bottom_in[1]
  PIN chany_bottom_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.83 0 52.97 1.36 ;
    END
  END chany_bottom_in[2]
  PIN chany_bottom_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.55 0 44.69 1.36 ;
    END
  END chany_bottom_in[3]
  PIN chany_bottom_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.71 0 42.85 1.36 ;
    END
  END chany_bottom_in[4]
  PIN chany_bottom_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.07 0 50.21 1.36 ;
    END
  END chany_bottom_in[5]
  PIN chany_bottom_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.17 0 20.31 1.36 ;
    END
  END chany_bottom_in[6]
  PIN chany_bottom_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.93 0 23.07 1.36 ;
    END
  END chany_bottom_in[7]
  PIN chany_bottom_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.21 0 8.35 1.36 ;
    END
  END chany_bottom_in[8]
  PIN chany_bottom_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.09 0 21.23 1.36 ;
    END
  END chany_bottom_in[9]
  PIN chany_bottom_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.51 0 33.65 1.36 ;
    END
  END chany_bottom_in[10]
  PIN chany_bottom_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.37 0 29.51 1.36 ;
    END
  END chany_bottom_in[11]
  PIN chany_bottom_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.99 0 51.13 1.36 ;
    END
  END chany_bottom_in[12]
  PIN chany_bottom_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.29 0 30.43 1.36 ;
    END
  END chany_bottom_in[13]
  PIN chany_bottom_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.45 0 28.59 1.36 ;
    END
  END chany_bottom_in[14]
  PIN chany_bottom_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.01 0 22.15 1.36 ;
    END
  END chany_bottom_in[15]
  PIN chany_bottom_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.27 0 36.41 1.36 ;
    END
  END chany_bottom_in[16]
  PIN chany_bottom_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.37 0 6.51 1.36 ;
    END
  END chany_bottom_in[17]
  PIN chany_bottom_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.21 0 31.35 1.36 ;
    END
  END chany_bottom_in[18]
  PIN chany_bottom_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.29 0 7.43 1.36 ;
    END
  END chany_bottom_in[19]
  PIN bottom_left_grid_pin_1_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.87 0 64.01 1.36 ;
    END
  END bottom_left_grid_pin_1_[0]
  PIN ccff_head[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 83.26 47.45 84.64 47.75 ;
    END
  END ccff_head[0]
  PIN chanx_right_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 83.26 52.89 84.64 53.19 ;
    END
  END chanx_right_out[0]
  PIN chanx_right_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 83.26 29.09 84.64 29.39 ;
    END
  END chanx_right_out[1]
  PIN chanx_right_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 83.26 50.17 84.64 50.47 ;
    END
  END chanx_right_out[2]
  PIN chanx_right_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 83.26 31.81 84.64 32.11 ;
    END
  END chanx_right_out[3]
  PIN chanx_right_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 83.26 70.57 84.64 70.87 ;
    END
  END chanx_right_out[4]
  PIN chanx_right_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 83.26 24.33 84.64 24.63 ;
    END
  END chanx_right_out[5]
  PIN chanx_right_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 83.26 66.49 84.64 66.79 ;
    END
  END chanx_right_out[6]
  PIN chanx_right_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 83.26 51.53 84.64 51.83 ;
    END
  END chanx_right_out[7]
  PIN chanx_right_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 83.26 34.53 84.64 34.83 ;
    END
  END chanx_right_out[8]
  PIN chanx_right_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 83.26 20.25 84.64 20.55 ;
    END
  END chanx_right_out[9]
  PIN chanx_right_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 83.26 71.93 84.64 72.23 ;
    END
  END chanx_right_out[10]
  PIN chanx_right_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 83.26 30.45 84.64 30.75 ;
    END
  END chanx_right_out[11]
  PIN chanx_right_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 83.26 39.29 84.64 39.59 ;
    END
  END chanx_right_out[12]
  PIN chanx_right_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 83.26 27.73 84.64 28.03 ;
    END
  END chanx_right_out[13]
  PIN chanx_right_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 83.26 48.81 84.64 49.11 ;
    END
  END chanx_right_out[14]
  PIN chanx_right_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 83.26 74.65 84.64 74.95 ;
    END
  END chanx_right_out[15]
  PIN chanx_right_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 83.26 57.65 84.64 57.95 ;
    END
  END chanx_right_out[16]
  PIN chanx_right_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 83.26 46.09 84.64 46.39 ;
    END
  END chanx_right_out[17]
  PIN chanx_right_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 83.26 73.29 84.64 73.59 ;
    END
  END chanx_right_out[18]
  PIN chanx_right_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 83.26 62.41 84.64 62.71 ;
    END
  END chanx_right_out[19]
  PIN chany_bottom_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.21 0 54.35 1.36 ;
    END
  END chany_bottom_out[0]
  PIN chany_bottom_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.23 0 48.37 1.36 ;
    END
  END chany_bottom_out[1]
  PIN chany_bottom_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.43 0 57.57 1.36 ;
    END
  END chany_bottom_out[2]
  PIN chany_bottom_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.53 0 27.67 1.36 ;
    END
  END chany_bottom_out[3]
  PIN chany_bottom_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.05 0 56.19 1.36 ;
    END
  END chany_bottom_out[4]
  PIN chany_bottom_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.85 0 23.99 1.36 ;
    END
  END chany_bottom_out[5]
  PIN chany_bottom_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.61 0 26.75 1.36 ;
    END
  END chany_bottom_out[6]
  PIN chany_bottom_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.39 0 46.53 1.36 ;
    END
  END chany_bottom_out[7]
  PIN chany_bottom_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.31 0 47.45 1.36 ;
    END
  END chany_bottom_out[8]
  PIN chany_bottom_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.77 0 24.91 1.36 ;
    END
  END chany_bottom_out[9]
  PIN chany_bottom_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.03 0 62.17 1.36 ;
    END
  END chany_bottom_out[10]
  PIN chany_bottom_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 44.93 0 45.23 1.36 ;
    END
  END chany_bottom_out[11]
  PIN chany_bottom_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.15 0 49.29 1.36 ;
    END
  END chany_bottom_out[12]
  PIN chany_bottom_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 9.05 0 9.35 1.36 ;
    END
  END chany_bottom_out[13]
  PIN chany_bottom_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 48.61 0 48.91 1.36 ;
    END
  END chany_bottom_out[14]
  PIN chany_bottom_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 46.77 0 47.07 1.36 ;
    END
  END chany_bottom_out[15]
  PIN chany_bottom_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.87 0 41.01 1.36 ;
    END
  END chany_bottom_out[16]
  PIN chany_bottom_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 5.37 0 5.67 1.36 ;
    END
  END chany_bottom_out[17]
  PIN chany_bottom_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 23.77 0 24.07 1.36 ;
    END
  END chany_bottom_out[18]
  PIN chany_bottom_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 7.21 0 7.51 1.36 ;
    END
  END chany_bottom_out[19]
  PIN ccff_tail[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.63 0 43.77 1.36 ;
    END
  END ccff_tail[0]
  PIN SC_IN_TOP
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 64.45 1.38 64.75 ;
    END
  END SC_IN_TOP
  PIN SC_IN_BOT
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.17 80.24 43.31 81.6 ;
    END
  END SC_IN_BOT
  PIN SC_OUT_TOP
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.25 80.24 42.39 81.6 ;
    END
  END SC_OUT_TOP
  PIN SC_OUT_BOT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 83.26 40.65 84.64 40.95 ;
    END
  END SC_OUT_BOT
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 0.48 2.96 ;
        RECT 65.76 2.48 66.24 2.96 ;
        RECT 0 7.92 0.48 8.4 ;
        RECT 65.76 7.92 66.24 8.4 ;
        RECT 0 13.36 0.48 13.84 ;
        RECT 65.76 13.36 66.24 13.84 ;
        RECT 0 18.8 0.48 19.28 ;
        RECT 84.16 18.8 84.64 19.28 ;
        RECT 0 24.24 0.48 24.72 ;
        RECT 84.16 24.24 84.64 24.72 ;
        RECT 0 29.68 0.48 30.16 ;
        RECT 84.16 29.68 84.64 30.16 ;
        RECT 0 35.12 0.48 35.6 ;
        RECT 84.16 35.12 84.64 35.6 ;
        RECT 0 40.56 0.48 41.04 ;
        RECT 84.16 40.56 84.64 41.04 ;
        RECT 0 46 0.48 46.48 ;
        RECT 84.16 46 84.64 46.48 ;
        RECT 0 51.44 0.48 51.92 ;
        RECT 84.16 51.44 84.64 51.92 ;
        RECT 0 56.88 0.48 57.36 ;
        RECT 84.16 56.88 84.64 57.36 ;
        RECT 0 62.32 0.48 62.8 ;
        RECT 84.16 62.32 84.64 62.8 ;
        RECT 0 67.76 0.48 68.24 ;
        RECT 84.16 67.76 84.64 68.24 ;
        RECT 0 73.2 0.48 73.68 ;
        RECT 84.16 73.2 84.64 73.68 ;
        RECT 0 78.64 0.48 79.12 ;
        RECT 84.16 78.64 84.64 79.12 ;
      LAYER met4 ;
        RECT 10.74 0 11.34 0.6 ;
        RECT 40.18 0 40.78 0.6 ;
        RECT 10.74 81 11.34 81.6 ;
        RECT 40.18 81 40.78 81.6 ;
      LAYER met5 ;
        RECT 0 26.96 3.2 30.16 ;
        RECT 81.44 26.96 84.64 30.16 ;
        RECT 0 67.76 3.2 70.96 ;
        RECT 81.44 67.76 84.64 70.96 ;
    END
  END VDD
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 0 66.24 0.24 ;
        RECT 0 5.2 0.48 5.68 ;
        RECT 65.76 5.2 66.24 5.68 ;
        RECT 0 10.64 0.48 11.12 ;
        RECT 65.76 10.64 66.24 11.12 ;
        RECT 0 16.08 84.64 16.56 ;
        RECT 0 21.52 0.48 22 ;
        RECT 84.16 21.52 84.64 22 ;
        RECT 0 26.96 0.48 27.44 ;
        RECT 84.16 26.96 84.64 27.44 ;
        RECT 0 32.4 0.48 32.88 ;
        RECT 84.16 32.4 84.64 32.88 ;
        RECT 0 37.84 0.48 38.32 ;
        RECT 84.16 37.84 84.64 38.32 ;
        RECT 0 43.28 0.48 43.76 ;
        RECT 84.16 43.28 84.64 43.76 ;
        RECT 0 48.72 0.48 49.2 ;
        RECT 84.16 48.72 84.64 49.2 ;
        RECT 0 54.16 0.48 54.64 ;
        RECT 84.16 54.16 84.64 54.64 ;
        RECT 0 59.6 0.48 60.08 ;
        RECT 84.16 59.6 84.64 60.08 ;
        RECT 0 65.04 0.48 65.52 ;
        RECT 84.16 65.04 84.64 65.52 ;
        RECT 0 70.48 0.48 70.96 ;
        RECT 84.16 70.48 84.64 70.96 ;
        RECT 0 75.92 0.48 76.4 ;
        RECT 84.16 75.92 84.64 76.4 ;
        RECT 0 81.36 84.64 81.6 ;
      LAYER met4 ;
        RECT 25.46 0 26.06 0.6 ;
        RECT 54.9 0 55.5 0.6 ;
        RECT 25.46 81 26.06 81.6 ;
        RECT 54.9 81 55.5 81.6 ;
      LAYER met5 ;
        RECT 0 47.36 3.2 50.56 ;
        RECT 81.44 47.36 84.64 50.56 ;
    END
  END VSS
  OBS
    LAYER li1 ;
      RECT 0 81.515 84.64 81.685 ;
      RECT 80.96 78.795 84.64 78.965 ;
      RECT 0 78.795 3.68 78.965 ;
      RECT 80.96 76.075 84.64 76.245 ;
      RECT 0 76.075 3.68 76.245 ;
      RECT 83.72 73.355 84.64 73.525 ;
      RECT 0 73.355 3.68 73.525 ;
      RECT 83.72 70.635 84.64 70.805 ;
      RECT 0 70.635 3.68 70.805 ;
      RECT 84.18 67.915 84.64 68.085 ;
      RECT 0 67.915 3.68 68.085 ;
      RECT 83.72 65.195 84.64 65.365 ;
      RECT 0 65.195 3.68 65.365 ;
      RECT 83.72 62.475 84.64 62.645 ;
      RECT 0 62.475 3.68 62.645 ;
      RECT 83.72 59.755 84.64 59.925 ;
      RECT 0 59.755 3.68 59.925 ;
      RECT 83.72 57.035 84.64 57.205 ;
      RECT 0 57.035 3.68 57.205 ;
      RECT 84.18 54.315 84.64 54.485 ;
      RECT 0 54.315 3.68 54.485 ;
      RECT 84.18 51.595 84.64 51.765 ;
      RECT 0 51.595 3.68 51.765 ;
      RECT 83.72 48.875 84.64 49.045 ;
      RECT 0 48.875 3.68 49.045 ;
      RECT 83.72 46.155 84.64 46.325 ;
      RECT 0 46.155 3.68 46.325 ;
      RECT 83.72 43.435 84.64 43.605 ;
      RECT 0 43.435 3.68 43.605 ;
      RECT 83.72 40.715 84.64 40.885 ;
      RECT 0 40.715 3.68 40.885 ;
      RECT 83.72 37.995 84.64 38.165 ;
      RECT 0 37.995 3.68 38.165 ;
      RECT 83.72 35.275 84.64 35.445 ;
      RECT 0 35.275 3.68 35.445 ;
      RECT 83.72 32.555 84.64 32.725 ;
      RECT 0 32.555 3.68 32.725 ;
      RECT 83.72 29.835 84.64 30.005 ;
      RECT 0 29.835 3.68 30.005 ;
      RECT 80.96 27.115 84.64 27.285 ;
      RECT 0 27.115 3.68 27.285 ;
      RECT 80.96 24.395 84.64 24.565 ;
      RECT 0 24.395 3.68 24.565 ;
      RECT 83.72 21.675 84.64 21.845 ;
      RECT 0 21.675 3.68 21.845 ;
      RECT 83.72 18.955 84.64 19.125 ;
      RECT 0 18.955 3.68 19.125 ;
      RECT 65.32 16.235 84.64 16.405 ;
      RECT 0 16.235 3.68 16.405 ;
      RECT 65.32 13.515 66.24 13.685 ;
      RECT 0 13.515 3.68 13.685 ;
      RECT 62.56 10.795 66.24 10.965 ;
      RECT 0 10.795 3.68 10.965 ;
      RECT 62.56 8.075 66.24 8.245 ;
      RECT 0 8.075 3.68 8.245 ;
      RECT 65.32 5.355 66.24 5.525 ;
      RECT 0 5.355 3.68 5.525 ;
      RECT 65.32 2.635 66.24 2.805 ;
      RECT 0 2.635 3.68 2.805 ;
      RECT 0 -0.085 66.24 0.085 ;
    LAYER met2 ;
      RECT 55.06 81.415 55.34 81.785 ;
      RECT 25.62 81.415 25.9 81.785 ;
      POLYGON 66.31 27.27 66.31 16.59 64.79 16.59 64.79 16.73 66.17 16.73 66.17 27.27 ;
      RECT 80.83 17.86 81.09 18.18 ;
      RECT 32.99 1.54 33.25 1.86 ;
      RECT 27.01 1.54 27.27 1.86 ;
      RECT 55.06 -0.185 55.34 0.185 ;
      RECT 25.62 -0.185 25.9 0.185 ;
      POLYGON 84.36 81.32 84.36 16.6 82.69 16.6 82.69 17.96 81.99 17.96 81.99 16.6 81.77 16.6 81.77 17.96 81.07 17.96 81.07 16.6 80.85 16.6 80.85 17.96 80.15 17.96 80.15 16.6 78.55 16.6 78.55 17.96 77.85 17.96 77.85 16.6 77.17 16.6 77.17 17.96 76.47 17.96 76.47 16.6 76.25 16.6 76.25 17.96 75.55 17.96 75.55 16.6 65.96 16.6 65.96 0.28 64.29 0.28 64.29 1.64 63.59 1.64 63.59 0.28 63.37 0.28 63.37 1.64 62.67 1.64 62.67 0.28 62.45 0.28 62.45 1.64 61.75 1.64 61.75 0.28 57.85 0.28 57.85 1.64 57.15 1.64 57.15 0.28 56.47 0.28 56.47 1.64 55.77 1.64 55.77 0.28 54.63 0.28 54.63 1.64 53.93 1.64 53.93 0.28 53.25 0.28 53.25 1.64 52.55 1.64 52.55 0.28 52.33 0.28 52.33 1.64 51.63 1.64 51.63 0.28 51.41 0.28 51.41 1.64 50.71 1.64 50.71 0.28 50.49 0.28 50.49 1.64 49.79 1.64 49.79 0.28 49.57 0.28 49.57 1.64 48.87 1.64 48.87 0.28 48.65 0.28 48.65 1.64 47.95 1.64 47.95 0.28 47.73 0.28 47.73 1.64 47.03 1.64 47.03 0.28 46.81 0.28 46.81 1.64 46.11 1.64 46.11 0.28 45.89 0.28 45.89 1.64 45.19 1.64 45.19 0.28 44.97 0.28 44.97 1.64 44.27 1.64 44.27 0.28 44.05 0.28 44.05 1.64 43.35 1.64 43.35 0.28 43.13 0.28 43.13 1.64 42.43 1.64 42.43 0.28 41.29 0.28 41.29 1.64 40.59 1.64 40.59 0.28 36.69 0.28 36.69 1.64 35.99 1.64 35.99 0.28 33.93 0.28 33.93 1.64 33.23 1.64 33.23 0.28 31.63 0.28 31.63 1.64 30.93 1.64 30.93 0.28 30.71 0.28 30.71 1.64 30.01 1.64 30.01 0.28 29.79 0.28 29.79 1.64 29.09 1.64 29.09 0.28 28.87 0.28 28.87 1.64 28.17 1.64 28.17 0.28 27.95 0.28 27.95 1.64 27.25 1.64 27.25 0.28 27.03 0.28 27.03 1.64 26.33 1.64 26.33 0.28 25.19 0.28 25.19 1.64 24.49 1.64 24.49 0.28 24.27 0.28 24.27 1.64 23.57 1.64 23.57 0.28 23.35 0.28 23.35 1.64 22.65 1.64 22.65 0.28 22.43 0.28 22.43 1.64 21.73 1.64 21.73 0.28 21.51 0.28 21.51 1.64 20.81 1.64 20.81 0.28 20.59 0.28 20.59 1.64 19.89 1.64 19.89 0.28 14.61 0.28 14.61 1.64 13.91 1.64 13.91 0.28 8.63 0.28 8.63 1.64 7.93 1.64 7.93 0.28 7.71 0.28 7.71 1.64 7.01 1.64 7.01 0.28 6.79 0.28 6.79 1.64 6.09 1.64 6.09 0.28 0.28 0.28 0.28 81.32 41.97 81.32 41.97 79.96 42.67 79.96 42.67 81.32 42.89 81.32 42.89 79.96 43.59 79.96 43.59 81.32 ;
    LAYER met3 ;
      POLYGON 55.365 81.765 55.365 81.76 55.58 81.76 55.58 81.44 55.365 81.44 55.365 81.435 55.035 81.435 55.035 81.44 54.82 81.44 54.82 81.76 55.035 81.76 55.035 81.765 ;
      POLYGON 25.925 81.765 25.925 81.76 26.14 81.76 26.14 81.44 25.925 81.44 25.925 81.435 25.595 81.435 25.595 81.44 25.38 81.44 25.38 81.76 25.595 81.76 25.595 81.765 ;
      POLYGON 83.425 38.245 83.425 37.915 83.095 37.915 83.095 37.93 72.07 37.93 72.07 38.23 83.095 38.23 83.095 38.245 ;
      POLYGON 83.41 23.95 83.41 23.67 82.86 23.67 82.86 23.65 30.21 23.65 30.21 23.95 ;
      POLYGON 64.565 9.005 64.565 8.675 64.235 8.675 64.235 8.69 57.35 8.69 57.35 8.99 64.235 8.99 64.235 9.005 ;
      POLYGON 55.365 0.165 55.365 0.16 55.58 0.16 55.58 -0.16 55.365 -0.16 55.365 -0.165 55.035 -0.165 55.035 -0.16 54.82 -0.16 54.82 0.16 55.035 0.16 55.035 0.165 ;
      POLYGON 25.925 0.165 25.925 0.16 26.14 0.16 26.14 -0.16 25.925 -0.16 25.925 -0.165 25.595 -0.165 25.595 -0.16 25.38 -0.16 25.38 0.16 25.595 0.16 25.595 0.165 ;
      POLYGON 84.24 81.2 84.24 78.07 82.86 78.07 82.86 76.97 84.24 76.97 84.24 76.71 82.86 76.71 82.86 75.61 84.24 75.61 84.24 75.35 82.86 75.35 82.86 74.25 84.24 74.25 84.24 73.99 82.86 73.99 82.86 72.89 84.24 72.89 84.24 72.63 82.86 72.63 82.86 71.53 84.24 71.53 84.24 71.27 82.86 71.27 82.86 70.17 84.24 70.17 84.24 69.91 82.86 69.91 82.86 68.81 84.24 68.81 84.24 68.55 82.86 68.55 82.86 67.45 84.24 67.45 84.24 67.19 82.86 67.19 82.86 66.09 84.24 66.09 84.24 65.83 82.86 65.83 82.86 64.73 84.24 64.73 84.24 64.47 82.86 64.47 82.86 63.37 84.24 63.37 84.24 63.11 82.86 63.11 82.86 62.01 84.24 62.01 84.24 61.75 82.86 61.75 82.86 60.65 84.24 60.65 84.24 59.71 82.86 59.71 82.86 58.61 84.24 58.61 84.24 58.35 82.86 58.35 82.86 57.25 84.24 57.25 84.24 56.99 82.86 56.99 82.86 55.89 84.24 55.89 84.24 54.95 82.86 54.95 82.86 53.85 84.24 53.85 84.24 53.59 82.86 53.59 82.86 52.49 84.24 52.49 84.24 52.23 82.86 52.23 82.86 51.13 84.24 51.13 84.24 50.87 82.86 50.87 82.86 49.77 84.24 49.77 84.24 49.51 82.86 49.51 82.86 48.41 84.24 48.41 84.24 48.15 82.86 48.15 82.86 47.05 84.24 47.05 84.24 46.79 82.86 46.79 82.86 45.69 84.24 45.69 84.24 45.43 82.86 45.43 82.86 44.33 84.24 44.33 84.24 44.07 82.86 44.07 82.86 42.97 84.24 42.97 84.24 42.71 82.86 42.71 82.86 41.61 84.24 41.61 84.24 41.35 82.86 41.35 82.86 40.25 84.24 40.25 84.24 39.99 82.86 39.99 82.86 38.89 84.24 38.89 84.24 37.95 82.86 37.95 82.86 36.85 84.24 36.85 84.24 36.59 82.86 36.59 82.86 35.49 84.24 35.49 84.24 35.23 82.86 35.23 82.86 34.13 84.24 34.13 84.24 33.87 82.86 33.87 82.86 32.77 84.24 32.77 84.24 32.51 82.86 32.51 82.86 31.41 84.24 31.41 84.24 31.15 82.86 31.15 82.86 30.05 84.24 30.05 84.24 29.79 82.86 29.79 82.86 28.69 84.24 28.69 84.24 28.43 82.86 28.43 82.86 27.33 84.24 27.33 84.24 27.07 82.86 27.07 82.86 25.97 84.24 25.97 84.24 25.03 82.86 25.03 82.86 23.93 84.24 23.93 84.24 23.67 82.86 23.67 82.86 22.57 84.24 22.57 84.24 22.31 82.86 22.31 82.86 21.21 84.24 21.21 84.24 20.95 82.86 20.95 82.86 19.85 84.24 19.85 84.24 16.72 65.84 16.72 65.84 8.71 64.46 8.71 64.46 7.61 65.84 7.61 65.84 7.35 64.46 7.35 64.46 6.25 65.84 6.25 65.84 5.99 64.46 5.99 64.46 4.89 65.84 4.89 65.84 0.4 0.4 0.4 0.4 64.05 1.78 64.05 1.78 65.15 0.4 65.15 0.4 81.2 ;
    LAYER met4 ;
      POLYGON 84.24 81.2 84.24 16.72 65.84 16.72 65.84 0.4 55.9 0.4 55.9 1 54.5 1 54.5 0.4 49.31 0.4 49.31 1.76 48.21 1.76 48.21 0.4 47.47 0.4 47.47 1.76 46.37 1.76 46.37 0.4 45.63 0.4 45.63 1.76 44.53 1.76 44.53 0.4 41.18 0.4 41.18 1 39.78 1 39.78 0.4 26.46 0.4 26.46 1 25.06 1 25.06 0.4 24.47 0.4 24.47 1.76 23.37 1.76 23.37 0.4 11.74 0.4 11.74 1 10.34 1 10.34 0.4 9.75 0.4 9.75 1.76 8.65 1.76 8.65 0.4 7.91 0.4 7.91 1.76 6.81 1.76 6.81 0.4 6.07 0.4 6.07 1.76 4.97 1.76 4.97 0.4 0.4 0.4 0.4 81.2 10.34 81.2 10.34 80.6 11.74 80.6 11.74 81.2 25.06 81.2 25.06 80.6 26.46 80.6 26.46 81.2 39.78 81.2 39.78 80.6 41.18 80.6 41.18 81.2 54.5 81.2 54.5 80.6 55.9 80.6 55.9 81.2 ;
    LAYER met5 ;
      POLYGON 83.04 80 83.04 72.56 79.84 72.56 79.84 66.16 83.04 66.16 83.04 52.16 79.84 52.16 79.84 45.76 83.04 45.76 83.04 31.76 79.84 31.76 79.84 25.36 83.04 25.36 83.04 17.92 64.64 17.92 64.64 1.6 1.6 1.6 1.6 25.36 4.8 25.36 4.8 31.76 1.6 31.76 1.6 45.76 4.8 45.76 4.8 52.16 1.6 52.16 1.6 66.16 4.8 66.16 4.8 72.56 1.6 72.56 1.6 80 ;
    LAYER met1 ;
      POLYGON 84.36 81.08 84.36 79.4 83.88 79.4 83.88 78.36 84.36 78.36 84.36 76.68 83.88 76.68 83.88 75.64 84.36 75.64 84.36 73.96 83.88 73.96 83.88 72.92 84.36 72.92 84.36 71.24 83.88 71.24 83.88 70.2 84.36 70.2 84.36 68.52 83.88 68.52 83.88 67.48 84.36 67.48 84.36 65.8 83.88 65.8 83.88 64.76 84.36 64.76 84.36 63.08 83.88 63.08 83.88 62.04 84.36 62.04 84.36 60.36 83.88 60.36 83.88 59.32 84.36 59.32 84.36 57.64 83.88 57.64 83.88 56.6 84.36 56.6 84.36 54.92 83.88 54.92 83.88 53.88 84.36 53.88 84.36 52.2 83.88 52.2 83.88 51.16 84.36 51.16 84.36 49.48 83.88 49.48 83.88 48.44 84.36 48.44 84.36 46.76 83.88 46.76 83.88 45.72 84.36 45.72 84.36 44.04 83.88 44.04 83.88 43 84.36 43 84.36 41.32 83.88 41.32 83.88 40.28 84.36 40.28 84.36 38.6 83.88 38.6 83.88 37.56 84.36 37.56 84.36 35.88 83.88 35.88 83.88 34.84 84.36 34.84 84.36 33.16 83.88 33.16 83.88 32.12 84.36 32.12 84.36 30.44 83.88 30.44 83.88 29.4 84.36 29.4 84.36 27.72 83.88 27.72 83.88 26.68 84.36 26.68 84.36 25 83.88 25 83.88 23.96 84.36 23.96 84.36 22.28 83.88 22.28 83.88 21.24 84.36 21.24 84.36 19.56 83.88 19.56 83.88 18.52 84.36 18.52 84.36 16.84 0.28 16.84 0.28 18.52 0.76 18.52 0.76 19.56 0.28 19.56 0.28 21.24 0.76 21.24 0.76 22.28 0.28 22.28 0.28 23.96 0.76 23.96 0.76 25 0.28 25 0.28 26.68 0.76 26.68 0.76 27.72 0.28 27.72 0.28 29.4 0.76 29.4 0.76 30.44 0.28 30.44 0.28 32.12 0.76 32.12 0.76 33.16 0.28 33.16 0.28 34.84 0.76 34.84 0.76 35.88 0.28 35.88 0.28 37.56 0.76 37.56 0.76 38.6 0.28 38.6 0.28 40.28 0.76 40.28 0.76 41.32 0.28 41.32 0.28 43 0.76 43 0.76 44.04 0.28 44.04 0.28 45.72 0.76 45.72 0.76 46.76 0.28 46.76 0.28 48.44 0.76 48.44 0.76 49.48 0.28 49.48 0.28 51.16 0.76 51.16 0.76 52.2 0.28 52.2 0.28 53.88 0.76 53.88 0.76 54.92 0.28 54.92 0.28 56.6 0.76 56.6 0.76 57.64 0.28 57.64 0.28 59.32 0.76 59.32 0.76 60.36 0.28 60.36 0.28 62.04 0.76 62.04 0.76 63.08 0.28 63.08 0.28 64.76 0.76 64.76 0.76 65.8 0.28 65.8 0.28 67.48 0.76 67.48 0.76 68.52 0.28 68.52 0.28 70.2 0.76 70.2 0.76 71.24 0.28 71.24 0.28 72.92 0.76 72.92 0.76 73.96 0.28 73.96 0.28 75.64 0.76 75.64 0.76 76.68 0.28 76.68 0.28 78.36 0.76 78.36 0.76 79.4 0.28 79.4 0.28 81.08 ;
      POLYGON 65.96 15.8 65.96 14.12 65.48 14.12 65.48 13.08 65.96 13.08 65.96 11.4 65.48 11.4 65.48 10.36 65.96 10.36 65.96 8.68 65.48 8.68 65.48 7.64 65.96 7.64 65.96 5.96 65.48 5.96 65.48 4.92 65.96 4.92 65.96 3.24 65.48 3.24 65.48 2.2 65.96 2.2 65.96 0.52 0.28 0.52 0.28 2.2 0.76 2.2 0.76 3.24 0.28 3.24 0.28 4.92 0.76 4.92 0.76 5.96 0.28 5.96 0.28 7.64 0.76 7.64 0.76 8.68 0.28 8.68 0.28 10.36 0.76 10.36 0.76 11.4 0.28 11.4 0.28 13.08 0.76 13.08 0.76 14.12 0.28 14.12 0.28 15.8 ;
    LAYER li1 ;
      POLYGON 84.47 81.43 84.47 16.49 66.07 16.49 66.07 0.17 0.17 0.17 0.17 81.43 ;
    LAYER mcon ;
      RECT 84.325 81.515 84.495 81.685 ;
      RECT 83.865 81.515 84.035 81.685 ;
      RECT 83.405 81.515 83.575 81.685 ;
      RECT 82.945 81.515 83.115 81.685 ;
      RECT 82.485 81.515 82.655 81.685 ;
      RECT 82.025 81.515 82.195 81.685 ;
      RECT 81.565 81.515 81.735 81.685 ;
      RECT 81.105 81.515 81.275 81.685 ;
      RECT 80.645 81.515 80.815 81.685 ;
      RECT 80.185 81.515 80.355 81.685 ;
      RECT 79.725 81.515 79.895 81.685 ;
      RECT 79.265 81.515 79.435 81.685 ;
      RECT 78.805 81.515 78.975 81.685 ;
      RECT 78.345 81.515 78.515 81.685 ;
      RECT 77.885 81.515 78.055 81.685 ;
      RECT 77.425 81.515 77.595 81.685 ;
      RECT 76.965 81.515 77.135 81.685 ;
      RECT 76.505 81.515 76.675 81.685 ;
      RECT 76.045 81.515 76.215 81.685 ;
      RECT 75.585 81.515 75.755 81.685 ;
      RECT 75.125 81.515 75.295 81.685 ;
      RECT 74.665 81.515 74.835 81.685 ;
      RECT 74.205 81.515 74.375 81.685 ;
      RECT 73.745 81.515 73.915 81.685 ;
      RECT 73.285 81.515 73.455 81.685 ;
      RECT 72.825 81.515 72.995 81.685 ;
      RECT 72.365 81.515 72.535 81.685 ;
      RECT 71.905 81.515 72.075 81.685 ;
      RECT 71.445 81.515 71.615 81.685 ;
      RECT 70.985 81.515 71.155 81.685 ;
      RECT 70.525 81.515 70.695 81.685 ;
      RECT 70.065 81.515 70.235 81.685 ;
      RECT 69.605 81.515 69.775 81.685 ;
      RECT 69.145 81.515 69.315 81.685 ;
      RECT 68.685 81.515 68.855 81.685 ;
      RECT 68.225 81.515 68.395 81.685 ;
      RECT 67.765 81.515 67.935 81.685 ;
      RECT 67.305 81.515 67.475 81.685 ;
      RECT 66.845 81.515 67.015 81.685 ;
      RECT 66.385 81.515 66.555 81.685 ;
      RECT 65.925 81.515 66.095 81.685 ;
      RECT 65.465 81.515 65.635 81.685 ;
      RECT 65.005 81.515 65.175 81.685 ;
      RECT 64.545 81.515 64.715 81.685 ;
      RECT 64.085 81.515 64.255 81.685 ;
      RECT 63.625 81.515 63.795 81.685 ;
      RECT 63.165 81.515 63.335 81.685 ;
      RECT 62.705 81.515 62.875 81.685 ;
      RECT 62.245 81.515 62.415 81.685 ;
      RECT 61.785 81.515 61.955 81.685 ;
      RECT 61.325 81.515 61.495 81.685 ;
      RECT 60.865 81.515 61.035 81.685 ;
      RECT 60.405 81.515 60.575 81.685 ;
      RECT 59.945 81.515 60.115 81.685 ;
      RECT 59.485 81.515 59.655 81.685 ;
      RECT 59.025 81.515 59.195 81.685 ;
      RECT 58.565 81.515 58.735 81.685 ;
      RECT 58.105 81.515 58.275 81.685 ;
      RECT 57.645 81.515 57.815 81.685 ;
      RECT 57.185 81.515 57.355 81.685 ;
      RECT 56.725 81.515 56.895 81.685 ;
      RECT 56.265 81.515 56.435 81.685 ;
      RECT 55.805 81.515 55.975 81.685 ;
      RECT 55.345 81.515 55.515 81.685 ;
      RECT 54.885 81.515 55.055 81.685 ;
      RECT 54.425 81.515 54.595 81.685 ;
      RECT 53.965 81.515 54.135 81.685 ;
      RECT 53.505 81.515 53.675 81.685 ;
      RECT 53.045 81.515 53.215 81.685 ;
      RECT 52.585 81.515 52.755 81.685 ;
      RECT 52.125 81.515 52.295 81.685 ;
      RECT 51.665 81.515 51.835 81.685 ;
      RECT 51.205 81.515 51.375 81.685 ;
      RECT 50.745 81.515 50.915 81.685 ;
      RECT 50.285 81.515 50.455 81.685 ;
      RECT 49.825 81.515 49.995 81.685 ;
      RECT 49.365 81.515 49.535 81.685 ;
      RECT 48.905 81.515 49.075 81.685 ;
      RECT 48.445 81.515 48.615 81.685 ;
      RECT 47.985 81.515 48.155 81.685 ;
      RECT 47.525 81.515 47.695 81.685 ;
      RECT 47.065 81.515 47.235 81.685 ;
      RECT 46.605 81.515 46.775 81.685 ;
      RECT 46.145 81.515 46.315 81.685 ;
      RECT 45.685 81.515 45.855 81.685 ;
      RECT 45.225 81.515 45.395 81.685 ;
      RECT 44.765 81.515 44.935 81.685 ;
      RECT 44.305 81.515 44.475 81.685 ;
      RECT 43.845 81.515 44.015 81.685 ;
      RECT 43.385 81.515 43.555 81.685 ;
      RECT 42.925 81.515 43.095 81.685 ;
      RECT 42.465 81.515 42.635 81.685 ;
      RECT 42.005 81.515 42.175 81.685 ;
      RECT 41.545 81.515 41.715 81.685 ;
      RECT 41.085 81.515 41.255 81.685 ;
      RECT 40.625 81.515 40.795 81.685 ;
      RECT 40.165 81.515 40.335 81.685 ;
      RECT 39.705 81.515 39.875 81.685 ;
      RECT 39.245 81.515 39.415 81.685 ;
      RECT 38.785 81.515 38.955 81.685 ;
      RECT 38.325 81.515 38.495 81.685 ;
      RECT 37.865 81.515 38.035 81.685 ;
      RECT 37.405 81.515 37.575 81.685 ;
      RECT 36.945 81.515 37.115 81.685 ;
      RECT 36.485 81.515 36.655 81.685 ;
      RECT 36.025 81.515 36.195 81.685 ;
      RECT 35.565 81.515 35.735 81.685 ;
      RECT 35.105 81.515 35.275 81.685 ;
      RECT 34.645 81.515 34.815 81.685 ;
      RECT 34.185 81.515 34.355 81.685 ;
      RECT 33.725 81.515 33.895 81.685 ;
      RECT 33.265 81.515 33.435 81.685 ;
      RECT 32.805 81.515 32.975 81.685 ;
      RECT 32.345 81.515 32.515 81.685 ;
      RECT 31.885 81.515 32.055 81.685 ;
      RECT 31.425 81.515 31.595 81.685 ;
      RECT 30.965 81.515 31.135 81.685 ;
      RECT 30.505 81.515 30.675 81.685 ;
      RECT 30.045 81.515 30.215 81.685 ;
      RECT 29.585 81.515 29.755 81.685 ;
      RECT 29.125 81.515 29.295 81.685 ;
      RECT 28.665 81.515 28.835 81.685 ;
      RECT 28.205 81.515 28.375 81.685 ;
      RECT 27.745 81.515 27.915 81.685 ;
      RECT 27.285 81.515 27.455 81.685 ;
      RECT 26.825 81.515 26.995 81.685 ;
      RECT 26.365 81.515 26.535 81.685 ;
      RECT 25.905 81.515 26.075 81.685 ;
      RECT 25.445 81.515 25.615 81.685 ;
      RECT 24.985 81.515 25.155 81.685 ;
      RECT 24.525 81.515 24.695 81.685 ;
      RECT 24.065 81.515 24.235 81.685 ;
      RECT 23.605 81.515 23.775 81.685 ;
      RECT 23.145 81.515 23.315 81.685 ;
      RECT 22.685 81.515 22.855 81.685 ;
      RECT 22.225 81.515 22.395 81.685 ;
      RECT 21.765 81.515 21.935 81.685 ;
      RECT 21.305 81.515 21.475 81.685 ;
      RECT 20.845 81.515 21.015 81.685 ;
      RECT 20.385 81.515 20.555 81.685 ;
      RECT 19.925 81.515 20.095 81.685 ;
      RECT 19.465 81.515 19.635 81.685 ;
      RECT 19.005 81.515 19.175 81.685 ;
      RECT 18.545 81.515 18.715 81.685 ;
      RECT 18.085 81.515 18.255 81.685 ;
      RECT 17.625 81.515 17.795 81.685 ;
      RECT 17.165 81.515 17.335 81.685 ;
      RECT 16.705 81.515 16.875 81.685 ;
      RECT 16.245 81.515 16.415 81.685 ;
      RECT 15.785 81.515 15.955 81.685 ;
      RECT 15.325 81.515 15.495 81.685 ;
      RECT 14.865 81.515 15.035 81.685 ;
      RECT 14.405 81.515 14.575 81.685 ;
      RECT 13.945 81.515 14.115 81.685 ;
      RECT 13.485 81.515 13.655 81.685 ;
      RECT 13.025 81.515 13.195 81.685 ;
      RECT 12.565 81.515 12.735 81.685 ;
      RECT 12.105 81.515 12.275 81.685 ;
      RECT 11.645 81.515 11.815 81.685 ;
      RECT 11.185 81.515 11.355 81.685 ;
      RECT 10.725 81.515 10.895 81.685 ;
      RECT 10.265 81.515 10.435 81.685 ;
      RECT 9.805 81.515 9.975 81.685 ;
      RECT 9.345 81.515 9.515 81.685 ;
      RECT 8.885 81.515 9.055 81.685 ;
      RECT 8.425 81.515 8.595 81.685 ;
      RECT 7.965 81.515 8.135 81.685 ;
      RECT 7.505 81.515 7.675 81.685 ;
      RECT 7.045 81.515 7.215 81.685 ;
      RECT 6.585 81.515 6.755 81.685 ;
      RECT 6.125 81.515 6.295 81.685 ;
      RECT 5.665 81.515 5.835 81.685 ;
      RECT 5.205 81.515 5.375 81.685 ;
      RECT 4.745 81.515 4.915 81.685 ;
      RECT 4.285 81.515 4.455 81.685 ;
      RECT 3.825 81.515 3.995 81.685 ;
      RECT 3.365 81.515 3.535 81.685 ;
      RECT 2.905 81.515 3.075 81.685 ;
      RECT 2.445 81.515 2.615 81.685 ;
      RECT 1.985 81.515 2.155 81.685 ;
      RECT 1.525 81.515 1.695 81.685 ;
      RECT 1.065 81.515 1.235 81.685 ;
      RECT 0.605 81.515 0.775 81.685 ;
      RECT 0.145 81.515 0.315 81.685 ;
      RECT 84.325 78.795 84.495 78.965 ;
      RECT 83.865 78.795 84.035 78.965 ;
      RECT 0.605 78.795 0.775 78.965 ;
      RECT 0.145 78.795 0.315 78.965 ;
      RECT 84.325 76.075 84.495 76.245 ;
      RECT 83.865 76.075 84.035 76.245 ;
      RECT 0.605 76.075 0.775 76.245 ;
      RECT 0.145 76.075 0.315 76.245 ;
      RECT 84.325 73.355 84.495 73.525 ;
      RECT 83.865 73.355 84.035 73.525 ;
      RECT 0.605 73.355 0.775 73.525 ;
      RECT 0.145 73.355 0.315 73.525 ;
      RECT 84.325 70.635 84.495 70.805 ;
      RECT 83.865 70.635 84.035 70.805 ;
      RECT 0.605 70.635 0.775 70.805 ;
      RECT 0.145 70.635 0.315 70.805 ;
      RECT 84.325 67.915 84.495 68.085 ;
      RECT 83.865 67.915 84.035 68.085 ;
      RECT 0.605 67.915 0.775 68.085 ;
      RECT 0.145 67.915 0.315 68.085 ;
      RECT 84.325 65.195 84.495 65.365 ;
      RECT 83.865 65.195 84.035 65.365 ;
      RECT 0.605 65.195 0.775 65.365 ;
      RECT 0.145 65.195 0.315 65.365 ;
      RECT 84.325 62.475 84.495 62.645 ;
      RECT 83.865 62.475 84.035 62.645 ;
      RECT 0.605 62.475 0.775 62.645 ;
      RECT 0.145 62.475 0.315 62.645 ;
      RECT 84.325 59.755 84.495 59.925 ;
      RECT 83.865 59.755 84.035 59.925 ;
      RECT 0.605 59.755 0.775 59.925 ;
      RECT 0.145 59.755 0.315 59.925 ;
      RECT 84.325 57.035 84.495 57.205 ;
      RECT 83.865 57.035 84.035 57.205 ;
      RECT 0.605 57.035 0.775 57.205 ;
      RECT 0.145 57.035 0.315 57.205 ;
      RECT 84.325 54.315 84.495 54.485 ;
      RECT 83.865 54.315 84.035 54.485 ;
      RECT 0.605 54.315 0.775 54.485 ;
      RECT 0.145 54.315 0.315 54.485 ;
      RECT 84.325 51.595 84.495 51.765 ;
      RECT 83.865 51.595 84.035 51.765 ;
      RECT 0.605 51.595 0.775 51.765 ;
      RECT 0.145 51.595 0.315 51.765 ;
      RECT 84.325 48.875 84.495 49.045 ;
      RECT 83.865 48.875 84.035 49.045 ;
      RECT 0.605 48.875 0.775 49.045 ;
      RECT 0.145 48.875 0.315 49.045 ;
      RECT 84.325 46.155 84.495 46.325 ;
      RECT 83.865 46.155 84.035 46.325 ;
      RECT 0.605 46.155 0.775 46.325 ;
      RECT 0.145 46.155 0.315 46.325 ;
      RECT 84.325 43.435 84.495 43.605 ;
      RECT 83.865 43.435 84.035 43.605 ;
      RECT 0.605 43.435 0.775 43.605 ;
      RECT 0.145 43.435 0.315 43.605 ;
      RECT 84.325 40.715 84.495 40.885 ;
      RECT 83.865 40.715 84.035 40.885 ;
      RECT 0.605 40.715 0.775 40.885 ;
      RECT 0.145 40.715 0.315 40.885 ;
      RECT 84.325 37.995 84.495 38.165 ;
      RECT 83.865 37.995 84.035 38.165 ;
      RECT 0.605 37.995 0.775 38.165 ;
      RECT 0.145 37.995 0.315 38.165 ;
      RECT 84.325 35.275 84.495 35.445 ;
      RECT 83.865 35.275 84.035 35.445 ;
      RECT 0.605 35.275 0.775 35.445 ;
      RECT 0.145 35.275 0.315 35.445 ;
      RECT 84.325 32.555 84.495 32.725 ;
      RECT 83.865 32.555 84.035 32.725 ;
      RECT 0.605 32.555 0.775 32.725 ;
      RECT 0.145 32.555 0.315 32.725 ;
      RECT 84.325 29.835 84.495 30.005 ;
      RECT 83.865 29.835 84.035 30.005 ;
      RECT 0.605 29.835 0.775 30.005 ;
      RECT 0.145 29.835 0.315 30.005 ;
      RECT 84.325 27.115 84.495 27.285 ;
      RECT 83.865 27.115 84.035 27.285 ;
      RECT 0.605 27.115 0.775 27.285 ;
      RECT 0.145 27.115 0.315 27.285 ;
      RECT 84.325 24.395 84.495 24.565 ;
      RECT 83.865 24.395 84.035 24.565 ;
      RECT 0.605 24.395 0.775 24.565 ;
      RECT 0.145 24.395 0.315 24.565 ;
      RECT 84.325 21.675 84.495 21.845 ;
      RECT 83.865 21.675 84.035 21.845 ;
      RECT 0.605 21.675 0.775 21.845 ;
      RECT 0.145 21.675 0.315 21.845 ;
      RECT 84.325 18.955 84.495 19.125 ;
      RECT 83.865 18.955 84.035 19.125 ;
      RECT 0.605 18.955 0.775 19.125 ;
      RECT 0.145 18.955 0.315 19.125 ;
      RECT 84.325 16.235 84.495 16.405 ;
      RECT 83.865 16.235 84.035 16.405 ;
      RECT 83.405 16.235 83.575 16.405 ;
      RECT 82.945 16.235 83.115 16.405 ;
      RECT 82.485 16.235 82.655 16.405 ;
      RECT 82.025 16.235 82.195 16.405 ;
      RECT 81.565 16.235 81.735 16.405 ;
      RECT 81.105 16.235 81.275 16.405 ;
      RECT 80.645 16.235 80.815 16.405 ;
      RECT 80.185 16.235 80.355 16.405 ;
      RECT 79.725 16.235 79.895 16.405 ;
      RECT 79.265 16.235 79.435 16.405 ;
      RECT 78.805 16.235 78.975 16.405 ;
      RECT 78.345 16.235 78.515 16.405 ;
      RECT 77.885 16.235 78.055 16.405 ;
      RECT 77.425 16.235 77.595 16.405 ;
      RECT 76.965 16.235 77.135 16.405 ;
      RECT 76.505 16.235 76.675 16.405 ;
      RECT 76.045 16.235 76.215 16.405 ;
      RECT 75.585 16.235 75.755 16.405 ;
      RECT 75.125 16.235 75.295 16.405 ;
      RECT 74.665 16.235 74.835 16.405 ;
      RECT 74.205 16.235 74.375 16.405 ;
      RECT 73.745 16.235 73.915 16.405 ;
      RECT 73.285 16.235 73.455 16.405 ;
      RECT 72.825 16.235 72.995 16.405 ;
      RECT 72.365 16.235 72.535 16.405 ;
      RECT 71.905 16.235 72.075 16.405 ;
      RECT 71.445 16.235 71.615 16.405 ;
      RECT 70.985 16.235 71.155 16.405 ;
      RECT 70.525 16.235 70.695 16.405 ;
      RECT 70.065 16.235 70.235 16.405 ;
      RECT 69.605 16.235 69.775 16.405 ;
      RECT 69.145 16.235 69.315 16.405 ;
      RECT 68.685 16.235 68.855 16.405 ;
      RECT 68.225 16.235 68.395 16.405 ;
      RECT 67.765 16.235 67.935 16.405 ;
      RECT 67.305 16.235 67.475 16.405 ;
      RECT 66.845 16.235 67.015 16.405 ;
      RECT 66.385 16.235 66.555 16.405 ;
      RECT 65.925 16.235 66.095 16.405 ;
      RECT 65.465 16.235 65.635 16.405 ;
      RECT 65.005 16.235 65.175 16.405 ;
      RECT 64.545 16.235 64.715 16.405 ;
      RECT 64.085 16.235 64.255 16.405 ;
      RECT 63.625 16.235 63.795 16.405 ;
      RECT 63.165 16.235 63.335 16.405 ;
      RECT 62.705 16.235 62.875 16.405 ;
      RECT 62.245 16.235 62.415 16.405 ;
      RECT 61.785 16.235 61.955 16.405 ;
      RECT 61.325 16.235 61.495 16.405 ;
      RECT 60.865 16.235 61.035 16.405 ;
      RECT 60.405 16.235 60.575 16.405 ;
      RECT 59.945 16.235 60.115 16.405 ;
      RECT 59.485 16.235 59.655 16.405 ;
      RECT 59.025 16.235 59.195 16.405 ;
      RECT 58.565 16.235 58.735 16.405 ;
      RECT 58.105 16.235 58.275 16.405 ;
      RECT 57.645 16.235 57.815 16.405 ;
      RECT 57.185 16.235 57.355 16.405 ;
      RECT 56.725 16.235 56.895 16.405 ;
      RECT 56.265 16.235 56.435 16.405 ;
      RECT 55.805 16.235 55.975 16.405 ;
      RECT 55.345 16.235 55.515 16.405 ;
      RECT 54.885 16.235 55.055 16.405 ;
      RECT 54.425 16.235 54.595 16.405 ;
      RECT 53.965 16.235 54.135 16.405 ;
      RECT 53.505 16.235 53.675 16.405 ;
      RECT 53.045 16.235 53.215 16.405 ;
      RECT 52.585 16.235 52.755 16.405 ;
      RECT 52.125 16.235 52.295 16.405 ;
      RECT 51.665 16.235 51.835 16.405 ;
      RECT 51.205 16.235 51.375 16.405 ;
      RECT 50.745 16.235 50.915 16.405 ;
      RECT 50.285 16.235 50.455 16.405 ;
      RECT 49.825 16.235 49.995 16.405 ;
      RECT 49.365 16.235 49.535 16.405 ;
      RECT 48.905 16.235 49.075 16.405 ;
      RECT 48.445 16.235 48.615 16.405 ;
      RECT 47.985 16.235 48.155 16.405 ;
      RECT 47.525 16.235 47.695 16.405 ;
      RECT 47.065 16.235 47.235 16.405 ;
      RECT 46.605 16.235 46.775 16.405 ;
      RECT 46.145 16.235 46.315 16.405 ;
      RECT 45.685 16.235 45.855 16.405 ;
      RECT 45.225 16.235 45.395 16.405 ;
      RECT 44.765 16.235 44.935 16.405 ;
      RECT 44.305 16.235 44.475 16.405 ;
      RECT 43.845 16.235 44.015 16.405 ;
      RECT 43.385 16.235 43.555 16.405 ;
      RECT 42.925 16.235 43.095 16.405 ;
      RECT 42.465 16.235 42.635 16.405 ;
      RECT 42.005 16.235 42.175 16.405 ;
      RECT 41.545 16.235 41.715 16.405 ;
      RECT 41.085 16.235 41.255 16.405 ;
      RECT 40.625 16.235 40.795 16.405 ;
      RECT 40.165 16.235 40.335 16.405 ;
      RECT 39.705 16.235 39.875 16.405 ;
      RECT 39.245 16.235 39.415 16.405 ;
      RECT 38.785 16.235 38.955 16.405 ;
      RECT 38.325 16.235 38.495 16.405 ;
      RECT 37.865 16.235 38.035 16.405 ;
      RECT 37.405 16.235 37.575 16.405 ;
      RECT 36.945 16.235 37.115 16.405 ;
      RECT 36.485 16.235 36.655 16.405 ;
      RECT 36.025 16.235 36.195 16.405 ;
      RECT 35.565 16.235 35.735 16.405 ;
      RECT 35.105 16.235 35.275 16.405 ;
      RECT 34.645 16.235 34.815 16.405 ;
      RECT 34.185 16.235 34.355 16.405 ;
      RECT 33.725 16.235 33.895 16.405 ;
      RECT 33.265 16.235 33.435 16.405 ;
      RECT 32.805 16.235 32.975 16.405 ;
      RECT 32.345 16.235 32.515 16.405 ;
      RECT 31.885 16.235 32.055 16.405 ;
      RECT 31.425 16.235 31.595 16.405 ;
      RECT 30.965 16.235 31.135 16.405 ;
      RECT 30.505 16.235 30.675 16.405 ;
      RECT 30.045 16.235 30.215 16.405 ;
      RECT 29.585 16.235 29.755 16.405 ;
      RECT 29.125 16.235 29.295 16.405 ;
      RECT 28.665 16.235 28.835 16.405 ;
      RECT 28.205 16.235 28.375 16.405 ;
      RECT 27.745 16.235 27.915 16.405 ;
      RECT 27.285 16.235 27.455 16.405 ;
      RECT 26.825 16.235 26.995 16.405 ;
      RECT 26.365 16.235 26.535 16.405 ;
      RECT 25.905 16.235 26.075 16.405 ;
      RECT 25.445 16.235 25.615 16.405 ;
      RECT 24.985 16.235 25.155 16.405 ;
      RECT 24.525 16.235 24.695 16.405 ;
      RECT 24.065 16.235 24.235 16.405 ;
      RECT 23.605 16.235 23.775 16.405 ;
      RECT 23.145 16.235 23.315 16.405 ;
      RECT 22.685 16.235 22.855 16.405 ;
      RECT 22.225 16.235 22.395 16.405 ;
      RECT 21.765 16.235 21.935 16.405 ;
      RECT 21.305 16.235 21.475 16.405 ;
      RECT 20.845 16.235 21.015 16.405 ;
      RECT 20.385 16.235 20.555 16.405 ;
      RECT 19.925 16.235 20.095 16.405 ;
      RECT 19.465 16.235 19.635 16.405 ;
      RECT 19.005 16.235 19.175 16.405 ;
      RECT 18.545 16.235 18.715 16.405 ;
      RECT 18.085 16.235 18.255 16.405 ;
      RECT 17.625 16.235 17.795 16.405 ;
      RECT 17.165 16.235 17.335 16.405 ;
      RECT 16.705 16.235 16.875 16.405 ;
      RECT 16.245 16.235 16.415 16.405 ;
      RECT 15.785 16.235 15.955 16.405 ;
      RECT 15.325 16.235 15.495 16.405 ;
      RECT 14.865 16.235 15.035 16.405 ;
      RECT 14.405 16.235 14.575 16.405 ;
      RECT 13.945 16.235 14.115 16.405 ;
      RECT 13.485 16.235 13.655 16.405 ;
      RECT 13.025 16.235 13.195 16.405 ;
      RECT 12.565 16.235 12.735 16.405 ;
      RECT 12.105 16.235 12.275 16.405 ;
      RECT 11.645 16.235 11.815 16.405 ;
      RECT 11.185 16.235 11.355 16.405 ;
      RECT 10.725 16.235 10.895 16.405 ;
      RECT 10.265 16.235 10.435 16.405 ;
      RECT 9.805 16.235 9.975 16.405 ;
      RECT 9.345 16.235 9.515 16.405 ;
      RECT 8.885 16.235 9.055 16.405 ;
      RECT 8.425 16.235 8.595 16.405 ;
      RECT 7.965 16.235 8.135 16.405 ;
      RECT 7.505 16.235 7.675 16.405 ;
      RECT 7.045 16.235 7.215 16.405 ;
      RECT 6.585 16.235 6.755 16.405 ;
      RECT 6.125 16.235 6.295 16.405 ;
      RECT 5.665 16.235 5.835 16.405 ;
      RECT 5.205 16.235 5.375 16.405 ;
      RECT 4.745 16.235 4.915 16.405 ;
      RECT 4.285 16.235 4.455 16.405 ;
      RECT 3.825 16.235 3.995 16.405 ;
      RECT 3.365 16.235 3.535 16.405 ;
      RECT 2.905 16.235 3.075 16.405 ;
      RECT 2.445 16.235 2.615 16.405 ;
      RECT 1.985 16.235 2.155 16.405 ;
      RECT 1.525 16.235 1.695 16.405 ;
      RECT 1.065 16.235 1.235 16.405 ;
      RECT 0.605 16.235 0.775 16.405 ;
      RECT 0.145 16.235 0.315 16.405 ;
      RECT 65.925 13.515 66.095 13.685 ;
      RECT 65.465 13.515 65.635 13.685 ;
      RECT 0.605 13.515 0.775 13.685 ;
      RECT 0.145 13.515 0.315 13.685 ;
      RECT 65.925 10.795 66.095 10.965 ;
      RECT 65.465 10.795 65.635 10.965 ;
      RECT 0.605 10.795 0.775 10.965 ;
      RECT 0.145 10.795 0.315 10.965 ;
      RECT 65.925 8.075 66.095 8.245 ;
      RECT 65.465 8.075 65.635 8.245 ;
      RECT 0.605 8.075 0.775 8.245 ;
      RECT 0.145 8.075 0.315 8.245 ;
      RECT 65.925 5.355 66.095 5.525 ;
      RECT 65.465 5.355 65.635 5.525 ;
      RECT 0.605 5.355 0.775 5.525 ;
      RECT 0.145 5.355 0.315 5.525 ;
      RECT 65.925 2.635 66.095 2.805 ;
      RECT 65.465 2.635 65.635 2.805 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 65.925 -0.085 66.095 0.085 ;
      RECT 65.465 -0.085 65.635 0.085 ;
      RECT 65.005 -0.085 65.175 0.085 ;
      RECT 64.545 -0.085 64.715 0.085 ;
      RECT 64.085 -0.085 64.255 0.085 ;
      RECT 63.625 -0.085 63.795 0.085 ;
      RECT 63.165 -0.085 63.335 0.085 ;
      RECT 62.705 -0.085 62.875 0.085 ;
      RECT 62.245 -0.085 62.415 0.085 ;
      RECT 61.785 -0.085 61.955 0.085 ;
      RECT 61.325 -0.085 61.495 0.085 ;
      RECT 60.865 -0.085 61.035 0.085 ;
      RECT 60.405 -0.085 60.575 0.085 ;
      RECT 59.945 -0.085 60.115 0.085 ;
      RECT 59.485 -0.085 59.655 0.085 ;
      RECT 59.025 -0.085 59.195 0.085 ;
      RECT 58.565 -0.085 58.735 0.085 ;
      RECT 58.105 -0.085 58.275 0.085 ;
      RECT 57.645 -0.085 57.815 0.085 ;
      RECT 57.185 -0.085 57.355 0.085 ;
      RECT 56.725 -0.085 56.895 0.085 ;
      RECT 56.265 -0.085 56.435 0.085 ;
      RECT 55.805 -0.085 55.975 0.085 ;
      RECT 55.345 -0.085 55.515 0.085 ;
      RECT 54.885 -0.085 55.055 0.085 ;
      RECT 54.425 -0.085 54.595 0.085 ;
      RECT 53.965 -0.085 54.135 0.085 ;
      RECT 53.505 -0.085 53.675 0.085 ;
      RECT 53.045 -0.085 53.215 0.085 ;
      RECT 52.585 -0.085 52.755 0.085 ;
      RECT 52.125 -0.085 52.295 0.085 ;
      RECT 51.665 -0.085 51.835 0.085 ;
      RECT 51.205 -0.085 51.375 0.085 ;
      RECT 50.745 -0.085 50.915 0.085 ;
      RECT 50.285 -0.085 50.455 0.085 ;
      RECT 49.825 -0.085 49.995 0.085 ;
      RECT 49.365 -0.085 49.535 0.085 ;
      RECT 48.905 -0.085 49.075 0.085 ;
      RECT 48.445 -0.085 48.615 0.085 ;
      RECT 47.985 -0.085 48.155 0.085 ;
      RECT 47.525 -0.085 47.695 0.085 ;
      RECT 47.065 -0.085 47.235 0.085 ;
      RECT 46.605 -0.085 46.775 0.085 ;
      RECT 46.145 -0.085 46.315 0.085 ;
      RECT 45.685 -0.085 45.855 0.085 ;
      RECT 45.225 -0.085 45.395 0.085 ;
      RECT 44.765 -0.085 44.935 0.085 ;
      RECT 44.305 -0.085 44.475 0.085 ;
      RECT 43.845 -0.085 44.015 0.085 ;
      RECT 43.385 -0.085 43.555 0.085 ;
      RECT 42.925 -0.085 43.095 0.085 ;
      RECT 42.465 -0.085 42.635 0.085 ;
      RECT 42.005 -0.085 42.175 0.085 ;
      RECT 41.545 -0.085 41.715 0.085 ;
      RECT 41.085 -0.085 41.255 0.085 ;
      RECT 40.625 -0.085 40.795 0.085 ;
      RECT 40.165 -0.085 40.335 0.085 ;
      RECT 39.705 -0.085 39.875 0.085 ;
      RECT 39.245 -0.085 39.415 0.085 ;
      RECT 38.785 -0.085 38.955 0.085 ;
      RECT 38.325 -0.085 38.495 0.085 ;
      RECT 37.865 -0.085 38.035 0.085 ;
      RECT 37.405 -0.085 37.575 0.085 ;
      RECT 36.945 -0.085 37.115 0.085 ;
      RECT 36.485 -0.085 36.655 0.085 ;
      RECT 36.025 -0.085 36.195 0.085 ;
      RECT 35.565 -0.085 35.735 0.085 ;
      RECT 35.105 -0.085 35.275 0.085 ;
      RECT 34.645 -0.085 34.815 0.085 ;
      RECT 34.185 -0.085 34.355 0.085 ;
      RECT 33.725 -0.085 33.895 0.085 ;
      RECT 33.265 -0.085 33.435 0.085 ;
      RECT 32.805 -0.085 32.975 0.085 ;
      RECT 32.345 -0.085 32.515 0.085 ;
      RECT 31.885 -0.085 32.055 0.085 ;
      RECT 31.425 -0.085 31.595 0.085 ;
      RECT 30.965 -0.085 31.135 0.085 ;
      RECT 30.505 -0.085 30.675 0.085 ;
      RECT 30.045 -0.085 30.215 0.085 ;
      RECT 29.585 -0.085 29.755 0.085 ;
      RECT 29.125 -0.085 29.295 0.085 ;
      RECT 28.665 -0.085 28.835 0.085 ;
      RECT 28.205 -0.085 28.375 0.085 ;
      RECT 27.745 -0.085 27.915 0.085 ;
      RECT 27.285 -0.085 27.455 0.085 ;
      RECT 26.825 -0.085 26.995 0.085 ;
      RECT 26.365 -0.085 26.535 0.085 ;
      RECT 25.905 -0.085 26.075 0.085 ;
      RECT 25.445 -0.085 25.615 0.085 ;
      RECT 24.985 -0.085 25.155 0.085 ;
      RECT 24.525 -0.085 24.695 0.085 ;
      RECT 24.065 -0.085 24.235 0.085 ;
      RECT 23.605 -0.085 23.775 0.085 ;
      RECT 23.145 -0.085 23.315 0.085 ;
      RECT 22.685 -0.085 22.855 0.085 ;
      RECT 22.225 -0.085 22.395 0.085 ;
      RECT 21.765 -0.085 21.935 0.085 ;
      RECT 21.305 -0.085 21.475 0.085 ;
      RECT 20.845 -0.085 21.015 0.085 ;
      RECT 20.385 -0.085 20.555 0.085 ;
      RECT 19.925 -0.085 20.095 0.085 ;
      RECT 19.465 -0.085 19.635 0.085 ;
      RECT 19.005 -0.085 19.175 0.085 ;
      RECT 18.545 -0.085 18.715 0.085 ;
      RECT 18.085 -0.085 18.255 0.085 ;
      RECT 17.625 -0.085 17.795 0.085 ;
      RECT 17.165 -0.085 17.335 0.085 ;
      RECT 16.705 -0.085 16.875 0.085 ;
      RECT 16.245 -0.085 16.415 0.085 ;
      RECT 15.785 -0.085 15.955 0.085 ;
      RECT 15.325 -0.085 15.495 0.085 ;
      RECT 14.865 -0.085 15.035 0.085 ;
      RECT 14.405 -0.085 14.575 0.085 ;
      RECT 13.945 -0.085 14.115 0.085 ;
      RECT 13.485 -0.085 13.655 0.085 ;
      RECT 13.025 -0.085 13.195 0.085 ;
      RECT 12.565 -0.085 12.735 0.085 ;
      RECT 12.105 -0.085 12.275 0.085 ;
      RECT 11.645 -0.085 11.815 0.085 ;
      RECT 11.185 -0.085 11.355 0.085 ;
      RECT 10.725 -0.085 10.895 0.085 ;
      RECT 10.265 -0.085 10.435 0.085 ;
      RECT 9.805 -0.085 9.975 0.085 ;
      RECT 9.345 -0.085 9.515 0.085 ;
      RECT 8.885 -0.085 9.055 0.085 ;
      RECT 8.425 -0.085 8.595 0.085 ;
      RECT 7.965 -0.085 8.135 0.085 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.145 -0.085 0.315 0.085 ;
    LAYER via ;
      RECT 55.125 81.525 55.275 81.675 ;
      RECT 25.685 81.525 25.835 81.675 ;
      RECT 82.265 17.945 82.415 18.095 ;
      RECT 76.745 17.945 76.895 18.095 ;
      RECT 55.125 16.245 55.275 16.395 ;
      RECT 25.685 16.245 25.835 16.395 ;
      RECT 55.125 -0.075 55.275 0.075 ;
      RECT 25.685 -0.075 25.835 0.075 ;
    LAYER via2 ;
      RECT 55.1 81.5 55.3 81.7 ;
      RECT 25.66 81.5 25.86 81.7 ;
      RECT 83.16 50.22 83.36 50.42 ;
      RECT 83.16 44.78 83.36 44.98 ;
      RECT 82.7 40.7 82.9 40.9 ;
      RECT 83.16 31.86 83.36 32.06 ;
      RECT 55.1 -0.1 55.3 0.1 ;
      RECT 25.66 -0.1 25.86 0.1 ;
    LAYER via3 ;
      RECT 55.1 81.5 55.3 81.7 ;
      RECT 25.66 81.5 25.86 81.7 ;
      RECT 55.1 -0.1 55.3 0.1 ;
      RECT 25.66 -0.1 25.86 0.1 ;
    LAYER OVERLAP ;
      POLYGON 0 0 0 81.6 84.64 81.6 84.64 16.32 66.24 16.32 66.24 0 ;
  END
END sb_0__2_

END LIBRARY
