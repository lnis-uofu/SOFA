//Generated from netlist by SpyDrNet
//netlist name: FPGA88_SOFA_A
module sky130_fd_sc_hd__dfrtp_1
(
    CLK,
    D,
    RESET_B,
    Q
);

    input CLK;
    input D;
    input RESET_B;
    output Q;

    wire CLK;
    wire D;
    wire Q;
    wire RESET_B;

endmodule

