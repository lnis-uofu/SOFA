VERSION 5.7 ;
BUSBITCHARS "[]" ;

UNITS
  DATABASE MICRONS 1000 ;
END UNITS

MANUFACTURINGGRID 0.005 ;

LAYER li1
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.46 ;
  WIDTH 0.17 ;
END li1

LAYER mcon
  TYPE CUT ;
END mcon

LAYER met1
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.34 ;
  WIDTH 0.14 ;
END met1

LAYER via
  TYPE CUT ;
END via

LAYER met2
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.46 ;
  WIDTH 0.14 ;
END met2

LAYER via2
  TYPE CUT ;
END via2

LAYER met3
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.68 ;
  WIDTH 0.3 ;
END met3

LAYER via3
  TYPE CUT ;
END via3

LAYER met4
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.92 ;
  WIDTH 0.3 ;
END met4

LAYER via4
  TYPE CUT ;
END via4

LAYER met5
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 3.4 ;
  WIDTH 1.6 ;
END met5

LAYER nwell
  TYPE MASTERSLICE ;
END nwell

LAYER pwell
  TYPE MASTERSLICE ;
END pwell

LAYER OVERLAP
  TYPE OVERLAP ;
END OVERLAP

VIA L1M1_PR
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.145 -0.115 0.145 0.115 ;
END L1M1_PR

VIA L1M1_PR_R
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.115 -0.145 0.115 0.145 ;
END L1M1_PR_R

VIA L1M1_PR_M
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.115 -0.145 0.115 0.145 ;
END L1M1_PR_M

VIA L1M1_PR_MR
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.145 -0.115 0.145 0.115 ;
END L1M1_PR_MR

VIA L1M1_PR_C
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.145 -0.145 0.145 0.145 ;
END L1M1_PR_C

VIA M1M2_PR
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR

VIA M1M2_PR_Enc
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_Enc

VIA M1M2_PR_R
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_R

VIA M1M2_PR_R_Enc
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR_R_Enc

VIA M1M2_PR_M
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_M

VIA M1M2_PR_M_Enc
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR_M_Enc

VIA M1M2_PR_MR
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR_MR

VIA M1M2_PR_MR_Enc
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_MR_Enc

VIA M1M2_PR_C
  LAYER met1 ;
    RECT -0.16 -0.16 0.16 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.16 0.16 0.16 ;
END M1M2_PR_C

VIA M2M3_PR
  LAYER met2 ;
    RECT -0.14 -0.185 0.14 0.185 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR

VIA M2M3_PR_R
  LAYER met2 ;
    RECT -0.185 -0.14 0.185 0.14 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_R

VIA M2M3_PR_M
  LAYER met2 ;
    RECT -0.14 -0.185 0.14 0.185 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_M

VIA M2M3_PR_MR
  LAYER met2 ;
    RECT -0.185 -0.14 0.185 0.14 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_MR

VIA M2M3_PR_C
  LAYER met2 ;
    RECT -0.185 -0.185 0.185 0.185 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_C

VIA M3M4_PR
  LAYER met3 ;
    RECT -0.19 -0.16 0.19 0.16 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR

VIA M3M4_PR_R
  LAYER met3 ;
    RECT -0.16 -0.19 0.16 0.19 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_R

VIA M3M4_PR_M
  LAYER met3 ;
    RECT -0.19 -0.16 0.19 0.16 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_M

VIA M3M4_PR_MR
  LAYER met3 ;
    RECT -0.16 -0.19 0.16 0.19 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_MR

VIA M3M4_PR_C
  LAYER met3 ;
    RECT -0.19 -0.19 0.19 0.19 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_C

VIA M4M5_PR
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR

VIA M4M5_PR_R
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_R

VIA M4M5_PR_M
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_M

VIA M4M5_PR_MR
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_MR

VIA M4M5_PR_C
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_C

SITE unit
  CLASS CORE ;
  SYMMETRY Y ;
  SIZE 0.46 BY 2.72 ;
END unit

SITE unithddbl
  CLASS CORE ;
  SIZE 0.46 BY 5.44 ;
END unithddbl

MACRO sb_1__1_
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  SIZE 117.76 BY 108.8 ;
  SYMMETRY X Y ;
  PIN chany_top_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 63.79 108 64.09 108.8 ;
    END
  END chany_top_in[0]
  PIN chany_top_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.34 108.315 84.48 108.8 ;
    END
  END chany_top_in[1]
  PIN chany_top_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.42 108.315 83.56 108.8 ;
    END
  END chany_top_in[2]
  PIN chany_top_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 73.91 108 74.21 108.8 ;
    END
  END chany_top_in[3]
  PIN chany_top_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.58 108.315 81.72 108.8 ;
    END
  END chany_top_in[4]
  PIN chany_top_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 56.43 108 56.73 108.8 ;
    END
  END chany_top_in[5]
  PIN chany_top_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.36 108.315 55.5 108.8 ;
    END
  END chany_top_in[6]
  PIN chany_top_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 60.11 108 60.41 108.8 ;
    END
  END chany_top_in[7]
  PIN chany_top_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.26 108.315 85.4 108.8 ;
    END
  END chany_top_in[8]
  PIN chany_top_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.02 108.315 88.16 108.8 ;
    END
  END chany_top_in[9]
  PIN chany_top_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.5 108.315 82.64 108.8 ;
    END
  END chany_top_in[10]
  PIN chany_top_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.94 108.315 89.08 108.8 ;
    END
  END chany_top_in[11]
  PIN chany_top_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 67.47 108 67.77 108.8 ;
    END
  END chany_top_in[12]
  PIN chany_top_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.32 108.315 67.46 108.8 ;
    END
  END chany_top_in[13]
  PIN chany_top_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 52.75 108 53.05 108.8 ;
    END
  END chany_top_in[14]
  PIN chany_top_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 58.27 108 58.57 108.8 ;
    END
  END chany_top_in[15]
  PIN chany_top_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.58 108.315 58.72 108.8 ;
    END
  END chany_top_in[16]
  PIN chany_top_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 54.59 108 54.89 108.8 ;
    END
  END chany_top_in[17]
  PIN chany_top_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.1 108.315 64.24 108.8 ;
    END
  END chany_top_in[18]
  PIN chany_top_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 69.31 108 69.61 108.8 ;
    END
  END chany_top_in[19]
  PIN top_left_grid_pin_42_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.5 97.435 13.64 97.92 ;
    END
  END top_left_grid_pin_42_[0]
  PIN top_left_grid_pin_43_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.66 97.435 11.8 97.92 ;
    END
  END top_left_grid_pin_43_[0]
  PIN top_left_grid_pin_44_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.44 97.435 8.58 97.92 ;
    END
  END top_left_grid_pin_44_[0]
  PIN top_left_grid_pin_45_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.58 97.435 12.72 97.92 ;
    END
  END top_left_grid_pin_45_[0]
  PIN top_left_grid_pin_46_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.28 97.435 10.42 97.92 ;
    END
  END top_left_grid_pin_46_[0]
  PIN top_left_grid_pin_47_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.3 97.435 4.44 97.92 ;
    END
  END top_left_grid_pin_47_[0]
  PIN top_left_grid_pin_48_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.36 97.435 9.5 97.92 ;
    END
  END top_left_grid_pin_48_[0]
  PIN top_left_grid_pin_49_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.06 97.435 7.2 97.92 ;
    END
  END top_left_grid_pin_49_[0]
  PIN chanx_right_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.96 66.15 117.76 66.45 ;
    END
  END chanx_right_in[0]
  PIN chanx_right_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.96 87.91 117.76 88.21 ;
    END
  END chanx_right_in[1]
  PIN chanx_right_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.96 36.23 117.76 36.53 ;
    END
  END chanx_right_in[2]
  PIN chanx_right_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.96 48.47 117.76 48.77 ;
    END
  END chanx_right_in[3]
  PIN chanx_right_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.96 71.59 117.76 71.89 ;
    END
  END chanx_right_in[4]
  PIN chanx_right_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.96 86.55 117.76 86.85 ;
    END
  END chanx_right_in[5]
  PIN chanx_right_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.96 62.07 117.76 62.37 ;
    END
  END chanx_right_in[6]
  PIN chanx_right_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.96 22.63 117.76 22.93 ;
    END
  END chanx_right_in[7]
  PIN chanx_right_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.96 34.87 117.76 35.17 ;
    END
  END chanx_right_in[8]
  PIN chanx_right_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.96 41.67 117.76 41.97 ;
    END
  END chanx_right_in[9]
  PIN chanx_right_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.96 64.79 117.76 65.09 ;
    END
  END chanx_right_in[10]
  PIN chanx_right_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.96 51.19 117.76 51.49 ;
    END
  END chanx_right_in[11]
  PIN chanx_right_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.96 23.99 117.76 24.29 ;
    END
  END chanx_right_in[12]
  PIN chanx_right_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.96 44.39 117.76 44.69 ;
    END
  END chanx_right_in[13]
  PIN chanx_right_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.96 60.71 117.76 61.01 ;
    END
  END chanx_right_in[14]
  PIN chanx_right_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.96 57.99 117.76 58.29 ;
    END
  END chanx_right_in[15]
  PIN chanx_right_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.96 67.51 117.76 67.81 ;
    END
  END chanx_right_in[16]
  PIN chanx_right_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.96 45.75 117.76 46.05 ;
    END
  END chanx_right_in[17]
  PIN chanx_right_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.96 63.43 117.76 63.73 ;
    END
  END chanx_right_in[18]
  PIN chanx_right_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.96 43.03 117.76 43.33 ;
    END
  END chanx_right_in[19]
  PIN right_bottom_grid_pin_34_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.04 10.88 105.18 11.365 ;
    END
  END right_bottom_grid_pin_34_[0]
  PIN right_bottom_grid_pin_35_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.48 10.88 111.62 11.365 ;
    END
  END right_bottom_grid_pin_35_[0]
  PIN right_bottom_grid_pin_36_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.8 10.88 107.94 11.365 ;
    END
  END right_bottom_grid_pin_36_[0]
  PIN right_bottom_grid_pin_37_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.86 10.88 113 11.365 ;
    END
  END right_bottom_grid_pin_37_[0]
  PIN right_bottom_grid_pin_38_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.88 10.88 107.02 11.365 ;
    END
  END right_bottom_grid_pin_38_[0]
  PIN right_bottom_grid_pin_39_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.12 10.88 104.26 11.365 ;
    END
  END right_bottom_grid_pin_39_[0]
  PIN right_bottom_grid_pin_40_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.96 10.88 106.1 11.365 ;
    END
  END right_bottom_grid_pin_40_[0]
  PIN right_bottom_grid_pin_41_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.72 10.88 108.86 11.365 ;
    END
  END right_bottom_grid_pin_41_[0]
  PIN chany_bottom_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.4 0 89.54 0.485 ;
    END
  END chany_bottom_in[0]
  PIN chany_bottom_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 52.75 0 53.05 0.8 ;
    END
  END chany_bottom_in[1]
  PIN chany_bottom_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.34 0 84.48 0.485 ;
    END
  END chany_bottom_in[2]
  PIN chany_bottom_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.2 0 80.34 0.485 ;
    END
  END chany_bottom_in[3]
  PIN chany_bottom_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.58 0 81.72 0.485 ;
    END
  END chany_bottom_in[4]
  PIN chany_bottom_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.26 0 39.4 0.485 ;
    END
  END chany_bottom_in[5]
  PIN chany_bottom_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 74.83 0 75.13 0.8 ;
    END
  END chany_bottom_in[6]
  PIN chany_bottom_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.66 0 34.8 0.485 ;
    END
  END chany_bottom_in[7]
  PIN chany_bottom_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.28 0 79.42 0.485 ;
    END
  END chany_bottom_in[8]
  PIN chany_bottom_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.86 0 67 0.485 ;
    END
  END chany_bottom_in[9]
  PIN chany_bottom_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.98 0 77.12 0.485 ;
    END
  END chany_bottom_in[10]
  PIN chany_bottom_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.14 0 75.28 0.485 ;
    END
  END chany_bottom_in[11]
  PIN chany_bottom_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.18 0 86.32 0.485 ;
    END
  END chany_bottom_in[12]
  PIN chany_bottom_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.18 0 40.32 0.485 ;
    END
  END chany_bottom_in[13]
  PIN chany_bottom_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.82 0 32.96 0.485 ;
    END
  END chany_bottom_in[14]
  PIN chany_bottom_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.5 0 36.64 0.485 ;
    END
  END chany_bottom_in[15]
  PIN chany_bottom_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.5 0 82.64 0.485 ;
    END
  END chany_bottom_in[16]
  PIN chany_bottom_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.66 0 57.8 0.485 ;
    END
  END chany_bottom_in[17]
  PIN chany_bottom_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.26 0 62.4 0.485 ;
    END
  END chany_bottom_in[18]
  PIN chany_bottom_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.82 0 55.96 0.485 ;
    END
  END chany_bottom_in[19]
  PIN bottom_left_grid_pin_42_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.42 10.88 14.56 11.365 ;
    END
  END bottom_left_grid_pin_42_[0]
  PIN bottom_left_grid_pin_43_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.34 10.88 15.48 11.365 ;
    END
  END bottom_left_grid_pin_43_[0]
  PIN bottom_left_grid_pin_44_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.92 10.88 3.06 11.365 ;
    END
  END bottom_left_grid_pin_44_[0]
  PIN bottom_left_grid_pin_45_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.28 10.88 10.42 11.365 ;
    END
  END bottom_left_grid_pin_45_[0]
  PIN bottom_left_grid_pin_46_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.22 10.88 5.36 11.365 ;
    END
  END bottom_left_grid_pin_46_[0]
  PIN bottom_left_grid_pin_47_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.3 10.88 4.44 11.365 ;
    END
  END bottom_left_grid_pin_47_[0]
  PIN bottom_left_grid_pin_48_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.5 10.88 13.64 11.365 ;
    END
  END bottom_left_grid_pin_48_[0]
  PIN bottom_left_grid_pin_49_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.06 10.88 7.2 11.365 ;
    END
  END bottom_left_grid_pin_49_[0]
  PIN chanx_left_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 59.35 0.8 59.65 ;
    END
  END chanx_left_in[0]
  PIN chanx_left_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 53.91 0.8 54.21 ;
    END
  END chanx_left_in[1]
  PIN chanx_left_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 62.07 0.8 62.37 ;
    END
  END chanx_left_in[2]
  PIN chanx_left_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 56.63 0.8 56.93 ;
    END
  END chanx_left_in[3]
  PIN chanx_left_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 22.63 0.8 22.93 ;
    END
  END chanx_left_in[4]
  PIN chanx_left_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 47.11 0.8 47.41 ;
    END
  END chanx_left_in[5]
  PIN chanx_left_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 43.03 0.8 43.33 ;
    END
  END chanx_left_in[6]
  PIN chanx_left_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 48.47 0.8 48.77 ;
    END
  END chanx_left_in[7]
  PIN chanx_left_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 66.83 0.8 67.13 ;
    END
  END chanx_left_in[8]
  PIN chanx_left_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 72.27 0.8 72.57 ;
    END
  END chanx_left_in[9]
  PIN chanx_left_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 41.67 0.8 41.97 ;
    END
  END chanx_left_in[10]
  PIN chanx_left_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 57.99 0.8 58.29 ;
    END
  END chanx_left_in[11]
  PIN chanx_left_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 60.71 0.8 61.01 ;
    END
  END chanx_left_in[12]
  PIN chanx_left_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 87.91 0.8 88.21 ;
    END
  END chanx_left_in[13]
  PIN chanx_left_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 45.75 0.8 46.05 ;
    END
  END chanx_left_in[14]
  PIN chanx_left_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 69.55 0.8 69.85 ;
    END
  END chanx_left_in[15]
  PIN chanx_left_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 63.43 0.8 63.73 ;
    END
  END chanx_left_in[16]
  PIN chanx_left_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 70.91 0.8 71.21 ;
    END
  END chanx_left_in[17]
  PIN chanx_left_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 85.19 0.8 85.49 ;
    END
  END chanx_left_in[18]
  PIN chanx_left_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 68.19 0.8 68.49 ;
    END
  END chanx_left_in[19]
  PIN left_bottom_grid_pin_34_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 6.75 10.88 7.05 11.68 ;
    END
  END left_bottom_grid_pin_34_[0]
  PIN left_bottom_grid_pin_35_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 8.59 10.88 8.89 11.68 ;
    END
  END left_bottom_grid_pin_35_[0]
  PIN left_bottom_grid_pin_36_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.9 10.88 9.04 11.365 ;
    END
  END left_bottom_grid_pin_36_[0]
  PIN left_bottom_grid_pin_37_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.98 10.88 8.12 11.365 ;
    END
  END left_bottom_grid_pin_37_[0]
  PIN left_bottom_grid_pin_38_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.66 10.88 11.8 11.365 ;
    END
  END left_bottom_grid_pin_38_[0]
  PIN left_bottom_grid_pin_39_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.58 10.88 12.72 11.365 ;
    END
  END left_bottom_grid_pin_39_[0]
  PIN left_bottom_grid_pin_40_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.22 0 28.36 0.485 ;
    END
  END left_bottom_grid_pin_40_[0]
  PIN left_bottom_grid_pin_41_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.14 10.88 6.28 11.365 ;
    END
  END left_bottom_grid_pin_41_[0]
  PIN ccff_head[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.96 29.43 117.76 29.73 ;
    END
  END ccff_head[0]
  PIN chany_top_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71 108.315 71.14 108.8 ;
    END
  END chany_top_out[0]
  PIN chany_top_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.44 108.315 77.58 108.8 ;
    END
  END chany_top_out[1]
  PIN chany_top_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.68 108.315 74.82 108.8 ;
    END
  END chany_top_out[2]
  PIN chany_top_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.36 108.315 78.5 108.8 ;
    END
  END chany_top_out[3]
  PIN chany_top_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.26 108.315 39.4 108.8 ;
    END
  END chany_top_out[4]
  PIN chany_top_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.42 108.315 60.56 108.8 ;
    END
  END chany_top_out[5]
  PIN chany_top_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.44 108.315 54.58 108.8 ;
    END
  END chany_top_out[6]
  PIN chany_top_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.76 108.315 50.9 108.8 ;
    END
  END chany_top_out[7]
  PIN chany_top_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.4 108.315 66.54 108.8 ;
    END
  END chany_top_out[8]
  PIN chany_top_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.28 108.315 79.42 108.8 ;
    END
  END chany_top_out[9]
  PIN chany_top_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.66 108.315 57.8 108.8 ;
    END
  END chany_top_out[10]
  PIN chany_top_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.18 108.315 63.32 108.8 ;
    END
  END chany_top_out[11]
  PIN chany_top_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.16 108.315 69.3 108.8 ;
    END
  END chany_top_out[12]
  PIN chany_top_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.52 108.315 76.66 108.8 ;
    END
  END chany_top_out[13]
  PIN chany_top_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.14 108.315 52.28 108.8 ;
    END
  END chany_top_out[14]
  PIN chany_top_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.02 108.315 65.16 108.8 ;
    END
  END chany_top_out[15]
  PIN chany_top_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.06 108.315 53.2 108.8 ;
    END
  END chany_top_out[16]
  PIN chany_top_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.08 108.315 70.22 108.8 ;
    END
  END chany_top_out[17]
  PIN chany_top_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.5 108.315 59.64 108.8 ;
    END
  END chany_top_out[18]
  PIN chany_top_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.6 108.315 75.74 108.8 ;
    END
  END chany_top_out[19]
  PIN chanx_right_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.96 70.23 117.76 70.53 ;
    END
  END chanx_right_out[0]
  PIN chanx_right_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.96 72.95 117.76 73.25 ;
    END
  END chanx_right_out[1]
  PIN chanx_right_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.96 25.35 117.76 25.65 ;
    END
  END chanx_right_out[2]
  PIN chanx_right_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.96 49.83 117.76 50.13 ;
    END
  END chanx_right_out[3]
  PIN chanx_right_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.96 56.63 117.76 56.93 ;
    END
  END chanx_right_out[4]
  PIN chanx_right_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.96 53.91 117.76 54.21 ;
    END
  END chanx_right_out[5]
  PIN chanx_right_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.96 85.19 117.76 85.49 ;
    END
  END chanx_right_out[6]
  PIN chanx_right_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.96 33.51 117.76 33.81 ;
    END
  END chanx_right_out[7]
  PIN chanx_right_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.96 32.15 117.76 32.45 ;
    END
  END chanx_right_out[8]
  PIN chanx_right_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.96 55.27 117.76 55.57 ;
    END
  END chanx_right_out[9]
  PIN chanx_right_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.96 26.71 117.76 27.01 ;
    END
  END chanx_right_out[10]
  PIN chanx_right_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.96 52.55 117.76 52.85 ;
    END
  END chanx_right_out[11]
  PIN chanx_right_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.96 15.83 117.76 16.13 ;
    END
  END chanx_right_out[12]
  PIN chanx_right_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.96 47.11 117.76 47.41 ;
    END
  END chanx_right_out[13]
  PIN chanx_right_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.96 30.79 117.76 31.09 ;
    END
  END chanx_right_out[14]
  PIN chanx_right_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.96 68.87 117.76 69.17 ;
    END
  END chanx_right_out[15]
  PIN chanx_right_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.96 14.47 117.76 14.77 ;
    END
  END chanx_right_out[16]
  PIN chanx_right_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.96 59.35 117.76 59.65 ;
    END
  END chanx_right_out[17]
  PIN chanx_right_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.96 28.07 117.76 28.37 ;
    END
  END chanx_right_out[18]
  PIN chanx_right_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.96 89.27 117.76 89.57 ;
    END
  END chanx_right_out[19]
  PIN chany_bottom_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.94 0 66.08 0.485 ;
    END
  END chany_bottom_out[0]
  PIN chany_bottom_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.26 0 85.4 0.485 ;
    END
  END chany_bottom_out[1]
  PIN chany_bottom_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.58 0 35.72 0.485 ;
    END
  END chany_bottom_out[2]
  PIN chany_bottom_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.42 0 83.56 0.485 ;
    END
  END chany_bottom_out[3]
  PIN chany_bottom_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.34 0 38.48 0.485 ;
    END
  END chany_bottom_out[4]
  PIN chany_bottom_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.3 0 73.44 0.485 ;
    END
  END chany_bottom_out[5]
  PIN chany_bottom_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.06 0 76.2 0.485 ;
    END
  END chany_bottom_out[6]
  PIN chany_bottom_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.42 0 37.56 0.485 ;
    END
  END chany_bottom_out[7]
  PIN chany_bottom_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.42 0 60.56 0.485 ;
    END
  END chany_bottom_out[8]
  PIN chany_bottom_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.1 0 64.24 0.485 ;
    END
  END chany_bottom_out[9]
  PIN chany_bottom_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.78 0 67.92 0.485 ;
    END
  END chany_bottom_out[10]
  PIN chany_bottom_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.22 0 74.36 0.485 ;
    END
  END chany_bottom_out[11]
  PIN chany_bottom_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.5 0 59.64 0.485 ;
    END
  END chany_bottom_out[12]
  PIN chany_bottom_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.9 0 55.04 0.485 ;
    END
  END chany_bottom_out[13]
  PIN chany_bottom_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.98 0 54.12 0.485 ;
    END
  END chany_bottom_out[14]
  PIN chany_bottom_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.02 0 65.16 0.485 ;
    END
  END chany_bottom_out[15]
  PIN chany_bottom_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.58 0 58.72 0.485 ;
    END
  END chany_bottom_out[16]
  PIN chany_bottom_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.18 0 63.32 0.485 ;
    END
  END chany_bottom_out[17]
  PIN chany_bottom_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.14 0 52.28 0.485 ;
    END
  END chany_bottom_out[18]
  PIN chany_bottom_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.06 0 53.2 0.485 ;
    END
  END chany_bottom_out[19]
  PIN chanx_left_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 23.99 0.8 24.29 ;
    END
  END chanx_left_out[0]
  PIN chanx_left_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 64.79 0.8 65.09 ;
    END
  END chanx_left_out[1]
  PIN chanx_left_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 34.87 0.8 35.17 ;
    END
  END chanx_left_out[2]
  PIN chanx_left_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 55.27 0.8 55.57 ;
    END
  END chanx_left_out[3]
  PIN chanx_left_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 15.83 0.8 16.13 ;
    END
  END chanx_left_out[4]
  PIN chanx_left_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 44.39 0.8 44.69 ;
    END
  END chanx_left_out[5]
  PIN chanx_left_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 33.51 0.8 33.81 ;
    END
  END chanx_left_out[6]
  PIN chanx_left_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 25.35 0.8 25.65 ;
    END
  END chanx_left_out[7]
  PIN chanx_left_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 30.79 0.8 31.09 ;
    END
  END chanx_left_out[8]
  PIN chanx_left_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 49.83 0.8 50.13 ;
    END
  END chanx_left_out[9]
  PIN chanx_left_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 36.23 0.8 36.53 ;
    END
  END chanx_left_out[10]
  PIN chanx_left_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 52.55 0.8 52.85 ;
    END
  END chanx_left_out[11]
  PIN chanx_left_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 17.19 0.8 17.49 ;
    END
  END chanx_left_out[12]
  PIN chanx_left_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 86.55 0.8 86.85 ;
    END
  END chanx_left_out[13]
  PIN chanx_left_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 37.59 0.8 37.89 ;
    END
  END chanx_left_out[14]
  PIN chanx_left_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 28.07 0.8 28.37 ;
    END
  END chanx_left_out[15]
  PIN chanx_left_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 14.47 0.8 14.77 ;
    END
  END chanx_left_out[16]
  PIN chanx_left_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 51.19 0.8 51.49 ;
    END
  END chanx_left_out[17]
  PIN chanx_left_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 32.15 0.8 32.45 ;
    END
  END chanx_left_out[18]
  PIN chanx_left_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 26.71 0.8 27.01 ;
    END
  END chanx_left_out[19]
  PIN ccff_tail[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 29.43 0.8 29.73 ;
    END
  END ccff_tail[0]
  PIN Test_en_S_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.36 0 78.5 0.485 ;
    END
  END Test_en_S_in
  PIN Test_en_N_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.76 108.315 73.9 108.8 ;
    END
  END Test_en_N_out
  PIN prog_clk_0_N_in
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER met2 ;
        RECT 38.34 108.315 38.48 108.8 ;
    END
  END prog_clk_0_N_in
  PIN prog_clk_1_N_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.34 108.315 61.48 108.8 ;
    END
  END prog_clk_1_N_in
  PIN prog_clk_1_S_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.34 0 61.48 0.485 ;
    END
  END prog_clk_1_S_in
  PIN prog_clk_1_E_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.96 37.59 117.76 37.89 ;
    END
  END prog_clk_1_E_out
  PIN prog_clk_1_W_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 40.31 0.8 40.61 ;
    END
  END prog_clk_1_W_out
  PIN prog_clk_2_N_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.38 108.315 72.52 108.8 ;
    END
  END prog_clk_2_N_in
  PIN prog_clk_2_E_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.96 82.47 117.76 82.77 ;
    END
  END prog_clk_2_E_in
  PIN prog_clk_2_S_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 70.23 0 70.53 0.8 ;
    END
  END prog_clk_2_S_in
  PIN prog_clk_2_W_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 74.99 0.8 75.29 ;
    END
  END prog_clk_2_W_in
  PIN prog_clk_2_W_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 73.63 0.8 73.93 ;
    END
  END prog_clk_2_W_out
  PIN prog_clk_2_S_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.16 0 69.3 0.485 ;
    END
  END prog_clk_2_S_out
  PIN prog_clk_2_N_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.1 108.315 87.24 108.8 ;
    END
  END prog_clk_2_N_out
  PIN prog_clk_2_E_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.96 74.31 117.76 74.61 ;
    END
  END prog_clk_2_E_out
  PIN prog_clk_3_W_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 76.35 0.8 76.65 ;
    END
  END prog_clk_3_W_in
  PIN prog_clk_3_E_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.96 77.03 117.76 77.33 ;
    END
  END prog_clk_3_E_in
  PIN prog_clk_3_S_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.56 0 87.7 0.485 ;
    END
  END prog_clk_3_S_in
  PIN prog_clk_3_N_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 72.07 108 72.37 108.8 ;
    END
  END prog_clk_3_N_in
  PIN prog_clk_3_E_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.96 81.11 117.76 81.41 ;
    END
  END prog_clk_3_E_out
  PIN prog_clk_3_W_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 81.79 0.8 82.09 ;
    END
  END prog_clk_3_W_out
  PIN prog_clk_3_N_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.18 108.315 86.32 108.8 ;
    END
  END prog_clk_3_N_out
  PIN prog_clk_3_S_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.08 0 70.22 0.485 ;
    END
  END prog_clk_3_S_out
  PIN clk_1_N_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.74 108.315 56.88 108.8 ;
    END
  END clk_1_N_in
  PIN clk_1_S_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.74 0 56.88 0.485 ;
    END
  END clk_1_S_in
  PIN clk_1_E_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.96 38.95 117.76 39.25 ;
    END
  END clk_1_E_out
  PIN clk_1_W_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 38.95 0.8 39.25 ;
    END
  END clk_1_W_out
  PIN clk_2_N_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 61.95 108 62.25 108.8 ;
    END
  END clk_2_N_in
  PIN clk_2_E_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.96 83.83 117.76 84.13 ;
    END
  END clk_2_E_in
  PIN clk_2_S_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 72.07 0 72.37 0.8 ;
    END
  END clk_2_S_in
  PIN clk_2_W_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 77.71 0.8 78.01 ;
    END
  END clk_2_W_in
  PIN clk_2_W_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 83.83 0.8 84.13 ;
    END
  END clk_2_W_out
  PIN clk_2_S_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71 0 71.14 0.485 ;
    END
  END clk_2_S_out
  PIN clk_2_N_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.2 108.315 80.34 108.8 ;
    END
  END clk_2_N_out
  PIN clk_2_E_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.96 75.67 117.76 75.97 ;
    END
  END clk_2_E_out
  PIN clk_3_W_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 79.07 0.8 79.37 ;
    END
  END clk_3_W_in
  PIN clk_3_E_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.96 79.75 117.76 80.05 ;
    END
  END clk_3_E_in
  PIN clk_3_S_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.48 0 88.62 0.485 ;
    END
  END clk_3_S_in
  PIN clk_3_N_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.26 108.315 62.4 108.8 ;
    END
  END clk_3_N_in
  PIN clk_3_E_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 116.96 78.39 117.76 78.69 ;
    END
  END clk_3_E_out
  PIN clk_3_W_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 80.43 0.8 80.73 ;
    END
  END clk_3_W_out
  PIN clk_3_N_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.24 108.315 68.38 108.8 ;
    END
  END clk_3_N_out
  PIN clk_3_S_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.38 0 72.52 0.485 ;
    END
  END clk_3_S_out
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 25.76 2.48 26.24 2.96 ;
        RECT 91.52 2.48 92 2.96 ;
        RECT 25.76 7.92 26.24 8.4 ;
        RECT 91.52 7.92 92 8.4 ;
        RECT 0 13.36 0.48 13.84 ;
        RECT 117.28 13.36 117.76 13.84 ;
        RECT 0 18.8 0.48 19.28 ;
        RECT 117.28 18.8 117.76 19.28 ;
        RECT 0 24.24 0.48 24.72 ;
        RECT 117.28 24.24 117.76 24.72 ;
        RECT 0 29.68 0.48 30.16 ;
        RECT 117.28 29.68 117.76 30.16 ;
        RECT 0 35.12 0.48 35.6 ;
        RECT 117.28 35.12 117.76 35.6 ;
        RECT 0 40.56 0.48 41.04 ;
        RECT 117.28 40.56 117.76 41.04 ;
        RECT 0 46 0.48 46.48 ;
        RECT 117.28 46 117.76 46.48 ;
        RECT 0 51.44 0.48 51.92 ;
        RECT 117.28 51.44 117.76 51.92 ;
        RECT 0 56.88 0.48 57.36 ;
        RECT 117.28 56.88 117.76 57.36 ;
        RECT 0 62.32 0.48 62.8 ;
        RECT 117.28 62.32 117.76 62.8 ;
        RECT 0 67.76 0.48 68.24 ;
        RECT 117.28 67.76 117.76 68.24 ;
        RECT 0 73.2 0.48 73.68 ;
        RECT 117.28 73.2 117.76 73.68 ;
        RECT 0 78.64 0.48 79.12 ;
        RECT 117.28 78.64 117.76 79.12 ;
        RECT 0 84.08 0.48 84.56 ;
        RECT 117.28 84.08 117.76 84.56 ;
        RECT 0 89.52 0.48 90 ;
        RECT 117.28 89.52 117.76 90 ;
        RECT 0 94.96 0.48 95.44 ;
        RECT 117.28 94.96 117.76 95.44 ;
        RECT 25.76 100.4 26.24 100.88 ;
        RECT 91.52 100.4 92 100.88 ;
        RECT 25.76 105.84 26.24 106.32 ;
        RECT 91.52 105.84 92 106.32 ;
      LAYER met5 ;
        RECT 0 22.2 3.2 25.4 ;
        RECT 114.56 22.2 117.76 25.4 ;
        RECT 0 63 3.2 66.2 ;
        RECT 114.56 63 117.76 66.2 ;
      LAYER met4 ;
        RECT 36.5 0 37.1 0.6 ;
        RECT 65.94 0 66.54 0.6 ;
        RECT 106.42 10.88 107.02 11.48 ;
        RECT 106.42 97.32 107.02 97.92 ;
        RECT 36.5 108.2 37.1 108.8 ;
        RECT 65.94 108.2 66.54 108.8 ;
    END
  END VDD
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 25.76 0 45.4 0.24 ;
        RECT 46.6 0 92 0.24 ;
        RECT 25.76 5.2 26.24 5.68 ;
        RECT 91.52 5.2 92 5.68 ;
        RECT 0 10.64 45.4 11.12 ;
        RECT 46.6 10.64 95.08 11.12 ;
        RECT 96.28 10.88 117.76 11.12 ;
        RECT 0 16.08 0.48 16.56 ;
        RECT 117.28 16.08 117.76 16.56 ;
        RECT 0 21.52 0.48 22 ;
        RECT 117.28 21.52 117.76 22 ;
        RECT 0 26.96 0.48 27.44 ;
        RECT 117.28 26.96 117.76 27.44 ;
        RECT 0 32.4 0.48 32.88 ;
        RECT 117.28 32.4 117.76 32.88 ;
        RECT 0 37.84 0.48 38.32 ;
        RECT 117.28 37.84 117.76 38.32 ;
        RECT 0 43.28 0.48 43.76 ;
        RECT 117.28 43.28 117.76 43.76 ;
        RECT 0 48.72 0.48 49.2 ;
        RECT 117.28 48.72 117.76 49.2 ;
        RECT 0 54.16 0.48 54.64 ;
        RECT 117.28 54.16 117.76 54.64 ;
        RECT 0 59.6 0.48 60.08 ;
        RECT 117.28 59.6 117.76 60.08 ;
        RECT 0 65.04 0.48 65.52 ;
        RECT 117.28 65.04 117.76 65.52 ;
        RECT 0 70.48 0.48 70.96 ;
        RECT 117.28 70.48 117.76 70.96 ;
        RECT 0 75.92 0.48 76.4 ;
        RECT 117.28 75.92 117.76 76.4 ;
        RECT 0 81.36 0.48 81.84 ;
        RECT 117.28 81.36 117.76 81.84 ;
        RECT 0 86.8 0.48 87.28 ;
        RECT 117.28 86.8 117.76 87.28 ;
        RECT 0 92.24 0.48 92.72 ;
        RECT 117.28 92.24 117.76 92.72 ;
        RECT 96.28 97.68 117.76 97.92 ;
        RECT 0 97.68 45.4 98.16 ;
        RECT 46.6 97.68 95.08 98.16 ;
        RECT 25.76 103.12 26.24 103.6 ;
        RECT 91.52 103.12 92 103.6 ;
        RECT 25.76 108.56 45.4 108.8 ;
        RECT 46.6 108.56 92 108.8 ;
      LAYER met5 ;
        RECT 0 42.6 3.2 45.8 ;
        RECT 114.56 42.6 117.76 45.8 ;
        RECT 0 83.4 3.2 86.6 ;
        RECT 114.56 83.4 117.76 86.6 ;
      LAYER met4 ;
        RECT 51.22 0 51.82 0.6 ;
        RECT 80.66 0 81.26 0.6 ;
        RECT 10.74 10.88 11.34 11.48 ;
        RECT 10.74 97.32 11.34 97.92 ;
        RECT 51.22 108.2 51.82 108.8 ;
        RECT 80.66 108.2 81.26 108.8 ;
    END
  END VSS
  OBS
    LAYER met4 ;
      POLYGON 91.69 36.53 91.69 11.385 91.705 11.385 91.705 11.055 91.375 11.055 91.375 11.385 91.39 11.385 91.39 36.53 ;
      POLYGON 91.6 108.4 91.6 97.52 106.02 97.52 106.02 96.92 107.42 96.92 107.42 97.52 117.36 97.52 117.36 11.28 107.42 11.28 107.42 11.88 106.02 11.88 106.02 11.28 91.6 11.28 91.6 0.4 81.66 0.4 81.66 1 80.26 1 80.26 0.4 75.53 0.4 75.53 1.2 74.43 1.2 74.43 0.4 72.77 0.4 72.77 1.2 71.67 1.2 71.67 0.4 70.93 0.4 70.93 1.2 69.83 1.2 69.83 0.4 66.94 0.4 66.94 1 65.54 1 65.54 0.4 53.45 0.4 53.45 1.2 52.35 1.2 52.35 0.4 52.22 0.4 52.22 1 50.82 1 50.82 0.4 37.5 0.4 37.5 1 36.1 1 36.1 0.4 26.16 0.4 26.16 11.28 11.74 11.28 11.74 11.88 10.34 11.88 10.34 11.28 9.29 11.28 9.29 12.08 8.19 12.08 8.19 11.28 7.45 11.28 7.45 12.08 6.35 12.08 6.35 11.28 0.4 11.28 0.4 97.52 10.34 97.52 10.34 96.92 11.74 96.92 11.74 97.52 26.16 97.52 26.16 108.4 36.1 108.4 36.1 107.8 37.5 107.8 37.5 108.4 50.82 108.4 50.82 107.8 52.22 107.8 52.22 108.4 52.35 108.4 52.35 107.6 53.45 107.6 53.45 108.4 54.19 108.4 54.19 107.6 55.29 107.6 55.29 108.4 56.03 108.4 56.03 107.6 57.13 107.6 57.13 108.4 57.87 108.4 57.87 107.6 58.97 107.6 58.97 108.4 59.71 108.4 59.71 107.6 60.81 107.6 60.81 108.4 61.55 108.4 61.55 107.6 62.65 107.6 62.65 108.4 63.39 108.4 63.39 107.6 64.49 107.6 64.49 108.4 65.54 108.4 65.54 107.8 66.94 107.8 66.94 108.4 67.07 108.4 67.07 107.6 68.17 107.6 68.17 108.4 68.91 108.4 68.91 107.6 70.01 107.6 70.01 108.4 71.67 108.4 71.67 107.6 72.77 107.6 72.77 108.4 73.51 108.4 73.51 107.6 74.61 107.6 74.61 108.4 80.26 108.4 80.26 107.8 81.66 107.8 81.66 108.4 ;
    LAYER met2 ;
      RECT 80.82 108.615 81.1 108.985 ;
      RECT 51.38 108.615 51.66 108.985 ;
      RECT 10.9 97.735 11.18 98.105 ;
      RECT 10.9 10.695 11.18 11.065 ;
      RECT 80.82 -0.185 81.1 0.185 ;
      RECT 51.38 -0.185 51.66 0.185 ;
      POLYGON 91.72 108.52 91.72 97.64 117.48 97.64 117.48 11.16 113.28 11.16 113.28 11.645 112.58 11.645 112.58 11.16 111.9 11.16 111.9 11.645 111.2 11.645 111.2 11.16 109.14 11.16 109.14 11.645 108.44 11.645 108.44 11.16 108.22 11.16 108.22 11.645 107.52 11.645 107.52 11.16 107.3 11.16 107.3 11.645 106.6 11.645 106.6 11.16 106.38 11.16 106.38 11.645 105.68 11.645 105.68 11.16 105.46 11.16 105.46 11.645 104.76 11.645 104.76 11.16 104.54 11.16 104.54 11.645 103.84 11.645 103.84 11.16 91.72 11.16 91.72 0.28 89.82 0.28 89.82 0.765 89.12 0.765 89.12 0.28 88.9 0.28 88.9 0.765 88.2 0.765 88.2 0.28 87.98 0.28 87.98 0.765 87.28 0.765 87.28 0.28 86.6 0.28 86.6 0.765 85.9 0.765 85.9 0.28 85.68 0.28 85.68 0.765 84.98 0.765 84.98 0.28 84.76 0.28 84.76 0.765 84.06 0.765 84.06 0.28 83.84 0.28 83.84 0.765 83.14 0.765 83.14 0.28 82.92 0.28 82.92 0.765 82.22 0.765 82.22 0.28 82 0.28 82 0.765 81.3 0.765 81.3 0.28 80.62 0.28 80.62 0.765 79.92 0.765 79.92 0.28 79.7 0.28 79.7 0.765 79 0.765 79 0.28 78.78 0.28 78.78 0.765 78.08 0.765 78.08 0.28 77.4 0.28 77.4 0.765 76.7 0.765 76.7 0.28 76.48 0.28 76.48 0.765 75.78 0.765 75.78 0.28 75.56 0.28 75.56 0.765 74.86 0.765 74.86 0.28 74.64 0.28 74.64 0.765 73.94 0.765 73.94 0.28 73.72 0.28 73.72 0.765 73.02 0.765 73.02 0.28 72.8 0.28 72.8 0.765 72.1 0.765 72.1 0.28 71.42 0.28 71.42 0.765 70.72 0.765 70.72 0.28 70.5 0.28 70.5 0.765 69.8 0.765 69.8 0.28 69.58 0.28 69.58 0.765 68.88 0.765 68.88 0.28 68.2 0.28 68.2 0.765 67.5 0.765 67.5 0.28 67.28 0.28 67.28 0.765 66.58 0.765 66.58 0.28 66.36 0.28 66.36 0.765 65.66 0.765 65.66 0.28 65.44 0.28 65.44 0.765 64.74 0.765 64.74 0.28 64.52 0.28 64.52 0.765 63.82 0.765 63.82 0.28 63.6 0.28 63.6 0.765 62.9 0.765 62.9 0.28 62.68 0.28 62.68 0.765 61.98 0.765 61.98 0.28 61.76 0.28 61.76 0.765 61.06 0.765 61.06 0.28 60.84 0.28 60.84 0.765 60.14 0.765 60.14 0.28 59.92 0.28 59.92 0.765 59.22 0.765 59.22 0.28 59 0.28 59 0.765 58.3 0.765 58.3 0.28 58.08 0.28 58.08 0.765 57.38 0.765 57.38 0.28 57.16 0.28 57.16 0.765 56.46 0.765 56.46 0.28 56.24 0.28 56.24 0.765 55.54 0.765 55.54 0.28 55.32 0.28 55.32 0.765 54.62 0.765 54.62 0.28 54.4 0.28 54.4 0.765 53.7 0.765 53.7 0.28 53.48 0.28 53.48 0.765 52.78 0.765 52.78 0.28 52.56 0.28 52.56 0.765 51.86 0.765 51.86 0.28 40.6 0.28 40.6 0.765 39.9 0.765 39.9 0.28 39.68 0.28 39.68 0.765 38.98 0.765 38.98 0.28 38.76 0.28 38.76 0.765 38.06 0.765 38.06 0.28 37.84 0.28 37.84 0.765 37.14 0.765 37.14 0.28 36.92 0.28 36.92 0.765 36.22 0.765 36.22 0.28 36 0.28 36 0.765 35.3 0.765 35.3 0.28 35.08 0.28 35.08 0.765 34.38 0.765 34.38 0.28 33.24 0.28 33.24 0.765 32.54 0.765 32.54 0.28 28.64 0.28 28.64 0.765 27.94 0.765 27.94 0.28 26.04 0.28 26.04 11.16 15.76 11.16 15.76 11.645 15.06 11.645 15.06 11.16 14.84 11.16 14.84 11.645 14.14 11.645 14.14 11.16 13.92 11.16 13.92 11.645 13.22 11.645 13.22 11.16 13 11.16 13 11.645 12.3 11.645 12.3 11.16 12.08 11.16 12.08 11.645 11.38 11.645 11.38 11.16 10.7 11.16 10.7 11.645 10 11.645 10 11.16 9.32 11.16 9.32 11.645 8.62 11.645 8.62 11.16 8.4 11.16 8.4 11.645 7.7 11.645 7.7 11.16 7.48 11.16 7.48 11.645 6.78 11.645 6.78 11.16 6.56 11.16 6.56 11.645 5.86 11.645 5.86 11.16 5.64 11.16 5.64 11.645 4.94 11.645 4.94 11.16 4.72 11.16 4.72 11.645 4.02 11.645 4.02 11.16 3.34 11.16 3.34 11.645 2.64 11.645 2.64 11.16 0.28 11.16 0.28 97.64 4.02 97.64 4.02 97.155 4.72 97.155 4.72 97.64 6.78 97.64 6.78 97.155 7.48 97.155 7.48 97.64 8.16 97.64 8.16 97.155 8.86 97.155 8.86 97.64 9.08 97.64 9.08 97.155 9.78 97.155 9.78 97.64 10 97.64 10 97.155 10.7 97.155 10.7 97.64 11.38 97.64 11.38 97.155 12.08 97.155 12.08 97.64 12.3 97.64 12.3 97.155 13 97.155 13 97.64 13.22 97.64 13.22 97.155 13.92 97.155 13.92 97.64 26.04 97.64 26.04 108.52 38.06 108.52 38.06 108.035 38.76 108.035 38.76 108.52 38.98 108.52 38.98 108.035 39.68 108.035 39.68 108.52 50.48 108.52 50.48 108.035 51.18 108.035 51.18 108.52 51.86 108.52 51.86 108.035 52.56 108.035 52.56 108.52 52.78 108.52 52.78 108.035 53.48 108.035 53.48 108.52 54.16 108.52 54.16 108.035 54.86 108.035 54.86 108.52 55.08 108.52 55.08 108.035 55.78 108.035 55.78 108.52 56.46 108.52 56.46 108.035 57.16 108.035 57.16 108.52 57.38 108.52 57.38 108.035 58.08 108.035 58.08 108.52 58.3 108.52 58.3 108.035 59 108.035 59 108.52 59.22 108.52 59.22 108.035 59.92 108.035 59.92 108.52 60.14 108.52 60.14 108.035 60.84 108.035 60.84 108.52 61.06 108.52 61.06 108.035 61.76 108.035 61.76 108.52 61.98 108.52 61.98 108.035 62.68 108.035 62.68 108.52 62.9 108.52 62.9 108.035 63.6 108.035 63.6 108.52 63.82 108.52 63.82 108.035 64.52 108.035 64.52 108.52 64.74 108.52 64.74 108.035 65.44 108.035 65.44 108.52 66.12 108.52 66.12 108.035 66.82 108.035 66.82 108.52 67.04 108.52 67.04 108.035 67.74 108.035 67.74 108.52 67.96 108.52 67.96 108.035 68.66 108.035 68.66 108.52 68.88 108.52 68.88 108.035 69.58 108.035 69.58 108.52 69.8 108.52 69.8 108.035 70.5 108.035 70.5 108.52 70.72 108.52 70.72 108.035 71.42 108.035 71.42 108.52 72.1 108.52 72.1 108.035 72.8 108.035 72.8 108.52 73.48 108.52 73.48 108.035 74.18 108.035 74.18 108.52 74.4 108.52 74.4 108.035 75.1 108.035 75.1 108.52 75.32 108.52 75.32 108.035 76.02 108.035 76.02 108.52 76.24 108.52 76.24 108.035 76.94 108.035 76.94 108.52 77.16 108.52 77.16 108.035 77.86 108.035 77.86 108.52 78.08 108.52 78.08 108.035 78.78 108.035 78.78 108.52 79 108.52 79 108.035 79.7 108.035 79.7 108.52 79.92 108.52 79.92 108.035 80.62 108.035 80.62 108.52 81.3 108.52 81.3 108.035 82 108.035 82 108.52 82.22 108.52 82.22 108.035 82.92 108.035 82.92 108.52 83.14 108.52 83.14 108.035 83.84 108.035 83.84 108.52 84.06 108.52 84.06 108.035 84.76 108.035 84.76 108.52 84.98 108.52 84.98 108.035 85.68 108.035 85.68 108.52 85.9 108.52 85.9 108.035 86.6 108.035 86.6 108.52 86.82 108.52 86.82 108.035 87.52 108.035 87.52 108.52 87.74 108.52 87.74 108.035 88.44 108.035 88.44 108.52 88.66 108.52 88.66 108.035 89.36 108.035 89.36 108.52 ;
    LAYER met3 ;
      POLYGON 81.125 108.965 81.125 108.96 81.34 108.96 81.34 108.64 81.125 108.64 81.125 108.635 80.795 108.635 80.795 108.64 80.58 108.64 80.58 108.96 80.795 108.96 80.795 108.965 ;
      POLYGON 51.685 108.965 51.685 108.96 51.9 108.96 51.9 108.64 51.685 108.64 51.685 108.635 51.355 108.635 51.355 108.64 51.14 108.64 51.14 108.96 51.355 108.96 51.355 108.965 ;
      POLYGON 11.205 98.085 11.205 98.08 11.42 98.08 11.42 97.76 11.205 97.76 11.205 97.755 10.875 97.755 10.875 97.76 10.66 97.76 10.66 98.08 10.875 98.08 10.875 98.085 ;
      POLYGON 26.37 12.05 26.37 11.37 34.88 11.37 34.88 11.07 26.07 11.07 26.07 12.05 ;
      POLYGON 91.73 11.38 91.73 11.06 91.35 11.06 91.35 11.07 89.32 11.07 89.32 11.37 91.35 11.37 91.35 11.38 ;
      POLYGON 11.205 11.045 11.205 11.04 11.42 11.04 11.42 10.72 11.205 10.72 11.205 10.715 10.875 10.715 10.875 10.72 10.66 10.72 10.66 11.04 10.875 11.04 10.875 11.045 ;
      POLYGON 81.125 0.165 81.125 0.16 81.34 0.16 81.34 -0.16 81.125 -0.16 81.125 -0.165 80.795 -0.165 80.795 -0.16 80.58 -0.16 80.58 0.16 80.795 0.16 80.795 0.165 ;
      POLYGON 51.685 0.165 51.685 0.16 51.9 0.16 51.9 -0.16 51.685 -0.16 51.685 -0.165 51.355 -0.165 51.355 -0.16 51.14 -0.16 51.14 0.16 51.355 0.16 51.355 0.165 ;
      POLYGON 91.6 108.4 91.6 97.52 117.36 97.52 117.36 89.97 116.56 89.97 116.56 88.87 117.36 88.87 117.36 88.61 116.56 88.61 116.56 87.51 117.36 87.51 117.36 87.25 116.56 87.25 116.56 86.15 117.36 86.15 117.36 85.89 116.56 85.89 116.56 84.79 117.36 84.79 117.36 84.53 116.56 84.53 116.56 83.43 117.36 83.43 117.36 83.17 116.56 83.17 116.56 82.07 117.36 82.07 117.36 81.81 116.56 81.81 116.56 80.71 117.36 80.71 117.36 80.45 116.56 80.45 116.56 79.35 117.36 79.35 117.36 79.09 116.56 79.09 116.56 77.99 117.36 77.99 117.36 77.73 116.56 77.73 116.56 76.63 117.36 76.63 117.36 76.37 116.56 76.37 116.56 75.27 117.36 75.27 117.36 75.01 116.56 75.01 116.56 73.91 117.36 73.91 117.36 73.65 116.56 73.65 116.56 72.55 117.36 72.55 117.36 72.29 116.56 72.29 116.56 71.19 117.36 71.19 117.36 70.93 116.56 70.93 116.56 69.83 117.36 69.83 117.36 69.57 116.56 69.57 116.56 68.47 117.36 68.47 117.36 68.21 116.56 68.21 116.56 67.11 117.36 67.11 117.36 66.85 116.56 66.85 116.56 65.75 117.36 65.75 117.36 65.49 116.56 65.49 116.56 64.39 117.36 64.39 117.36 64.13 116.56 64.13 116.56 63.03 117.36 63.03 117.36 62.77 116.56 62.77 116.56 61.67 117.36 61.67 117.36 61.41 116.56 61.41 116.56 60.31 117.36 60.31 117.36 60.05 116.56 60.05 116.56 58.95 117.36 58.95 117.36 58.69 116.56 58.69 116.56 57.59 117.36 57.59 117.36 57.33 116.56 57.33 116.56 56.23 117.36 56.23 117.36 55.97 116.56 55.97 116.56 54.87 117.36 54.87 117.36 54.61 116.56 54.61 116.56 53.51 117.36 53.51 117.36 53.25 116.56 53.25 116.56 52.15 117.36 52.15 117.36 51.89 116.56 51.89 116.56 50.79 117.36 50.79 117.36 50.53 116.56 50.53 116.56 49.43 117.36 49.43 117.36 49.17 116.56 49.17 116.56 48.07 117.36 48.07 117.36 47.81 116.56 47.81 116.56 46.71 117.36 46.71 117.36 46.45 116.56 46.45 116.56 45.35 117.36 45.35 117.36 45.09 116.56 45.09 116.56 43.99 117.36 43.99 117.36 43.73 116.56 43.73 116.56 42.63 117.36 42.63 117.36 42.37 116.56 42.37 116.56 41.27 117.36 41.27 117.36 39.65 116.56 39.65 116.56 38.55 117.36 38.55 117.36 38.29 116.56 38.29 116.56 37.19 117.36 37.19 117.36 36.93 116.56 36.93 116.56 35.83 117.36 35.83 117.36 35.57 116.56 35.57 116.56 34.47 117.36 34.47 117.36 34.21 116.56 34.21 116.56 33.11 117.36 33.11 117.36 32.85 116.56 32.85 116.56 31.75 117.36 31.75 117.36 31.49 116.56 31.49 116.56 30.39 117.36 30.39 117.36 30.13 116.56 30.13 116.56 29.03 117.36 29.03 117.36 28.77 116.56 28.77 116.56 27.67 117.36 27.67 117.36 27.41 116.56 27.41 116.56 26.31 117.36 26.31 117.36 26.05 116.56 26.05 116.56 24.95 117.36 24.95 117.36 24.69 116.56 24.69 116.56 23.59 117.36 23.59 117.36 23.33 116.56 23.33 116.56 22.23 117.36 22.23 117.36 16.53 116.56 16.53 116.56 15.43 117.36 15.43 117.36 15.17 116.56 15.17 116.56 14.07 117.36 14.07 117.36 11.28 91.6 11.28 91.6 0.4 26.16 0.4 26.16 11.28 0.4 11.28 0.4 14.07 1.2 14.07 1.2 15.17 0.4 15.17 0.4 15.43 1.2 15.43 1.2 16.53 0.4 16.53 0.4 16.79 1.2 16.79 1.2 17.89 0.4 17.89 0.4 22.23 1.2 22.23 1.2 23.33 0.4 23.33 0.4 23.59 1.2 23.59 1.2 24.69 0.4 24.69 0.4 24.95 1.2 24.95 1.2 26.05 0.4 26.05 0.4 26.31 1.2 26.31 1.2 27.41 0.4 27.41 0.4 27.67 1.2 27.67 1.2 28.77 0.4 28.77 0.4 29.03 1.2 29.03 1.2 30.13 0.4 30.13 0.4 30.39 1.2 30.39 1.2 31.49 0.4 31.49 0.4 31.75 1.2 31.75 1.2 32.85 0.4 32.85 0.4 33.11 1.2 33.11 1.2 34.21 0.4 34.21 0.4 34.47 1.2 34.47 1.2 35.57 0.4 35.57 0.4 35.83 1.2 35.83 1.2 36.93 0.4 36.93 0.4 37.19 1.2 37.19 1.2 38.29 0.4 38.29 0.4 38.55 1.2 38.55 1.2 39.65 0.4 39.65 0.4 39.91 1.2 39.91 1.2 41.01 0.4 41.01 0.4 41.27 1.2 41.27 1.2 42.37 0.4 42.37 0.4 42.63 1.2 42.63 1.2 43.73 0.4 43.73 0.4 43.99 1.2 43.99 1.2 45.09 0.4 45.09 0.4 45.35 1.2 45.35 1.2 46.45 0.4 46.45 0.4 46.71 1.2 46.71 1.2 47.81 0.4 47.81 0.4 48.07 1.2 48.07 1.2 49.17 0.4 49.17 0.4 49.43 1.2 49.43 1.2 50.53 0.4 50.53 0.4 50.79 1.2 50.79 1.2 51.89 0.4 51.89 0.4 52.15 1.2 52.15 1.2 53.25 0.4 53.25 0.4 53.51 1.2 53.51 1.2 54.61 0.4 54.61 0.4 54.87 1.2 54.87 1.2 55.97 0.4 55.97 0.4 56.23 1.2 56.23 1.2 57.33 0.4 57.33 0.4 57.59 1.2 57.59 1.2 58.69 0.4 58.69 0.4 58.95 1.2 58.95 1.2 60.05 0.4 60.05 0.4 60.31 1.2 60.31 1.2 61.41 0.4 61.41 0.4 61.67 1.2 61.67 1.2 62.77 0.4 62.77 0.4 63.03 1.2 63.03 1.2 64.13 0.4 64.13 0.4 64.39 1.2 64.39 1.2 65.49 0.4 65.49 0.4 66.43 1.2 66.43 1.2 67.53 0.4 67.53 0.4 67.79 1.2 67.79 1.2 68.89 0.4 68.89 0.4 69.15 1.2 69.15 1.2 70.25 0.4 70.25 0.4 70.51 1.2 70.51 1.2 71.61 0.4 71.61 0.4 71.87 1.2 71.87 1.2 72.97 0.4 72.97 0.4 73.23 1.2 73.23 1.2 74.33 0.4 74.33 0.4 74.59 1.2 74.59 1.2 75.69 0.4 75.69 0.4 75.95 1.2 75.95 1.2 77.05 0.4 77.05 0.4 77.31 1.2 77.31 1.2 78.41 0.4 78.41 0.4 78.67 1.2 78.67 1.2 79.77 0.4 79.77 0.4 80.03 1.2 80.03 1.2 81.13 0.4 81.13 0.4 81.39 1.2 81.39 1.2 82.49 0.4 82.49 0.4 83.43 1.2 83.43 1.2 84.53 0.4 84.53 0.4 84.79 1.2 84.79 1.2 85.89 0.4 85.89 0.4 86.15 1.2 86.15 1.2 87.25 0.4 87.25 0.4 87.51 1.2 87.51 1.2 88.61 0.4 88.61 0.4 97.52 26.16 97.52 26.16 108.4 ;
    LAYER met5 ;
      POLYGON 90.4 107.2 90.4 96.32 116.16 96.32 116.16 88.2 112.96 88.2 112.96 81.8 116.16 81.8 116.16 67.8 112.96 67.8 112.96 61.4 116.16 61.4 116.16 47.4 112.96 47.4 112.96 41 116.16 41 116.16 27 112.96 27 112.96 20.6 116.16 20.6 116.16 12.48 90.4 12.48 90.4 1.6 27.36 1.6 27.36 12.48 1.6 12.48 1.6 20.6 4.8 20.6 4.8 27 1.6 27 1.6 41 4.8 41 4.8 47.4 1.6 47.4 1.6 61.4 4.8 61.4 4.8 67.8 1.6 67.8 1.6 81.8 4.8 81.8 4.8 88.2 1.6 88.2 1.6 96.32 27.36 96.32 27.36 107.2 ;
    LAYER met1 ;
      RECT 45.68 108.56 46.32 109.04 ;
      POLYGON 90.92 108.36 90.92 107.2 90.78 107.2 90.78 108.22 68.38 108.22 68.38 106.86 68.24 106.86 68.24 108.36 ;
      POLYGON 39.95 98.56 39.95 98.5 40.545 98.5 40.545 98.545 40.835 98.545 40.835 98.315 40.545 98.315 40.545 98.36 39.95 98.36 39.95 98.3 39.63 98.3 39.63 98.56 ;
      POLYGON 75.83 97.54 75.83 97.28 75.51 97.28 75.51 97.34 74.895 97.34 74.895 97.295 74.605 97.295 74.605 97.525 74.895 97.525 74.895 97.48 75.51 97.48 75.51 97.54 ;
      POLYGON 71.69 97.54 71.69 97.48 72.305 97.48 72.305 97.525 72.595 97.525 72.595 97.295 72.305 97.295 72.305 97.34 71.69 97.34 71.69 97.28 71.37 97.28 71.37 97.54 ;
      POLYGON 62.03 97.54 62.03 97.28 61.71 97.28 61.71 97.34 27.07 97.34 27.07 97.28 26.75 97.28 26.75 97.54 27.07 97.54 27.07 97.48 61.71 97.48 61.71 97.54 ;
      POLYGON 26.15 97.54 26.15 97.28 25.83 97.28 25.83 97.34 20.54 97.34 20.54 95.98 20.4 95.98 20.4 97.48 25.83 97.48 25.83 97.54 ;
      POLYGON 12.26 12.48 12.26 11.46 30.43 11.46 30.43 11.52 30.52 11.52 30.52 11.8 30.66 11.8 30.66 11.52 30.75 11.52 30.75 11.26 30.43 11.26 30.43 11.32 12.12 11.32 12.12 12.48 ;
      POLYGON 53.66 11.8 53.66 11.46 64.47 11.46 64.47 11.52 64.79 11.52 64.79 11.26 64.47 11.26 64.47 11.32 53.52 11.32 53.52 11.8 ;
      POLYGON 79.05 11.52 79.05 11.26 78.73 11.26 78.73 11.32 76.275 11.32 76.275 11.275 75.985 11.275 75.985 11.32 75.37 11.32 75.37 11.26 75.05 11.26 75.05 11.52 75.37 11.52 75.37 11.46 75.985 11.46 75.985 11.505 76.275 11.505 76.275 11.46 78.73 11.46 78.73 11.52 ;
      POLYGON 52.37 11.52 52.37 11.26 52.05 11.26 52.05 11.32 51.435 11.32 51.435 11.275 51.145 11.275 51.145 11.505 51.435 11.505 51.435 11.46 52.05 11.46 52.05 11.52 ;
      RECT 50.67 11.26 50.99 11.52 ;
      POLYGON 40.41 11.52 40.41 11.26 40.09 11.26 40.09 11.32 34.875 11.32 34.875 11.275 34.585 11.275 34.585 11.505 34.875 11.505 34.875 11.46 40.09 11.46 40.09 11.52 ;
      POLYGON 33.97 11.52 33.97 11.26 33.65 11.26 33.65 11.32 32.575 11.32 32.575 11.275 32.285 11.275 32.285 11.505 32.575 11.505 32.575 11.46 33.65 11.46 33.65 11.52 ;
      POLYGON 46.39 10.5 46.39 10.44 47.005 10.44 47.005 10.485 47.295 10.485 47.295 10.255 47.005 10.255 47.005 10.3 46.39 10.3 46.39 10.24 46.07 10.24 46.07 10.3 44.135 10.3 44.135 10.255 44.09 10.255 44.09 10.24 43.77 10.24 43.77 10.5 44.09 10.5 44.09 10.485 44.135 10.485 44.135 10.44 46.07 10.44 46.07 10.5 ;
      POLYGON 37.65 10.5 37.65 10.44 37.805 10.44 37.805 10.485 38.095 10.485 38.095 10.255 37.805 10.255 37.805 10.3 37.65 10.3 37.65 10.24 37.33 10.24 37.33 10.5 ;
      POLYGON 34.89 10.5 34.89 10.44 35.965 10.44 35.965 10.485 36.255 10.485 36.255 10.255 35.965 10.255 35.965 10.3 34.89 10.3 34.89 10.24 34.57 10.24 34.57 10.5 ;
      RECT 33.65 10.24 33.97 10.5 ;
      POLYGON 42.235 10.485 42.235 10.255 41.945 10.255 41.945 10.3 39.995 10.3 39.995 10.255 39.705 10.255 39.705 10.485 39.995 10.485 39.995 10.44 41.945 10.44 41.945 10.485 ;
      RECT 45.68 -0.24 46.32 0.24 ;
      POLYGON 46.32 108.52 46.32 108.28 91.72 108.28 91.72 106.6 91.24 106.6 91.24 105.56 91.72 105.56 91.72 103.88 91.24 103.88 91.24 102.84 91.72 102.84 91.72 101.16 91.24 101.16 91.24 100.12 91.72 100.12 91.72 98.44 46.32 98.44 46.32 97.4 95.36 97.4 95.36 97.64 96 97.64 96 97.4 117.48 97.4 117.48 95.72 117 95.72 117 94.68 117.48 94.68 117.48 93 117 93 117 91.96 117.48 91.96 117.48 90.28 117 90.28 117 89.24 117.48 89.24 117.48 87.56 117 87.56 117 86.52 117.48 86.52 117.48 84.84 117 84.84 117 83.8 117.48 83.8 117.48 82.12 117 82.12 117 81.08 117.48 81.08 117.48 79.4 117 79.4 117 78.36 117.48 78.36 117.48 76.68 117 76.68 117 75.64 117.48 75.64 117.48 73.96 117 73.96 117 72.92 117.48 72.92 117.48 71.24 117 71.24 117 70.2 117.48 70.2 117.48 68.52 117 68.52 117 67.48 117.48 67.48 117.48 65.8 117 65.8 117 64.76 117.48 64.76 117.48 63.08 117 63.08 117 62.04 117.48 62.04 117.48 60.36 117 60.36 117 59.32 117.48 59.32 117.48 57.64 117 57.64 117 56.6 117.48 56.6 117.48 54.92 117 54.92 117 53.88 117.48 53.88 117.48 52.2 117 52.2 117 51.16 117.48 51.16 117.48 49.48 117 49.48 117 48.44 117.48 48.44 117.48 46.76 117 46.76 117 45.72 117.48 45.72 117.48 44.04 117 44.04 117 43 117.48 43 117.48 41.32 117 41.32 117 40.28 117.48 40.28 117.48 38.6 117 38.6 117 37.56 117.48 37.56 117.48 35.88 117 35.88 117 34.84 117.48 34.84 117.48 33.16 117 33.16 117 32.12 117.48 32.12 117.48 30.44 117 30.44 117 29.4 117.48 29.4 117.48 27.72 117 27.72 117 26.68 117.48 26.68 117.48 25 117 25 117 23.96 117.48 23.96 117.48 22.28 117 22.28 117 21.24 117.48 21.24 117.48 19.56 117 19.56 117 18.52 117.48 18.52 117.48 16.84 117 16.84 117 15.8 117.48 15.8 117.48 14.12 117 14.12 117 13.08 117.48 13.08 117.48 11.4 96 11.4 96 11.16 95.36 11.16 95.36 11.4 46.32 11.4 46.32 10.36 91.72 10.36 91.72 8.68 91.24 8.68 91.24 7.64 91.72 7.64 91.72 5.96 91.24 5.96 91.24 4.92 91.72 4.92 91.72 3.24 91.24 3.24 91.24 2.2 91.72 2.2 91.72 0.52 46.32 0.52 46.32 0.28 45.68 0.28 45.68 0.52 26.04 0.52 26.04 2.2 26.52 2.2 26.52 3.24 26.04 3.24 26.04 4.92 26.52 4.92 26.52 5.96 26.04 5.96 26.04 7.64 26.52 7.64 26.52 8.68 26.04 8.68 26.04 10.36 45.68 10.36 45.68 11.4 0.28 11.4 0.28 13.08 0.76 13.08 0.76 14.12 0.28 14.12 0.28 15.8 0.76 15.8 0.76 16.84 0.28 16.84 0.28 18.52 0.76 18.52 0.76 19.56 0.28 19.56 0.28 21.24 0.76 21.24 0.76 22.28 0.28 22.28 0.28 23.96 0.76 23.96 0.76 25 0.28 25 0.28 26.68 0.76 26.68 0.76 27.72 0.28 27.72 0.28 29.4 0.76 29.4 0.76 30.44 0.28 30.44 0.28 32.12 0.76 32.12 0.76 33.16 0.28 33.16 0.28 34.84 0.76 34.84 0.76 35.88 0.28 35.88 0.28 37.56 0.76 37.56 0.76 38.6 0.28 38.6 0.28 40.28 0.76 40.28 0.76 41.32 0.28 41.32 0.28 43 0.76 43 0.76 44.04 0.28 44.04 0.28 45.72 0.76 45.72 0.76 46.76 0.28 46.76 0.28 48.44 0.76 48.44 0.76 49.48 0.28 49.48 0.28 51.16 0.76 51.16 0.76 52.2 0.28 52.2 0.28 53.88 0.76 53.88 0.76 54.92 0.28 54.92 0.28 56.6 0.76 56.6 0.76 57.64 0.28 57.64 0.28 59.32 0.76 59.32 0.76 60.36 0.28 60.36 0.28 62.04 0.76 62.04 0.76 63.08 0.28 63.08 0.28 64.76 0.76 64.76 0.76 65.8 0.28 65.8 0.28 67.48 0.76 67.48 0.76 68.52 0.28 68.52 0.28 70.2 0.76 70.2 0.76 71.24 0.28 71.24 0.28 72.92 0.76 72.92 0.76 73.96 0.28 73.96 0.28 75.64 0.76 75.64 0.76 76.68 0.28 76.68 0.28 78.36 0.76 78.36 0.76 79.4 0.28 79.4 0.28 81.08 0.76 81.08 0.76 82.12 0.28 82.12 0.28 83.8 0.76 83.8 0.76 84.84 0.28 84.84 0.28 86.52 0.76 86.52 0.76 87.56 0.28 87.56 0.28 89.24 0.76 89.24 0.76 90.28 0.28 90.28 0.28 91.96 0.76 91.96 0.76 93 0.28 93 0.28 94.68 0.76 94.68 0.76 95.72 0.28 95.72 0.28 97.4 45.68 97.4 45.68 98.44 26.04 98.44 26.04 100.12 26.52 100.12 26.52 101.16 26.04 101.16 26.04 102.84 26.52 102.84 26.52 103.88 26.04 103.88 26.04 105.56 26.52 105.56 26.52 106.6 26.04 106.6 26.04 108.28 45.68 108.28 45.68 108.52 ;
    LAYER li1 ;
      RECT 25.76 108.715 92 108.885 ;
      RECT 88.32 105.995 92 106.165 ;
      RECT 25.76 105.995 29.44 106.165 ;
      RECT 91.54 103.275 92 103.445 ;
      RECT 25.76 103.275 29.44 103.445 ;
      RECT 91.08 100.555 92 100.725 ;
      RECT 25.76 100.555 29.44 100.725 ;
      RECT 89.24 97.835 117.76 98.005 ;
      RECT 0 97.835 29.44 98.005 ;
      RECT 116.84 95.115 117.76 95.285 ;
      RECT 0 95.115 3.68 95.285 ;
      RECT 116.84 92.395 117.76 92.565 ;
      RECT 0 92.395 3.68 92.565 ;
      RECT 116.84 89.675 117.76 89.845 ;
      RECT 0 89.675 3.68 89.845 ;
      RECT 116.84 86.955 117.76 87.125 ;
      RECT 0 86.955 3.68 87.125 ;
      RECT 116.84 84.235 117.76 84.405 ;
      RECT 0 84.235 3.68 84.405 ;
      RECT 116.84 81.515 117.76 81.685 ;
      RECT 0 81.515 3.68 81.685 ;
      RECT 114.08 78.795 117.76 78.965 ;
      RECT 0 78.795 1.84 78.965 ;
      RECT 114.08 76.075 117.76 76.245 ;
      RECT 0 76.075 3.68 76.245 ;
      RECT 116.84 73.355 117.76 73.525 ;
      RECT 0 73.355 3.68 73.525 ;
      RECT 116.84 70.635 117.76 70.805 ;
      RECT 0 70.635 1.84 70.805 ;
      RECT 116.84 67.915 117.76 68.085 ;
      RECT 0 67.915 1.84 68.085 ;
      RECT 116.84 65.195 117.76 65.365 ;
      RECT 0 65.195 3.68 65.365 ;
      RECT 116.84 62.475 117.76 62.645 ;
      RECT 0 62.475 3.68 62.645 ;
      RECT 116.84 59.755 117.76 59.925 ;
      RECT 0 59.755 3.68 59.925 ;
      RECT 116.84 57.035 117.76 57.205 ;
      RECT 0 57.035 3.68 57.205 ;
      RECT 114.08 54.315 117.76 54.485 ;
      RECT 0 54.315 3.68 54.485 ;
      RECT 114.08 51.595 117.76 51.765 ;
      RECT 0 51.595 3.68 51.765 ;
      RECT 116.84 48.875 117.76 49.045 ;
      RECT 0 48.875 1.84 49.045 ;
      RECT 116.84 46.155 117.76 46.325 ;
      RECT 0 46.155 1.84 46.325 ;
      RECT 116.84 43.435 117.76 43.605 ;
      RECT 0 43.435 3.68 43.605 ;
      RECT 114.08 40.715 117.76 40.885 ;
      RECT 0 40.715 3.68 40.885 ;
      RECT 114.08 37.995 117.76 38.165 ;
      RECT 0 37.995 3.68 38.165 ;
      RECT 116.84 35.275 117.76 35.445 ;
      RECT 0 35.275 3.68 35.445 ;
      RECT 114.08 32.555 117.76 32.725 ;
      RECT 0 32.555 1.84 32.725 ;
      RECT 114.08 29.835 117.76 30.005 ;
      RECT 0 29.835 1.84 30.005 ;
      RECT 116.84 27.115 117.76 27.285 ;
      RECT 0 27.115 1.84 27.285 ;
      RECT 116.84 24.395 117.76 24.565 ;
      RECT 0 24.395 3.68 24.565 ;
      RECT 114.08 21.675 117.76 21.845 ;
      RECT 0 21.675 3.68 21.845 ;
      RECT 114.08 18.955 117.76 19.125 ;
      RECT 0 18.955 3.68 19.125 ;
      RECT 117.3 16.235 117.76 16.405 ;
      RECT 0 16.235 3.68 16.405 ;
      RECT 117.3 13.515 117.76 13.685 ;
      RECT 0 13.515 3.68 13.685 ;
      RECT 88.78 10.795 117.76 10.965 ;
      RECT 0 10.795 29.44 10.965 ;
      RECT 90.16 8.075 92 8.245 ;
      RECT 25.76 8.075 29.44 8.245 ;
      RECT 91.54 5.355 92 5.525 ;
      RECT 25.76 5.355 29.44 5.525 ;
      RECT 88.32 2.635 92 2.805 ;
      RECT 25.76 2.635 29.44 2.805 ;
      RECT 25.76 -0.085 92 0.085 ;
      POLYGON 91.83 108.63 91.83 97.75 117.59 97.75 117.59 11.05 91.83 11.05 91.83 0.17 25.93 0.17 25.93 11.05 0.17 11.05 0.17 97.75 25.93 97.75 25.93 108.63 ;
    LAYER mcon ;
      RECT 40.605 98.345 40.775 98.515 ;
      RECT 74.665 97.325 74.835 97.495 ;
      RECT 72.365 97.325 72.535 97.495 ;
      RECT 76.045 11.305 76.215 11.475 ;
      RECT 51.205 11.305 51.375 11.475 ;
      RECT 50.755 11.305 50.925 11.475 ;
      RECT 34.645 11.305 34.815 11.475 ;
      RECT 32.345 11.305 32.515 11.475 ;
      RECT 47.065 10.285 47.235 10.455 ;
      RECT 43.905 10.285 44.075 10.455 ;
      RECT 42.005 10.285 42.175 10.455 ;
      RECT 39.765 10.285 39.935 10.455 ;
      RECT 37.865 10.285 38.035 10.455 ;
      RECT 36.025 10.285 36.195 10.455 ;
      RECT 33.725 10.285 33.895 10.455 ;
    LAYER via ;
      RECT 80.885 108.725 81.035 108.875 ;
      RECT 51.445 108.725 51.595 108.875 ;
      RECT 39.715 98.355 39.865 98.505 ;
      RECT 80.885 97.845 81.035 97.995 ;
      RECT 51.445 97.845 51.595 97.995 ;
      RECT 10.965 97.845 11.115 97.995 ;
      RECT 75.595 97.335 75.745 97.485 ;
      RECT 71.455 97.335 71.605 97.485 ;
      RECT 61.795 97.335 61.945 97.485 ;
      RECT 26.835 97.335 26.985 97.485 ;
      RECT 25.915 97.335 26.065 97.485 ;
      RECT 78.815 11.315 78.965 11.465 ;
      RECT 75.135 11.315 75.285 11.465 ;
      RECT 64.555 11.315 64.705 11.465 ;
      RECT 52.135 11.315 52.285 11.465 ;
      RECT 50.755 11.315 50.905 11.465 ;
      RECT 40.175 11.315 40.325 11.465 ;
      RECT 33.735 11.315 33.885 11.465 ;
      RECT 30.515 11.315 30.665 11.465 ;
      RECT 80.885 10.805 81.035 10.955 ;
      RECT 51.445 10.805 51.595 10.955 ;
      RECT 10.965 10.805 11.115 10.955 ;
      RECT 43.855 10.295 44.005 10.445 ;
      RECT 37.415 10.295 37.565 10.445 ;
      RECT 34.655 10.295 34.805 10.445 ;
      RECT 33.735 10.295 33.885 10.445 ;
      RECT 80.885 -0.075 81.035 0.075 ;
      RECT 51.445 -0.075 51.595 0.075 ;
    LAYER via2 ;
      RECT 80.86 108.7 81.06 108.9 ;
      RECT 51.42 108.7 51.62 108.9 ;
      RECT 10.94 97.82 11.14 98.02 ;
      RECT 1.05 72.32 1.25 72.52 ;
      RECT 116.51 44.44 116.71 44.64 ;
      RECT 10.94 10.78 11.14 10.98 ;
      RECT 80.86 -0.1 81.06 0.1 ;
      RECT 51.42 -0.1 51.62 0.1 ;
    LAYER via3 ;
      RECT 80.86 108.7 81.06 108.9 ;
      RECT 51.42 108.7 51.62 108.9 ;
      RECT 10.94 97.82 11.14 98.02 ;
      RECT 91.44 11.12 91.64 11.32 ;
      RECT 10.94 10.78 11.14 10.98 ;
      RECT 80.86 -0.1 81.06 0.1 ;
      RECT 51.42 -0.1 51.62 0.1 ;
    LAYER OVERLAP ;
      POLYGON 25.76 0 25.76 10.88 0 10.88 0 97.92 25.76 97.92 25.76 108.8 92 108.8 92 97.92 117.76 97.92 117.76 10.88 92 10.88 92 0 ;
  END
END sb_1__1_

END LIBRARY
