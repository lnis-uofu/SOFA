VERSION 5.7 ;
BUSBITCHARS "[]" ;

UNITS
  DATABASE MICRONS 1000 ;
END UNITS

MANUFACTURINGGRID 0.005 ;

LAYER li1
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.46 ;
  WIDTH 0.17 ;
END li1

LAYER mcon
  TYPE CUT ;
END mcon

LAYER met1
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.34 ;
  WIDTH 0.14 ;
END met1

LAYER via
  TYPE CUT ;
END via

LAYER met2
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.46 ;
  WIDTH 0.14 ;
END met2

LAYER via2
  TYPE CUT ;
END via2

LAYER met3
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.68 ;
  WIDTH 0.3 ;
END met3

LAYER via3
  TYPE CUT ;
END via3

LAYER met4
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.92 ;
  WIDTH 0.3 ;
END met4

LAYER via4
  TYPE CUT ;
END via4

LAYER met5
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 3.4 ;
  WIDTH 1.6 ;
END met5

LAYER nwell
  TYPE MASTERSLICE ;
END nwell

LAYER pwell
  TYPE MASTERSLICE ;
END pwell

LAYER OVERLAP
  TYPE OVERLAP ;
END OVERLAP

VIA L1M1_PR
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.145 -0.115 0.145 0.115 ;
END L1M1_PR

VIA L1M1_PR_R
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.115 -0.145 0.115 0.145 ;
END L1M1_PR_R

VIA L1M1_PR_M
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.115 -0.145 0.115 0.145 ;
END L1M1_PR_M

VIA L1M1_PR_MR
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.145 -0.115 0.145 0.115 ;
END L1M1_PR_MR

VIA L1M1_PR_C
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.145 -0.145 0.145 0.145 ;
END L1M1_PR_C

VIA M1M2_PR
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR

VIA M1M2_PR_Enc
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_Enc

VIA M1M2_PR_R
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_R

VIA M1M2_PR_R_Enc
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR_R_Enc

VIA M1M2_PR_M
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_M

VIA M1M2_PR_M_Enc
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR_M_Enc

VIA M1M2_PR_MR
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR_MR

VIA M1M2_PR_MR_Enc
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_MR_Enc

VIA M1M2_PR_C
  LAYER met1 ;
    RECT -0.16 -0.16 0.16 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.16 0.16 0.16 ;
END M1M2_PR_C

VIA M2M3_PR
  LAYER met2 ;
    RECT -0.14 -0.185 0.14 0.185 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR

VIA M2M3_PR_R
  LAYER met2 ;
    RECT -0.185 -0.14 0.185 0.14 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_R

VIA M2M3_PR_M
  LAYER met2 ;
    RECT -0.14 -0.185 0.14 0.185 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_M

VIA M2M3_PR_MR
  LAYER met2 ;
    RECT -0.185 -0.14 0.185 0.14 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_MR

VIA M2M3_PR_C
  LAYER met2 ;
    RECT -0.185 -0.185 0.185 0.185 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_C

VIA M3M4_PR
  LAYER met3 ;
    RECT -0.19 -0.16 0.19 0.16 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR

VIA M3M4_PR_R
  LAYER met3 ;
    RECT -0.16 -0.19 0.16 0.19 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_R

VIA M3M4_PR_M
  LAYER met3 ;
    RECT -0.19 -0.16 0.19 0.16 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_M

VIA M3M4_PR_MR
  LAYER met3 ;
    RECT -0.16 -0.19 0.16 0.19 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_MR

VIA M3M4_PR_C
  LAYER met3 ;
    RECT -0.19 -0.19 0.19 0.19 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_C

VIA M4M5_PR
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR

VIA M4M5_PR_R
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_R

VIA M4M5_PR_M
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_M

VIA M4M5_PR_MR
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_MR

VIA M4M5_PR_C
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_C

SITE unit
  CLASS CORE ;
  SYMMETRY Y ;
  SIZE 0.46 BY 2.72 ;
END unit

SITE unithddbl
  CLASS CORE ;
  SIZE 0.46 BY 5.44 ;
END unithddbl

MACRO cby_1__1_
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  SIZE 66.24 BY 76.16 ;
  SYMMETRY X Y ;
  PIN prog_clk[0]
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER met3 ;
        RECT 0 3.25 1.38 3.55 ;
    END
  END prog_clk[0]
  PIN chany_bottom_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.21 0 31.35 1.36 ;
    END
  END chany_bottom_in[0]
  PIN chany_bottom_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.05 0 33.19 1.36 ;
    END
  END chany_bottom_in[1]
  PIN chany_bottom_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.07 0 27.21 1.36 ;
    END
  END chany_bottom_in[2]
  PIN chany_bottom_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.47 0 45.61 1.36 ;
    END
  END chany_bottom_in[3]
  PIN chany_bottom_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.87 0 41.01 1.36 ;
    END
  END chany_bottom_in[4]
  PIN chany_bottom_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.61 0 49.75 1.36 ;
    END
  END chany_bottom_in[5]
  PIN chany_bottom_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.13 0 32.27 1.36 ;
    END
  END chany_bottom_in[6]
  PIN chany_bottom_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.71 0 42.85 1.36 ;
    END
  END chany_bottom_in[7]
  PIN chany_bottom_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.77 0 24.91 1.36 ;
    END
  END chany_bottom_in[8]
  PIN chany_bottom_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.79 0 41.93 1.36 ;
    END
  END chany_bottom_in[9]
  PIN chany_bottom_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.83 0 29.97 1.36 ;
    END
  END chany_bottom_in[10]
  PIN chany_bottom_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.29 0 53.43 1.36 ;
    END
  END chany_bottom_in[11]
  PIN chany_bottom_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.05 0 56.19 1.36 ;
    END
  END chany_bottom_in[12]
  PIN chany_bottom_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.09 0 44.23 1.36 ;
    END
  END chany_bottom_in[13]
  PIN chany_bottom_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.47 0 22.61 1.36 ;
    END
  END chany_bottom_in[14]
  PIN chany_bottom_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.39 0 46.53 1.36 ;
    END
  END chany_bottom_in[15]
  PIN chany_bottom_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.85 0 23.99 1.36 ;
    END
  END chany_bottom_in[16]
  PIN chany_bottom_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.23 0 48.37 1.36 ;
    END
  END chany_bottom_in[17]
  PIN chany_bottom_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.99 0 28.13 1.36 ;
    END
  END chany_bottom_in[18]
  PIN chany_bottom_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.27 0 59.41 1.36 ;
    END
  END chany_bottom_in[19]
  PIN chany_top_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.75 74.8 53.89 76.16 ;
    END
  END chany_top_in[0]
  PIN chany_top_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.73 74.8 36.87 76.16 ;
    END
  END chany_top_in[1]
  PIN chany_top_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.45 74.8 28.59 76.16 ;
    END
  END chany_top_in[2]
  PIN chany_top_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.01 74.8 45.15 76.16 ;
    END
  END chany_top_in[3]
  PIN chany_top_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.53 74.8 27.67 76.16 ;
    END
  END chany_top_in[4]
  PIN chany_top_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.91 74.8 52.05 76.16 ;
    END
  END chany_top_in[5]
  PIN chany_top_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.11 74.8 15.25 76.16 ;
    END
  END chany_top_in[6]
  PIN chany_top_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.39 74.8 46.53 76.16 ;
    END
  END chany_top_in[7]
  PIN chany_top_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.87 74.8 41.01 76.16 ;
    END
  END chany_top_in[8]
  PIN chany_top_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.31 74.8 47.45 76.16 ;
    END
  END chany_top_in[9]
  PIN chany_top_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.77 74.8 24.91 76.16 ;
    END
  END chany_top_in[10]
  PIN chany_top_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.23 74.8 48.37 76.16 ;
    END
  END chany_top_in[11]
  PIN chany_top_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.09 74.8 21.23 76.16 ;
    END
  END chany_top_in[12]
  PIN chany_top_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.15 74.8 49.29 76.16 ;
    END
  END chany_top_in[13]
  PIN chany_top_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.85 74.8 23.99 76.16 ;
    END
  END chany_top_in[14]
  PIN chany_top_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.49 74.8 62.63 76.16 ;
    END
  END chany_top_in[15]
  PIN chany_top_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.93 74.8 23.07 76.16 ;
    END
  END chany_top_in[16]
  PIN chany_top_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.07 74.8 50.21 76.16 ;
    END
  END chany_top_in[17]
  PIN chany_top_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.61 74.8 26.75 76.16 ;
    END
  END chany_top_in[18]
  PIN chany_top_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.99 74.8 51.13 76.16 ;
    END
  END chany_top_in[19]
  PIN ccff_head[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 58.33 1.38 58.63 ;
    END
  END ccff_head[0]
  PIN chany_bottom_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.21 0 54.35 1.36 ;
    END
  END chany_bottom_out[0]
  PIN chany_bottom_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.89 0 35.03 1.36 ;
    END
  END chany_bottom_out[1]
  PIN chany_bottom_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.97 0 34.11 1.36 ;
    END
  END chany_bottom_out[2]
  PIN chany_bottom_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.45 0 51.59 1.36 ;
    END
  END chany_bottom_out[3]
  PIN chany_bottom_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 42.17 0 42.47 1.36 ;
    END
  END chany_bottom_out[4]
  PIN chany_bottom_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.91 0 29.05 1.36 ;
    END
  END chany_bottom_out[5]
  PIN chany_bottom_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.89 0 58.03 1.36 ;
    END
  END chany_bottom_out[6]
  PIN chany_bottom_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.31 0 47.45 1.36 ;
    END
  END chany_bottom_out[7]
  PIN chany_bottom_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.65 0 37.79 1.36 ;
    END
  END chany_bottom_out[8]
  PIN chany_bottom_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.55 0 21.69 1.36 ;
    END
  END chany_bottom_out[9]
  PIN chany_bottom_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 37.57 0 37.87 1.36 ;
    END
  END chany_bottom_out[10]
  PIN chany_bottom_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.37 0 52.51 1.36 ;
    END
  END chany_bottom_out[11]
  PIN chany_bottom_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.97 0 57.11 1.36 ;
    END
  END chany_bottom_out[12]
  PIN chany_bottom_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.53 0 50.67 1.36 ;
    END
  END chany_bottom_out[13]
  PIN chany_bottom_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.81 0 35.95 1.36 ;
    END
  END chany_bottom_out[14]
  PIN chany_bottom_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.63 0 20.77 1.36 ;
    END
  END chany_bottom_out[15]
  PIN chany_bottom_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 44.01 0 44.31 1.36 ;
    END
  END chany_bottom_out[16]
  PIN chany_bottom_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.95 0 40.09 1.36 ;
    END
  END chany_bottom_out[17]
  PIN chany_bottom_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.73 0 36.87 1.36 ;
    END
  END chany_bottom_out[18]
  PIN chany_bottom_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.57 0 38.71 1.36 ;
    END
  END chany_bottom_out[19]
  PIN chany_top_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.13 74.8 32.27 76.16 ;
    END
  END chany_top_out[0]
  PIN chany_top_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.49 74.8 39.63 76.16 ;
    END
  END chany_top_out[1]
  PIN chany_top_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.57 74.8 38.71 76.16 ;
    END
  END chany_top_out[2]
  PIN chany_top_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.09 74.8 44.23 76.16 ;
    END
  END chany_top_out[3]
  PIN chany_top_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.29 74.8 30.43 76.16 ;
    END
  END chany_top_out[4]
  PIN chany_top_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.79 74.8 41.93 76.16 ;
    END
  END chany_top_out[5]
  PIN chany_top_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.81 74.8 58.95 76.16 ;
    END
  END chany_top_out[6]
  PIN chany_top_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.97 74.8 34.11 76.16 ;
    END
  END chany_top_out[7]
  PIN chany_top_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.71 74.8 42.85 76.16 ;
    END
  END chany_top_out[8]
  PIN chany_top_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.01 74.8 22.15 76.16 ;
    END
  END chany_top_out[9]
  PIN chany_top_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.65 74.8 37.79 76.16 ;
    END
  END chany_top_out[10]
  PIN chany_top_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.21 74.8 31.35 76.16 ;
    END
  END chany_top_out[11]
  PIN chany_top_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.37 74.8 29.51 76.16 ;
    END
  END chany_top_out[12]
  PIN chany_top_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.83 74.8 52.97 76.16 ;
    END
  END chany_top_out[13]
  PIN chany_top_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.97 74.8 57.11 76.16 ;
    END
  END chany_top_out[14]
  PIN chany_top_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.19 74.8 14.33 76.16 ;
    END
  END chany_top_out[15]
  PIN chany_top_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.05 74.8 33.19 76.16 ;
    END
  END chany_top_out[16]
  PIN chany_top_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.05 74.8 56.19 76.16 ;
    END
  END chany_top_out[17]
  PIN chany_top_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.89 74.8 58.03 76.16 ;
    END
  END chany_top_out[18]
  PIN chany_top_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.81 74.8 35.95 76.16 ;
    END
  END chany_top_out[19]
  PIN left_grid_pin_16_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 13.45 1.38 13.75 ;
    END
  END left_grid_pin_16_[0]
  PIN left_grid_pin_17_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 22.97 1.38 23.27 ;
    END
  END left_grid_pin_17_[0]
  PIN left_grid_pin_18_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 24.33 1.38 24.63 ;
    END
  END left_grid_pin_18_[0]
  PIN left_grid_pin_19_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 6.65 1.38 6.95 ;
    END
  END left_grid_pin_19_[0]
  PIN left_grid_pin_20_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 20.25 1.38 20.55 ;
    END
  END left_grid_pin_20_[0]
  PIN left_grid_pin_21_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 16.17 1.38 16.47 ;
    END
  END left_grid_pin_21_[0]
  PIN left_grid_pin_22_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 14.81 1.38 15.11 ;
    END
  END left_grid_pin_22_[0]
  PIN left_grid_pin_23_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 5.29 1.38 5.59 ;
    END
  END left_grid_pin_23_[0]
  PIN left_grid_pin_24_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 37.93 1.38 38.23 ;
    END
  END left_grid_pin_24_[0]
  PIN left_grid_pin_25_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 17.53 1.38 17.83 ;
    END
  END left_grid_pin_25_[0]
  PIN left_grid_pin_26_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 18.89 1.38 19.19 ;
    END
  END left_grid_pin_26_[0]
  PIN left_grid_pin_27_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 21.61 1.38 21.91 ;
    END
  END left_grid_pin_27_[0]
  PIN left_grid_pin_28_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 40.65 1.38 40.95 ;
    END
  END left_grid_pin_28_[0]
  PIN left_grid_pin_29_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 39.29 1.38 39.59 ;
    END
  END left_grid_pin_29_[0]
  PIN left_grid_pin_30_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 42.01 1.38 42.31 ;
    END
  END left_grid_pin_30_[0]
  PIN left_grid_pin_31_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 59.69 1.38 59.99 ;
    END
  END left_grid_pin_31_[0]
  PIN ccff_tail[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 64.86 40.65 66.24 40.95 ;
    END
  END ccff_tail[0]
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 0.48 2.96 ;
        RECT 65.76 2.48 66.24 2.96 ;
        RECT 0 7.92 0.48 8.4 ;
        RECT 65.76 7.92 66.24 8.4 ;
        RECT 0 13.36 0.48 13.84 ;
        RECT 65.76 13.36 66.24 13.84 ;
        RECT 0 18.8 0.48 19.28 ;
        RECT 65.76 18.8 66.24 19.28 ;
        RECT 0 24.24 0.48 24.72 ;
        RECT 65.76 24.24 66.24 24.72 ;
        RECT 0 29.68 0.48 30.16 ;
        RECT 65.76 29.68 66.24 30.16 ;
        RECT 0 35.12 0.48 35.6 ;
        RECT 65.76 35.12 66.24 35.6 ;
        RECT 0 40.56 0.48 41.04 ;
        RECT 65.76 40.56 66.24 41.04 ;
        RECT 0 46 0.48 46.48 ;
        RECT 65.76 46 66.24 46.48 ;
        RECT 0 51.44 0.48 51.92 ;
        RECT 65.76 51.44 66.24 51.92 ;
        RECT 0 56.88 0.48 57.36 ;
        RECT 65.76 56.88 66.24 57.36 ;
        RECT 0 62.32 0.48 62.8 ;
        RECT 65.76 62.32 66.24 62.8 ;
        RECT 0 67.76 0.48 68.24 ;
        RECT 65.76 67.76 66.24 68.24 ;
        RECT 0 73.2 0.48 73.68 ;
        RECT 65.76 73.2 66.24 73.68 ;
      LAYER met5 ;
        RECT 0 36.48 3.2 39.68 ;
        RECT 63.04 36.48 66.24 39.68 ;
      LAYER met4 ;
        RECT 10.74 0 11.34 0.6 ;
        RECT 40.18 0 40.78 0.6 ;
        RECT 10.74 75.56 11.34 76.16 ;
        RECT 40.18 75.56 40.78 76.16 ;
    END
  END VDD
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 0 66.24 0.24 ;
        RECT 0 5.2 0.48 5.68 ;
        RECT 65.76 5.2 66.24 5.68 ;
        RECT 0 10.64 0.48 11.12 ;
        RECT 65.76 10.64 66.24 11.12 ;
        RECT 0 16.08 0.48 16.56 ;
        RECT 65.76 16.08 66.24 16.56 ;
        RECT 0 21.52 0.48 22 ;
        RECT 65.76 21.52 66.24 22 ;
        RECT 0 26.96 0.48 27.44 ;
        RECT 65.76 26.96 66.24 27.44 ;
        RECT 0 32.4 0.48 32.88 ;
        RECT 65.76 32.4 66.24 32.88 ;
        RECT 0 37.84 0.48 38.32 ;
        RECT 65.76 37.84 66.24 38.32 ;
        RECT 0 43.28 0.48 43.76 ;
        RECT 65.76 43.28 66.24 43.76 ;
        RECT 0 48.72 0.48 49.2 ;
        RECT 65.76 48.72 66.24 49.2 ;
        RECT 0 54.16 0.48 54.64 ;
        RECT 65.76 54.16 66.24 54.64 ;
        RECT 0 59.6 0.48 60.08 ;
        RECT 65.76 59.6 66.24 60.08 ;
        RECT 0 65.04 0.48 65.52 ;
        RECT 65.76 65.04 66.24 65.52 ;
        RECT 0 70.48 0.48 70.96 ;
        RECT 65.76 70.48 66.24 70.96 ;
        RECT 0 75.92 66.24 76.16 ;
      LAYER met5 ;
        RECT 0 16.08 3.2 19.28 ;
        RECT 63.04 16.08 66.24 19.28 ;
        RECT 0 56.88 3.2 60.08 ;
        RECT 63.04 56.88 66.24 60.08 ;
      LAYER met4 ;
        RECT 25.46 0 26.06 0.6 ;
        RECT 54.9 0 55.5 0.6 ;
        RECT 25.46 75.56 26.06 76.16 ;
        RECT 54.9 75.56 55.5 76.16 ;
    END
  END VSS
  OBS
    LAYER li1 ;
      RECT 0 76.075 66.24 76.245 ;
      RECT 65.32 73.355 66.24 73.525 ;
      RECT 0 73.355 3.68 73.525 ;
      RECT 65.32 70.635 66.24 70.805 ;
      RECT 0 70.635 1.84 70.805 ;
      RECT 65.32 67.915 66.24 68.085 ;
      RECT 0 67.915 1.84 68.085 ;
      RECT 65.32 65.195 66.24 65.365 ;
      RECT 0 65.195 1.84 65.365 ;
      RECT 65.32 62.475 66.24 62.645 ;
      RECT 0 62.475 1.84 62.645 ;
      RECT 65.32 59.755 66.24 59.925 ;
      RECT 0 59.755 1.84 59.925 ;
      RECT 65.32 57.035 66.24 57.205 ;
      RECT 0 57.035 1.84 57.205 ;
      RECT 65.32 54.315 66.24 54.485 ;
      RECT 0 54.315 1.84 54.485 ;
      RECT 65.32 51.595 66.24 51.765 ;
      RECT 0 51.595 1.84 51.765 ;
      RECT 65.32 48.875 66.24 49.045 ;
      RECT 0 48.875 1.84 49.045 ;
      RECT 65.32 46.155 66.24 46.325 ;
      RECT 0 46.155 3.68 46.325 ;
      RECT 65.32 43.435 66.24 43.605 ;
      RECT 0 43.435 3.68 43.605 ;
      RECT 65.32 40.715 66.24 40.885 ;
      RECT 0 40.715 1.84 40.885 ;
      RECT 65.32 37.995 66.24 38.165 ;
      RECT 0 37.995 1.84 38.165 ;
      RECT 65.32 35.275 66.24 35.445 ;
      RECT 0 35.275 3.68 35.445 ;
      RECT 65.32 32.555 66.24 32.725 ;
      RECT 0 32.555 3.68 32.725 ;
      RECT 65.32 29.835 66.24 30.005 ;
      RECT 0 29.835 1.84 30.005 ;
      RECT 65.32 27.115 66.24 27.285 ;
      RECT 0 27.115 1.84 27.285 ;
      RECT 65.32 24.395 66.24 24.565 ;
      RECT 0 24.395 1.84 24.565 ;
      RECT 65.32 21.675 66.24 21.845 ;
      RECT 0 21.675 1.84 21.845 ;
      RECT 65.32 18.955 66.24 19.125 ;
      RECT 0 18.955 1.84 19.125 ;
      RECT 65.32 16.235 66.24 16.405 ;
      RECT 0 16.235 1.84 16.405 ;
      RECT 65.32 13.515 66.24 13.685 ;
      RECT 0 13.515 1.84 13.685 ;
      RECT 65.32 10.795 66.24 10.965 ;
      RECT 0 10.795 3.68 10.965 ;
      RECT 65.32 8.075 66.24 8.245 ;
      RECT 0 8.075 3.68 8.245 ;
      RECT 65.32 5.355 66.24 5.525 ;
      RECT 0 5.355 1.84 5.525 ;
      RECT 65.32 2.635 66.24 2.805 ;
      RECT 0 2.635 3.68 2.805 ;
      RECT 0 -0.085 66.24 0.085 ;
    LAYER met3 ;
      POLYGON 55.365 76.325 55.365 76.32 55.58 76.32 55.58 76 55.365 76 55.365 75.995 55.035 75.995 55.035 76 54.82 76 54.82 76.32 55.035 76.32 55.035 76.325 ;
      POLYGON 25.925 76.325 25.925 76.32 26.14 76.32 26.14 76 25.925 76 25.925 75.995 25.595 75.995 25.595 76 25.38 76 25.38 76.32 25.595 76.32 25.595 76.325 ;
      POLYGON 55.365 0.165 55.365 0.16 55.58 0.16 55.58 -0.16 55.365 -0.16 55.365 -0.165 55.035 -0.165 55.035 -0.16 54.82 -0.16 54.82 0.16 55.035 0.16 55.035 0.165 ;
      POLYGON 25.925 0.165 25.925 0.16 26.14 0.16 26.14 -0.16 25.925 -0.16 25.925 -0.165 25.595 -0.165 25.595 -0.16 25.38 -0.16 25.38 0.16 25.595 0.16 25.595 0.165 ;
      POLYGON 65.84 75.76 65.84 41.35 64.46 41.35 64.46 40.25 65.84 40.25 65.84 0.4 0.4 0.4 0.4 2.85 1.78 2.85 1.78 3.95 0.4 3.95 0.4 4.89 1.78 4.89 1.78 5.99 0.4 5.99 0.4 6.25 1.78 6.25 1.78 7.35 0.4 7.35 0.4 13.05 1.78 13.05 1.78 14.15 0.4 14.15 0.4 14.41 1.78 14.41 1.78 15.51 0.4 15.51 0.4 15.77 1.78 15.77 1.78 16.87 0.4 16.87 0.4 17.13 1.78 17.13 1.78 18.23 0.4 18.23 0.4 18.49 1.78 18.49 1.78 19.59 0.4 19.59 0.4 19.85 1.78 19.85 1.78 20.95 0.4 20.95 0.4 21.21 1.78 21.21 1.78 22.31 0.4 22.31 0.4 22.57 1.78 22.57 1.78 23.67 0.4 23.67 0.4 23.93 1.78 23.93 1.78 25.03 0.4 25.03 0.4 37.53 1.78 37.53 1.78 38.63 0.4 38.63 0.4 38.89 1.78 38.89 1.78 39.99 0.4 39.99 0.4 40.25 1.78 40.25 1.78 41.35 0.4 41.35 0.4 41.61 1.78 41.61 1.78 42.71 0.4 42.71 0.4 57.93 1.78 57.93 1.78 59.03 0.4 59.03 0.4 59.29 1.78 59.29 1.78 60.39 0.4 60.39 0.4 75.76 ;
    LAYER met2 ;
      RECT 55.06 75.975 55.34 76.345 ;
      RECT 25.62 75.975 25.9 76.345 ;
      RECT 56.45 74.3 56.71 74.62 ;
      RECT 45.41 74.3 45.67 74.62 ;
      RECT 23.33 74.3 23.59 74.62 ;
      RECT 34.37 1.54 34.63 1.86 ;
      RECT 55.06 -0.185 55.34 0.185 ;
      RECT 25.62 -0.185 25.9 0.185 ;
      POLYGON 65.96 75.88 65.96 0.28 59.69 0.28 59.69 1.64 58.99 1.64 58.99 0.28 58.31 0.28 58.31 1.64 57.61 1.64 57.61 0.28 57.39 0.28 57.39 1.64 56.69 1.64 56.69 0.28 56.47 0.28 56.47 1.64 55.77 1.64 55.77 0.28 54.63 0.28 54.63 1.64 53.93 1.64 53.93 0.28 53.71 0.28 53.71 1.64 53.01 1.64 53.01 0.28 52.79 0.28 52.79 1.64 52.09 1.64 52.09 0.28 51.87 0.28 51.87 1.64 51.17 1.64 51.17 0.28 50.95 0.28 50.95 1.64 50.25 1.64 50.25 0.28 50.03 0.28 50.03 1.64 49.33 1.64 49.33 0.28 48.65 0.28 48.65 1.64 47.95 1.64 47.95 0.28 47.73 0.28 47.73 1.64 47.03 1.64 47.03 0.28 46.81 0.28 46.81 1.64 46.11 1.64 46.11 0.28 45.89 0.28 45.89 1.64 45.19 1.64 45.19 0.28 44.51 0.28 44.51 1.64 43.81 1.64 43.81 0.28 43.13 0.28 43.13 1.64 42.43 1.64 42.43 0.28 42.21 0.28 42.21 1.64 41.51 1.64 41.51 0.28 41.29 0.28 41.29 1.64 40.59 1.64 40.59 0.28 40.37 0.28 40.37 1.64 39.67 1.64 39.67 0.28 38.99 0.28 38.99 1.64 38.29 1.64 38.29 0.28 38.07 0.28 38.07 1.64 37.37 1.64 37.37 0.28 37.15 0.28 37.15 1.64 36.45 1.64 36.45 0.28 36.23 0.28 36.23 1.64 35.53 1.64 35.53 0.28 35.31 0.28 35.31 1.64 34.61 1.64 34.61 0.28 34.39 0.28 34.39 1.64 33.69 1.64 33.69 0.28 33.47 0.28 33.47 1.64 32.77 1.64 32.77 0.28 32.55 0.28 32.55 1.64 31.85 1.64 31.85 0.28 31.63 0.28 31.63 1.64 30.93 1.64 30.93 0.28 30.25 0.28 30.25 1.64 29.55 1.64 29.55 0.28 29.33 0.28 29.33 1.64 28.63 1.64 28.63 0.28 28.41 0.28 28.41 1.64 27.71 1.64 27.71 0.28 27.49 0.28 27.49 1.64 26.79 1.64 26.79 0.28 25.19 0.28 25.19 1.64 24.49 1.64 24.49 0.28 24.27 0.28 24.27 1.64 23.57 1.64 23.57 0.28 22.89 0.28 22.89 1.64 22.19 1.64 22.19 0.28 21.97 0.28 21.97 1.64 21.27 1.64 21.27 0.28 21.05 0.28 21.05 1.64 20.35 1.64 20.35 0.28 0.28 0.28 0.28 75.88 13.91 75.88 13.91 74.52 14.61 74.52 14.61 75.88 14.83 75.88 14.83 74.52 15.53 74.52 15.53 75.88 20.81 75.88 20.81 74.52 21.51 74.52 21.51 75.88 21.73 75.88 21.73 74.52 22.43 74.52 22.43 75.88 22.65 75.88 22.65 74.52 23.35 74.52 23.35 75.88 23.57 75.88 23.57 74.52 24.27 74.52 24.27 75.88 24.49 75.88 24.49 74.52 25.19 74.52 25.19 75.88 26.33 75.88 26.33 74.52 27.03 74.52 27.03 75.88 27.25 75.88 27.25 74.52 27.95 74.52 27.95 75.88 28.17 75.88 28.17 74.52 28.87 74.52 28.87 75.88 29.09 75.88 29.09 74.52 29.79 74.52 29.79 75.88 30.01 75.88 30.01 74.52 30.71 74.52 30.71 75.88 30.93 75.88 30.93 74.52 31.63 74.52 31.63 75.88 31.85 75.88 31.85 74.52 32.55 74.52 32.55 75.88 32.77 75.88 32.77 74.52 33.47 74.52 33.47 75.88 33.69 75.88 33.69 74.52 34.39 74.52 34.39 75.88 35.53 75.88 35.53 74.52 36.23 74.52 36.23 75.88 36.45 75.88 36.45 74.52 37.15 74.52 37.15 75.88 37.37 75.88 37.37 74.52 38.07 74.52 38.07 75.88 38.29 75.88 38.29 74.52 38.99 74.52 38.99 75.88 39.21 75.88 39.21 74.52 39.91 74.52 39.91 75.88 40.59 75.88 40.59 74.52 41.29 74.52 41.29 75.88 41.51 75.88 41.51 74.52 42.21 74.52 42.21 75.88 42.43 75.88 42.43 74.52 43.13 74.52 43.13 75.88 43.81 75.88 43.81 74.52 44.51 74.52 44.51 75.88 44.73 75.88 44.73 74.52 45.43 74.52 45.43 75.88 46.11 75.88 46.11 74.52 46.81 74.52 46.81 75.88 47.03 75.88 47.03 74.52 47.73 74.52 47.73 75.88 47.95 75.88 47.95 74.52 48.65 74.52 48.65 75.88 48.87 75.88 48.87 74.52 49.57 74.52 49.57 75.88 49.79 75.88 49.79 74.52 50.49 74.52 50.49 75.88 50.71 75.88 50.71 74.52 51.41 74.52 51.41 75.88 51.63 75.88 51.63 74.52 52.33 74.52 52.33 75.88 52.55 75.88 52.55 74.52 53.25 74.52 53.25 75.88 53.47 75.88 53.47 74.52 54.17 74.52 54.17 75.88 55.77 75.88 55.77 74.52 56.47 74.52 56.47 75.88 56.69 75.88 56.69 74.52 57.39 74.52 57.39 75.88 57.61 75.88 57.61 74.52 58.31 74.52 58.31 75.88 58.53 75.88 58.53 74.52 59.23 74.52 59.23 75.88 62.21 75.88 62.21 74.52 62.91 74.52 62.91 75.88 ;
    LAYER met4 ;
      POLYGON 65.84 75.76 65.84 0.4 55.9 0.4 55.9 1 54.5 1 54.5 0.4 44.71 0.4 44.71 1.76 43.61 1.76 43.61 0.4 42.87 0.4 42.87 1.76 41.77 1.76 41.77 0.4 41.18 0.4 41.18 1 39.78 1 39.78 0.4 38.27 0.4 38.27 1.76 37.17 1.76 37.17 0.4 26.46 0.4 26.46 1 25.06 1 25.06 0.4 11.74 0.4 11.74 1 10.34 1 10.34 0.4 0.4 0.4 0.4 75.76 10.34 75.76 10.34 75.16 11.74 75.16 11.74 75.76 25.06 75.76 25.06 75.16 26.46 75.16 26.46 75.76 39.78 75.76 39.78 75.16 41.18 75.16 41.18 75.76 54.5 75.76 54.5 75.16 55.9 75.16 55.9 75.76 ;
    LAYER met5 ;
      POLYGON 64.64 74.56 64.64 61.68 61.44 61.68 61.44 55.28 64.64 55.28 64.64 41.28 61.44 41.28 61.44 34.88 64.64 34.88 64.64 20.88 61.44 20.88 61.44 14.48 64.64 14.48 64.64 1.6 1.6 1.6 1.6 14.48 4.8 14.48 4.8 20.88 1.6 20.88 1.6 34.88 4.8 34.88 4.8 41.28 1.6 41.28 1.6 55.28 4.8 55.28 4.8 61.68 1.6 61.68 1.6 74.56 ;
    LAYER met1 ;
      POLYGON 65.96 75.64 65.96 73.96 65.48 73.96 65.48 72.92 65.96 72.92 65.96 71.24 65.48 71.24 65.48 70.2 65.96 70.2 65.96 68.52 65.48 68.52 65.48 67.48 65.96 67.48 65.96 65.8 65.48 65.8 65.48 64.76 65.96 64.76 65.96 63.08 65.48 63.08 65.48 62.04 65.96 62.04 65.96 60.36 65.48 60.36 65.48 59.32 65.96 59.32 65.96 57.64 65.48 57.64 65.48 56.6 65.96 56.6 65.96 54.92 65.48 54.92 65.48 53.88 65.96 53.88 65.96 52.2 65.48 52.2 65.48 51.16 65.96 51.16 65.96 49.48 65.48 49.48 65.48 48.44 65.96 48.44 65.96 46.76 65.48 46.76 65.48 45.72 65.96 45.72 65.96 44.04 65.48 44.04 65.48 43 65.96 43 65.96 41.32 65.48 41.32 65.48 40.28 65.96 40.28 65.96 38.6 65.48 38.6 65.48 37.56 65.96 37.56 65.96 35.88 65.48 35.88 65.48 34.84 65.96 34.84 65.96 33.16 65.48 33.16 65.48 32.12 65.96 32.12 65.96 30.44 65.48 30.44 65.48 29.4 65.96 29.4 65.96 27.72 65.48 27.72 65.48 26.68 65.96 26.68 65.96 25 65.48 25 65.48 23.96 65.96 23.96 65.96 22.28 65.48 22.28 65.48 21.24 65.96 21.24 65.96 19.56 65.48 19.56 65.48 18.52 65.96 18.52 65.96 16.84 65.48 16.84 65.48 15.8 65.96 15.8 65.96 14.12 65.48 14.12 65.48 13.08 65.96 13.08 65.96 11.4 65.48 11.4 65.48 10.36 65.96 10.36 65.96 8.68 65.48 8.68 65.48 7.64 65.96 7.64 65.96 5.96 65.48 5.96 65.48 4.92 65.96 4.92 65.96 3.24 65.48 3.24 65.48 2.2 65.96 2.2 65.96 0.52 0.28 0.52 0.28 2.2 0.76 2.2 0.76 3.24 0.28 3.24 0.28 4.92 0.76 4.92 0.76 5.96 0.28 5.96 0.28 7.64 0.76 7.64 0.76 8.68 0.28 8.68 0.28 10.36 0.76 10.36 0.76 11.4 0.28 11.4 0.28 13.08 0.76 13.08 0.76 14.12 0.28 14.12 0.28 15.8 0.76 15.8 0.76 16.84 0.28 16.84 0.28 18.52 0.76 18.52 0.76 19.56 0.28 19.56 0.28 21.24 0.76 21.24 0.76 22.28 0.28 22.28 0.28 23.96 0.76 23.96 0.76 25 0.28 25 0.28 26.68 0.76 26.68 0.76 27.72 0.28 27.72 0.28 29.4 0.76 29.4 0.76 30.44 0.28 30.44 0.28 32.12 0.76 32.12 0.76 33.16 0.28 33.16 0.28 34.84 0.76 34.84 0.76 35.88 0.28 35.88 0.28 37.56 0.76 37.56 0.76 38.6 0.28 38.6 0.28 40.28 0.76 40.28 0.76 41.32 0.28 41.32 0.28 43 0.76 43 0.76 44.04 0.28 44.04 0.28 45.72 0.76 45.72 0.76 46.76 0.28 46.76 0.28 48.44 0.76 48.44 0.76 49.48 0.28 49.48 0.28 51.16 0.76 51.16 0.76 52.2 0.28 52.2 0.28 53.88 0.76 53.88 0.76 54.92 0.28 54.92 0.28 56.6 0.76 56.6 0.76 57.64 0.28 57.64 0.28 59.32 0.76 59.32 0.76 60.36 0.28 60.36 0.28 62.04 0.76 62.04 0.76 63.08 0.28 63.08 0.28 64.76 0.76 64.76 0.76 65.8 0.28 65.8 0.28 67.48 0.76 67.48 0.76 68.52 0.28 68.52 0.28 70.2 0.76 70.2 0.76 71.24 0.28 71.24 0.28 72.92 0.76 72.92 0.76 73.96 0.28 73.96 0.28 75.64 ;
    LAYER li1 ;
      RECT 0.17 0.17 66.07 75.99 ;
    LAYER mcon ;
      RECT 65.925 76.075 66.095 76.245 ;
      RECT 65.465 76.075 65.635 76.245 ;
      RECT 65.005 76.075 65.175 76.245 ;
      RECT 64.545 76.075 64.715 76.245 ;
      RECT 64.085 76.075 64.255 76.245 ;
      RECT 63.625 76.075 63.795 76.245 ;
      RECT 63.165 76.075 63.335 76.245 ;
      RECT 62.705 76.075 62.875 76.245 ;
      RECT 62.245 76.075 62.415 76.245 ;
      RECT 61.785 76.075 61.955 76.245 ;
      RECT 61.325 76.075 61.495 76.245 ;
      RECT 60.865 76.075 61.035 76.245 ;
      RECT 60.405 76.075 60.575 76.245 ;
      RECT 59.945 76.075 60.115 76.245 ;
      RECT 59.485 76.075 59.655 76.245 ;
      RECT 59.025 76.075 59.195 76.245 ;
      RECT 58.565 76.075 58.735 76.245 ;
      RECT 58.105 76.075 58.275 76.245 ;
      RECT 57.645 76.075 57.815 76.245 ;
      RECT 57.185 76.075 57.355 76.245 ;
      RECT 56.725 76.075 56.895 76.245 ;
      RECT 56.265 76.075 56.435 76.245 ;
      RECT 55.805 76.075 55.975 76.245 ;
      RECT 55.345 76.075 55.515 76.245 ;
      RECT 54.885 76.075 55.055 76.245 ;
      RECT 54.425 76.075 54.595 76.245 ;
      RECT 53.965 76.075 54.135 76.245 ;
      RECT 53.505 76.075 53.675 76.245 ;
      RECT 53.045 76.075 53.215 76.245 ;
      RECT 52.585 76.075 52.755 76.245 ;
      RECT 52.125 76.075 52.295 76.245 ;
      RECT 51.665 76.075 51.835 76.245 ;
      RECT 51.205 76.075 51.375 76.245 ;
      RECT 50.745 76.075 50.915 76.245 ;
      RECT 50.285 76.075 50.455 76.245 ;
      RECT 49.825 76.075 49.995 76.245 ;
      RECT 49.365 76.075 49.535 76.245 ;
      RECT 48.905 76.075 49.075 76.245 ;
      RECT 48.445 76.075 48.615 76.245 ;
      RECT 47.985 76.075 48.155 76.245 ;
      RECT 47.525 76.075 47.695 76.245 ;
      RECT 47.065 76.075 47.235 76.245 ;
      RECT 46.605 76.075 46.775 76.245 ;
      RECT 46.145 76.075 46.315 76.245 ;
      RECT 45.685 76.075 45.855 76.245 ;
      RECT 45.225 76.075 45.395 76.245 ;
      RECT 44.765 76.075 44.935 76.245 ;
      RECT 44.305 76.075 44.475 76.245 ;
      RECT 43.845 76.075 44.015 76.245 ;
      RECT 43.385 76.075 43.555 76.245 ;
      RECT 42.925 76.075 43.095 76.245 ;
      RECT 42.465 76.075 42.635 76.245 ;
      RECT 42.005 76.075 42.175 76.245 ;
      RECT 41.545 76.075 41.715 76.245 ;
      RECT 41.085 76.075 41.255 76.245 ;
      RECT 40.625 76.075 40.795 76.245 ;
      RECT 40.165 76.075 40.335 76.245 ;
      RECT 39.705 76.075 39.875 76.245 ;
      RECT 39.245 76.075 39.415 76.245 ;
      RECT 38.785 76.075 38.955 76.245 ;
      RECT 38.325 76.075 38.495 76.245 ;
      RECT 37.865 76.075 38.035 76.245 ;
      RECT 37.405 76.075 37.575 76.245 ;
      RECT 36.945 76.075 37.115 76.245 ;
      RECT 36.485 76.075 36.655 76.245 ;
      RECT 36.025 76.075 36.195 76.245 ;
      RECT 35.565 76.075 35.735 76.245 ;
      RECT 35.105 76.075 35.275 76.245 ;
      RECT 34.645 76.075 34.815 76.245 ;
      RECT 34.185 76.075 34.355 76.245 ;
      RECT 33.725 76.075 33.895 76.245 ;
      RECT 33.265 76.075 33.435 76.245 ;
      RECT 32.805 76.075 32.975 76.245 ;
      RECT 32.345 76.075 32.515 76.245 ;
      RECT 31.885 76.075 32.055 76.245 ;
      RECT 31.425 76.075 31.595 76.245 ;
      RECT 30.965 76.075 31.135 76.245 ;
      RECT 30.505 76.075 30.675 76.245 ;
      RECT 30.045 76.075 30.215 76.245 ;
      RECT 29.585 76.075 29.755 76.245 ;
      RECT 29.125 76.075 29.295 76.245 ;
      RECT 28.665 76.075 28.835 76.245 ;
      RECT 28.205 76.075 28.375 76.245 ;
      RECT 27.745 76.075 27.915 76.245 ;
      RECT 27.285 76.075 27.455 76.245 ;
      RECT 26.825 76.075 26.995 76.245 ;
      RECT 26.365 76.075 26.535 76.245 ;
      RECT 25.905 76.075 26.075 76.245 ;
      RECT 25.445 76.075 25.615 76.245 ;
      RECT 24.985 76.075 25.155 76.245 ;
      RECT 24.525 76.075 24.695 76.245 ;
      RECT 24.065 76.075 24.235 76.245 ;
      RECT 23.605 76.075 23.775 76.245 ;
      RECT 23.145 76.075 23.315 76.245 ;
      RECT 22.685 76.075 22.855 76.245 ;
      RECT 22.225 76.075 22.395 76.245 ;
      RECT 21.765 76.075 21.935 76.245 ;
      RECT 21.305 76.075 21.475 76.245 ;
      RECT 20.845 76.075 21.015 76.245 ;
      RECT 20.385 76.075 20.555 76.245 ;
      RECT 19.925 76.075 20.095 76.245 ;
      RECT 19.465 76.075 19.635 76.245 ;
      RECT 19.005 76.075 19.175 76.245 ;
      RECT 18.545 76.075 18.715 76.245 ;
      RECT 18.085 76.075 18.255 76.245 ;
      RECT 17.625 76.075 17.795 76.245 ;
      RECT 17.165 76.075 17.335 76.245 ;
      RECT 16.705 76.075 16.875 76.245 ;
      RECT 16.245 76.075 16.415 76.245 ;
      RECT 15.785 76.075 15.955 76.245 ;
      RECT 15.325 76.075 15.495 76.245 ;
      RECT 14.865 76.075 15.035 76.245 ;
      RECT 14.405 76.075 14.575 76.245 ;
      RECT 13.945 76.075 14.115 76.245 ;
      RECT 13.485 76.075 13.655 76.245 ;
      RECT 13.025 76.075 13.195 76.245 ;
      RECT 12.565 76.075 12.735 76.245 ;
      RECT 12.105 76.075 12.275 76.245 ;
      RECT 11.645 76.075 11.815 76.245 ;
      RECT 11.185 76.075 11.355 76.245 ;
      RECT 10.725 76.075 10.895 76.245 ;
      RECT 10.265 76.075 10.435 76.245 ;
      RECT 9.805 76.075 9.975 76.245 ;
      RECT 9.345 76.075 9.515 76.245 ;
      RECT 8.885 76.075 9.055 76.245 ;
      RECT 8.425 76.075 8.595 76.245 ;
      RECT 7.965 76.075 8.135 76.245 ;
      RECT 7.505 76.075 7.675 76.245 ;
      RECT 7.045 76.075 7.215 76.245 ;
      RECT 6.585 76.075 6.755 76.245 ;
      RECT 6.125 76.075 6.295 76.245 ;
      RECT 5.665 76.075 5.835 76.245 ;
      RECT 5.205 76.075 5.375 76.245 ;
      RECT 4.745 76.075 4.915 76.245 ;
      RECT 4.285 76.075 4.455 76.245 ;
      RECT 3.825 76.075 3.995 76.245 ;
      RECT 3.365 76.075 3.535 76.245 ;
      RECT 2.905 76.075 3.075 76.245 ;
      RECT 2.445 76.075 2.615 76.245 ;
      RECT 1.985 76.075 2.155 76.245 ;
      RECT 1.525 76.075 1.695 76.245 ;
      RECT 1.065 76.075 1.235 76.245 ;
      RECT 0.605 76.075 0.775 76.245 ;
      RECT 0.145 76.075 0.315 76.245 ;
      RECT 65.925 73.355 66.095 73.525 ;
      RECT 65.465 73.355 65.635 73.525 ;
      RECT 0.605 73.355 0.775 73.525 ;
      RECT 0.145 73.355 0.315 73.525 ;
      RECT 65.925 70.635 66.095 70.805 ;
      RECT 65.465 70.635 65.635 70.805 ;
      RECT 0.605 70.635 0.775 70.805 ;
      RECT 0.145 70.635 0.315 70.805 ;
      RECT 65.925 67.915 66.095 68.085 ;
      RECT 65.465 67.915 65.635 68.085 ;
      RECT 0.605 67.915 0.775 68.085 ;
      RECT 0.145 67.915 0.315 68.085 ;
      RECT 65.925 65.195 66.095 65.365 ;
      RECT 65.465 65.195 65.635 65.365 ;
      RECT 0.605 65.195 0.775 65.365 ;
      RECT 0.145 65.195 0.315 65.365 ;
      RECT 65.925 62.475 66.095 62.645 ;
      RECT 65.465 62.475 65.635 62.645 ;
      RECT 0.605 62.475 0.775 62.645 ;
      RECT 0.145 62.475 0.315 62.645 ;
      RECT 65.925 59.755 66.095 59.925 ;
      RECT 65.465 59.755 65.635 59.925 ;
      RECT 0.605 59.755 0.775 59.925 ;
      RECT 0.145 59.755 0.315 59.925 ;
      RECT 65.925 57.035 66.095 57.205 ;
      RECT 65.465 57.035 65.635 57.205 ;
      RECT 0.605 57.035 0.775 57.205 ;
      RECT 0.145 57.035 0.315 57.205 ;
      RECT 65.925 54.315 66.095 54.485 ;
      RECT 65.465 54.315 65.635 54.485 ;
      RECT 0.605 54.315 0.775 54.485 ;
      RECT 0.145 54.315 0.315 54.485 ;
      RECT 65.925 51.595 66.095 51.765 ;
      RECT 65.465 51.595 65.635 51.765 ;
      RECT 0.605 51.595 0.775 51.765 ;
      RECT 0.145 51.595 0.315 51.765 ;
      RECT 65.925 48.875 66.095 49.045 ;
      RECT 65.465 48.875 65.635 49.045 ;
      RECT 0.605 48.875 0.775 49.045 ;
      RECT 0.145 48.875 0.315 49.045 ;
      RECT 65.925 46.155 66.095 46.325 ;
      RECT 65.465 46.155 65.635 46.325 ;
      RECT 0.605 46.155 0.775 46.325 ;
      RECT 0.145 46.155 0.315 46.325 ;
      RECT 65.925 43.435 66.095 43.605 ;
      RECT 65.465 43.435 65.635 43.605 ;
      RECT 0.605 43.435 0.775 43.605 ;
      RECT 0.145 43.435 0.315 43.605 ;
      RECT 65.925 40.715 66.095 40.885 ;
      RECT 65.465 40.715 65.635 40.885 ;
      RECT 0.605 40.715 0.775 40.885 ;
      RECT 0.145 40.715 0.315 40.885 ;
      RECT 65.925 37.995 66.095 38.165 ;
      RECT 65.465 37.995 65.635 38.165 ;
      RECT 0.605 37.995 0.775 38.165 ;
      RECT 0.145 37.995 0.315 38.165 ;
      RECT 65.925 35.275 66.095 35.445 ;
      RECT 65.465 35.275 65.635 35.445 ;
      RECT 0.605 35.275 0.775 35.445 ;
      RECT 0.145 35.275 0.315 35.445 ;
      RECT 65.925 32.555 66.095 32.725 ;
      RECT 65.465 32.555 65.635 32.725 ;
      RECT 0.605 32.555 0.775 32.725 ;
      RECT 0.145 32.555 0.315 32.725 ;
      RECT 65.925 29.835 66.095 30.005 ;
      RECT 65.465 29.835 65.635 30.005 ;
      RECT 0.605 29.835 0.775 30.005 ;
      RECT 0.145 29.835 0.315 30.005 ;
      RECT 65.925 27.115 66.095 27.285 ;
      RECT 65.465 27.115 65.635 27.285 ;
      RECT 0.605 27.115 0.775 27.285 ;
      RECT 0.145 27.115 0.315 27.285 ;
      RECT 65.925 24.395 66.095 24.565 ;
      RECT 65.465 24.395 65.635 24.565 ;
      RECT 0.605 24.395 0.775 24.565 ;
      RECT 0.145 24.395 0.315 24.565 ;
      RECT 65.925 21.675 66.095 21.845 ;
      RECT 65.465 21.675 65.635 21.845 ;
      RECT 0.605 21.675 0.775 21.845 ;
      RECT 0.145 21.675 0.315 21.845 ;
      RECT 65.925 18.955 66.095 19.125 ;
      RECT 65.465 18.955 65.635 19.125 ;
      RECT 0.605 18.955 0.775 19.125 ;
      RECT 0.145 18.955 0.315 19.125 ;
      RECT 65.925 16.235 66.095 16.405 ;
      RECT 65.465 16.235 65.635 16.405 ;
      RECT 0.605 16.235 0.775 16.405 ;
      RECT 0.145 16.235 0.315 16.405 ;
      RECT 65.925 13.515 66.095 13.685 ;
      RECT 65.465 13.515 65.635 13.685 ;
      RECT 0.605 13.515 0.775 13.685 ;
      RECT 0.145 13.515 0.315 13.685 ;
      RECT 65.925 10.795 66.095 10.965 ;
      RECT 65.465 10.795 65.635 10.965 ;
      RECT 0.605 10.795 0.775 10.965 ;
      RECT 0.145 10.795 0.315 10.965 ;
      RECT 65.925 8.075 66.095 8.245 ;
      RECT 65.465 8.075 65.635 8.245 ;
      RECT 0.605 8.075 0.775 8.245 ;
      RECT 0.145 8.075 0.315 8.245 ;
      RECT 65.925 5.355 66.095 5.525 ;
      RECT 65.465 5.355 65.635 5.525 ;
      RECT 0.605 5.355 0.775 5.525 ;
      RECT 0.145 5.355 0.315 5.525 ;
      RECT 65.925 2.635 66.095 2.805 ;
      RECT 65.465 2.635 65.635 2.805 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 65.925 -0.085 66.095 0.085 ;
      RECT 65.465 -0.085 65.635 0.085 ;
      RECT 65.005 -0.085 65.175 0.085 ;
      RECT 64.545 -0.085 64.715 0.085 ;
      RECT 64.085 -0.085 64.255 0.085 ;
      RECT 63.625 -0.085 63.795 0.085 ;
      RECT 63.165 -0.085 63.335 0.085 ;
      RECT 62.705 -0.085 62.875 0.085 ;
      RECT 62.245 -0.085 62.415 0.085 ;
      RECT 61.785 -0.085 61.955 0.085 ;
      RECT 61.325 -0.085 61.495 0.085 ;
      RECT 60.865 -0.085 61.035 0.085 ;
      RECT 60.405 -0.085 60.575 0.085 ;
      RECT 59.945 -0.085 60.115 0.085 ;
      RECT 59.485 -0.085 59.655 0.085 ;
      RECT 59.025 -0.085 59.195 0.085 ;
      RECT 58.565 -0.085 58.735 0.085 ;
      RECT 58.105 -0.085 58.275 0.085 ;
      RECT 57.645 -0.085 57.815 0.085 ;
      RECT 57.185 -0.085 57.355 0.085 ;
      RECT 56.725 -0.085 56.895 0.085 ;
      RECT 56.265 -0.085 56.435 0.085 ;
      RECT 55.805 -0.085 55.975 0.085 ;
      RECT 55.345 -0.085 55.515 0.085 ;
      RECT 54.885 -0.085 55.055 0.085 ;
      RECT 54.425 -0.085 54.595 0.085 ;
      RECT 53.965 -0.085 54.135 0.085 ;
      RECT 53.505 -0.085 53.675 0.085 ;
      RECT 53.045 -0.085 53.215 0.085 ;
      RECT 52.585 -0.085 52.755 0.085 ;
      RECT 52.125 -0.085 52.295 0.085 ;
      RECT 51.665 -0.085 51.835 0.085 ;
      RECT 51.205 -0.085 51.375 0.085 ;
      RECT 50.745 -0.085 50.915 0.085 ;
      RECT 50.285 -0.085 50.455 0.085 ;
      RECT 49.825 -0.085 49.995 0.085 ;
      RECT 49.365 -0.085 49.535 0.085 ;
      RECT 48.905 -0.085 49.075 0.085 ;
      RECT 48.445 -0.085 48.615 0.085 ;
      RECT 47.985 -0.085 48.155 0.085 ;
      RECT 47.525 -0.085 47.695 0.085 ;
      RECT 47.065 -0.085 47.235 0.085 ;
      RECT 46.605 -0.085 46.775 0.085 ;
      RECT 46.145 -0.085 46.315 0.085 ;
      RECT 45.685 -0.085 45.855 0.085 ;
      RECT 45.225 -0.085 45.395 0.085 ;
      RECT 44.765 -0.085 44.935 0.085 ;
      RECT 44.305 -0.085 44.475 0.085 ;
      RECT 43.845 -0.085 44.015 0.085 ;
      RECT 43.385 -0.085 43.555 0.085 ;
      RECT 42.925 -0.085 43.095 0.085 ;
      RECT 42.465 -0.085 42.635 0.085 ;
      RECT 42.005 -0.085 42.175 0.085 ;
      RECT 41.545 -0.085 41.715 0.085 ;
      RECT 41.085 -0.085 41.255 0.085 ;
      RECT 40.625 -0.085 40.795 0.085 ;
      RECT 40.165 -0.085 40.335 0.085 ;
      RECT 39.705 -0.085 39.875 0.085 ;
      RECT 39.245 -0.085 39.415 0.085 ;
      RECT 38.785 -0.085 38.955 0.085 ;
      RECT 38.325 -0.085 38.495 0.085 ;
      RECT 37.865 -0.085 38.035 0.085 ;
      RECT 37.405 -0.085 37.575 0.085 ;
      RECT 36.945 -0.085 37.115 0.085 ;
      RECT 36.485 -0.085 36.655 0.085 ;
      RECT 36.025 -0.085 36.195 0.085 ;
      RECT 35.565 -0.085 35.735 0.085 ;
      RECT 35.105 -0.085 35.275 0.085 ;
      RECT 34.645 -0.085 34.815 0.085 ;
      RECT 34.185 -0.085 34.355 0.085 ;
      RECT 33.725 -0.085 33.895 0.085 ;
      RECT 33.265 -0.085 33.435 0.085 ;
      RECT 32.805 -0.085 32.975 0.085 ;
      RECT 32.345 -0.085 32.515 0.085 ;
      RECT 31.885 -0.085 32.055 0.085 ;
      RECT 31.425 -0.085 31.595 0.085 ;
      RECT 30.965 -0.085 31.135 0.085 ;
      RECT 30.505 -0.085 30.675 0.085 ;
      RECT 30.045 -0.085 30.215 0.085 ;
      RECT 29.585 -0.085 29.755 0.085 ;
      RECT 29.125 -0.085 29.295 0.085 ;
      RECT 28.665 -0.085 28.835 0.085 ;
      RECT 28.205 -0.085 28.375 0.085 ;
      RECT 27.745 -0.085 27.915 0.085 ;
      RECT 27.285 -0.085 27.455 0.085 ;
      RECT 26.825 -0.085 26.995 0.085 ;
      RECT 26.365 -0.085 26.535 0.085 ;
      RECT 25.905 -0.085 26.075 0.085 ;
      RECT 25.445 -0.085 25.615 0.085 ;
      RECT 24.985 -0.085 25.155 0.085 ;
      RECT 24.525 -0.085 24.695 0.085 ;
      RECT 24.065 -0.085 24.235 0.085 ;
      RECT 23.605 -0.085 23.775 0.085 ;
      RECT 23.145 -0.085 23.315 0.085 ;
      RECT 22.685 -0.085 22.855 0.085 ;
      RECT 22.225 -0.085 22.395 0.085 ;
      RECT 21.765 -0.085 21.935 0.085 ;
      RECT 21.305 -0.085 21.475 0.085 ;
      RECT 20.845 -0.085 21.015 0.085 ;
      RECT 20.385 -0.085 20.555 0.085 ;
      RECT 19.925 -0.085 20.095 0.085 ;
      RECT 19.465 -0.085 19.635 0.085 ;
      RECT 19.005 -0.085 19.175 0.085 ;
      RECT 18.545 -0.085 18.715 0.085 ;
      RECT 18.085 -0.085 18.255 0.085 ;
      RECT 17.625 -0.085 17.795 0.085 ;
      RECT 17.165 -0.085 17.335 0.085 ;
      RECT 16.705 -0.085 16.875 0.085 ;
      RECT 16.245 -0.085 16.415 0.085 ;
      RECT 15.785 -0.085 15.955 0.085 ;
      RECT 15.325 -0.085 15.495 0.085 ;
      RECT 14.865 -0.085 15.035 0.085 ;
      RECT 14.405 -0.085 14.575 0.085 ;
      RECT 13.945 -0.085 14.115 0.085 ;
      RECT 13.485 -0.085 13.655 0.085 ;
      RECT 13.025 -0.085 13.195 0.085 ;
      RECT 12.565 -0.085 12.735 0.085 ;
      RECT 12.105 -0.085 12.275 0.085 ;
      RECT 11.645 -0.085 11.815 0.085 ;
      RECT 11.185 -0.085 11.355 0.085 ;
      RECT 10.725 -0.085 10.895 0.085 ;
      RECT 10.265 -0.085 10.435 0.085 ;
      RECT 9.805 -0.085 9.975 0.085 ;
      RECT 9.345 -0.085 9.515 0.085 ;
      RECT 8.885 -0.085 9.055 0.085 ;
      RECT 8.425 -0.085 8.595 0.085 ;
      RECT 7.965 -0.085 8.135 0.085 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.145 -0.085 0.315 0.085 ;
    LAYER via ;
      RECT 55.125 76.085 55.275 76.235 ;
      RECT 25.685 76.085 25.835 76.235 ;
      RECT 50.985 74.385 51.135 74.535 ;
      RECT 48.225 74.385 48.375 74.535 ;
      RECT 33.045 74.385 33.195 74.535 ;
      RECT 40.865 1.625 41.015 1.775 ;
      RECT 55.125 -0.075 55.275 0.075 ;
      RECT 25.685 -0.075 25.835 0.075 ;
    LAYER via2 ;
      RECT 55.1 76.06 55.3 76.26 ;
      RECT 25.66 76.06 25.86 76.26 ;
      RECT 1.74 58.38 1.94 58.58 ;
      RECT 1.74 21.66 1.94 21.86 ;
      RECT 1.28 16.22 1.48 16.42 ;
      RECT 1.28 13.5 1.48 13.7 ;
      RECT 55.1 -0.1 55.3 0.1 ;
      RECT 25.66 -0.1 25.86 0.1 ;
    LAYER via3 ;
      RECT 55.1 76.06 55.3 76.26 ;
      RECT 25.66 76.06 25.86 76.26 ;
      RECT 55.1 -0.1 55.3 0.1 ;
      RECT 25.66 -0.1 25.86 0.1 ;
    LAYER OVERLAP ;
      POLYGON 0 0 0 76.16 66.24 76.16 66.24 0 ;
  END
END cby_1__1_

END LIBRARY
