VERSION 5.7 ;
BUSBITCHARS "[]" ;

UNITS
  DATABASE MICRONS 1000 ;
END UNITS

MANUFACTURINGGRID 0.005 ;

LAYER li1
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.46 ;
  WIDTH 0.17 ;
END li1

LAYER mcon
  TYPE CUT ;
END mcon

LAYER met1
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.34 ;
  WIDTH 0.14 ;
END met1

LAYER via
  TYPE CUT ;
END via

LAYER met2
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.46 ;
  WIDTH 0.14 ;
END met2

LAYER via2
  TYPE CUT ;
END via2

LAYER met3
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.68 ;
  WIDTH 0.3 ;
END met3

LAYER via3
  TYPE CUT ;
END via3

LAYER met4
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.92 ;
  WIDTH 0.3 ;
END met4

LAYER via4
  TYPE CUT ;
END via4

LAYER met5
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 3.4 ;
  WIDTH 1.6 ;
END met5

LAYER nwell
  TYPE MASTERSLICE ;
END nwell

LAYER pwell
  TYPE MASTERSLICE ;
END pwell

LAYER OVERLAP
  TYPE OVERLAP ;
END OVERLAP

VIA L1M1_PR
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.145 -0.115 0.145 0.115 ;
END L1M1_PR

VIA L1M1_PR_R
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.115 -0.145 0.115 0.145 ;
END L1M1_PR_R

VIA L1M1_PR_M
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.115 -0.145 0.115 0.145 ;
END L1M1_PR_M

VIA L1M1_PR_MR
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.145 -0.115 0.145 0.115 ;
END L1M1_PR_MR

VIA L1M1_PR_C
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.145 -0.145 0.145 0.145 ;
END L1M1_PR_C

VIA M1M2_PR
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR

VIA M1M2_PR_Enc
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_Enc

VIA M1M2_PR_R
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_R

VIA M1M2_PR_R_Enc
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR_R_Enc

VIA M1M2_PR_M
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_M

VIA M1M2_PR_M_Enc
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR_M_Enc

VIA M1M2_PR_MR
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR_MR

VIA M1M2_PR_MR_Enc
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_MR_Enc

VIA M1M2_PR_C
  LAYER met1 ;
    RECT -0.16 -0.16 0.16 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.16 0.16 0.16 ;
END M1M2_PR_C

VIA M2M3_PR
  LAYER met2 ;
    RECT -0.14 -0.185 0.14 0.185 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR

VIA M2M3_PR_R
  LAYER met2 ;
    RECT -0.185 -0.14 0.185 0.14 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_R

VIA M2M3_PR_M
  LAYER met2 ;
    RECT -0.14 -0.185 0.14 0.185 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_M

VIA M2M3_PR_MR
  LAYER met2 ;
    RECT -0.185 -0.14 0.185 0.14 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_MR

VIA M2M3_PR_C
  LAYER met2 ;
    RECT -0.185 -0.185 0.185 0.185 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_C

VIA M3M4_PR
  LAYER met3 ;
    RECT -0.19 -0.16 0.19 0.16 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR

VIA M3M4_PR_R
  LAYER met3 ;
    RECT -0.16 -0.19 0.16 0.19 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_R

VIA M3M4_PR_M
  LAYER met3 ;
    RECT -0.19 -0.16 0.19 0.16 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_M

VIA M3M4_PR_MR
  LAYER met3 ;
    RECT -0.16 -0.19 0.16 0.19 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_MR

VIA M3M4_PR_C
  LAYER met3 ;
    RECT -0.19 -0.19 0.19 0.19 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_C

VIA M4M5_PR
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR

VIA M4M5_PR_R
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_R

VIA M4M5_PR_M
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_M

VIA M4M5_PR_MR
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_MR

VIA M4M5_PR_C
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_C

SITE unit
  CLASS CORE ;
  SYMMETRY Y ;
  SIZE 0.46 BY 2.72 ;
END unit

SITE unithddbl
  CLASS CORE ;
  SIZE 0.46 BY 5.44 ;
END unithddbl

MACRO cbx_1__1_
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  SIZE 77.28 BY 65.28 ;
  SYMMETRY X Y ;
  PIN prog_clk[0]
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER met2 ;
        RECT 2.23 63.92 2.37 65.28 ;
    END
  END prog_clk[0]
  PIN chanx_left_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 8.01 1.38 8.31 ;
    END
  END chanx_left_in[0]
  PIN chanx_left_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 16.85 1.38 17.15 ;
    END
  END chanx_left_in[1]
  PIN chanx_left_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 26.37 1.38 26.67 ;
    END
  END chanx_left_in[2]
  PIN chanx_left_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 36.57 1.38 36.87 ;
    END
  END chanx_left_in[3]
  PIN chanx_left_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 43.37 1.38 43.67 ;
    END
  END chanx_left_in[4]
  PIN chanx_left_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 48.13 1.38 48.43 ;
    END
  END chanx_left_in[5]
  PIN chanx_left_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 34.53 1.38 34.83 ;
    END
  END chanx_left_in[6]
  PIN chanx_left_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 42.01 1.38 42.31 ;
    END
  END chanx_left_in[7]
  PIN chanx_left_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 60.37 1.38 60.67 ;
    END
  END chanx_left_in[8]
  PIN chanx_left_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 54.93 1.38 55.23 ;
    END
  END chanx_left_in[9]
  PIN chanx_left_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 31.13 1.38 31.43 ;
    END
  END chanx_left_in[10]
  PIN chanx_left_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 33.17 1.38 33.47 ;
    END
  END chanx_left_in[11]
  PIN chanx_left_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 59.01 1.38 59.31 ;
    END
  END chanx_left_in[12]
  PIN chanx_left_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 61.73 1.38 62.03 ;
    END
  END chanx_left_in[13]
  PIN chanx_left_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 15.49 1.38 15.79 ;
    END
  END chanx_left_in[14]
  PIN chanx_left_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 56.29 1.38 56.59 ;
    END
  END chanx_left_in[15]
  PIN chanx_left_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 28.41 1.38 28.71 ;
    END
  END chanx_left_in[16]
  PIN chanx_left_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 22.29 1.38 22.59 ;
    END
  END chanx_left_in[17]
  PIN chanx_left_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 37.93 1.38 38.23 ;
    END
  END chanx_left_in[18]
  PIN chanx_left_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 49.49 1.38 49.79 ;
    END
  END chanx_left_in[19]
  PIN chanx_right_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 75.9 29.09 77.28 29.39 ;
    END
  END chanx_right_in[0]
  PIN chanx_right_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 75.9 40.65 77.28 40.95 ;
    END
  END chanx_right_in[1]
  PIN chanx_right_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 75.9 54.93 77.28 55.23 ;
    END
  END chanx_right_in[2]
  PIN chanx_right_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 75.9 11.41 77.28 11.71 ;
    END
  END chanx_right_in[3]
  PIN chanx_right_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 75.9 32.49 77.28 32.79 ;
    END
  END chanx_right_in[4]
  PIN chanx_right_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 75.9 30.45 77.28 30.75 ;
    END
  END chanx_right_in[5]
  PIN chanx_right_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 75.9 22.29 77.28 22.59 ;
    END
  END chanx_right_in[6]
  PIN chanx_right_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 75.9 37.93 77.28 38.23 ;
    END
  END chanx_right_in[7]
  PIN chanx_right_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 75.9 27.73 77.28 28.03 ;
    END
  END chanx_right_in[8]
  PIN chanx_right_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 75.9 16.85 77.28 17.15 ;
    END
  END chanx_right_in[9]
  PIN chanx_right_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 75.9 50.85 77.28 51.15 ;
    END
  END chanx_right_in[10]
  PIN chanx_right_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 75.9 33.85 77.28 34.15 ;
    END
  END chanx_right_in[11]
  PIN chanx_right_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 75.9 10.05 77.28 10.35 ;
    END
  END chanx_right_in[12]
  PIN chanx_right_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 75.9 4.61 77.28 4.91 ;
    END
  END chanx_right_in[13]
  PIN chanx_right_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 75.9 8.69 77.28 8.99 ;
    END
  END chanx_right_in[14]
  PIN chanx_right_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 75.9 23.65 77.28 23.95 ;
    END
  END chanx_right_in[15]
  PIN chanx_right_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 75.9 43.37 77.28 43.67 ;
    END
  END chanx_right_in[16]
  PIN chanx_right_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 75.9 20.93 77.28 21.23 ;
    END
  END chanx_right_in[17]
  PIN chanx_right_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 75.9 15.49 77.28 15.79 ;
    END
  END chanx_right_in[18]
  PIN chanx_right_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 75.9 52.21 77.28 52.51 ;
    END
  END chanx_right_in[19]
  PIN ccff_head[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 75.9 46.77 77.28 47.07 ;
    END
  END ccff_head[0]
  PIN chanx_left_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 18.21 1.38 18.51 ;
    END
  END chanx_left_out[0]
  PIN chanx_left_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 6.65 1.38 6.95 ;
    END
  END chanx_left_out[1]
  PIN chanx_left_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 29.77 1.38 30.07 ;
    END
  END chanx_left_out[2]
  PIN chanx_left_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 3.93 1.38 4.23 ;
    END
  END chanx_left_out[3]
  PIN chanx_left_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 52.21 1.38 52.51 ;
    END
  END chanx_left_out[4]
  PIN chanx_left_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 50.85 1.38 51.15 ;
    END
  END chanx_left_out[5]
  PIN chanx_left_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 23.65 1.38 23.95 ;
    END
  END chanx_left_out[6]
  PIN chanx_left_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 20.93 1.38 21.23 ;
    END
  END chanx_left_out[7]
  PIN chanx_left_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 25.01 1.38 25.31 ;
    END
  END chanx_left_out[8]
  PIN chanx_left_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 44.73 1.38 45.03 ;
    END
  END chanx_left_out[9]
  PIN chanx_left_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 5.29 1.38 5.59 ;
    END
  END chanx_left_out[10]
  PIN chanx_left_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 39.29 1.38 39.59 ;
    END
  END chanx_left_out[11]
  PIN chanx_left_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 46.09 1.38 46.39 ;
    END
  END chanx_left_out[12]
  PIN chanx_left_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 10.73 1.38 11.03 ;
    END
  END chanx_left_out[13]
  PIN chanx_left_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 9.37 1.38 9.67 ;
    END
  END chanx_left_out[14]
  PIN chanx_left_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 12.09 1.38 12.39 ;
    END
  END chanx_left_out[15]
  PIN chanx_left_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 53.57 1.38 53.87 ;
    END
  END chanx_left_out[16]
  PIN chanx_left_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 19.57 1.38 19.87 ;
    END
  END chanx_left_out[17]
  PIN chanx_left_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 40.65 1.38 40.95 ;
    END
  END chanx_left_out[18]
  PIN chanx_left_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 13.45 1.38 13.75 ;
    END
  END chanx_left_out[19]
  PIN chanx_right_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 75.9 35.21 77.28 35.51 ;
    END
  END chanx_right_out[0]
  PIN chanx_right_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 75.9 7.33 77.28 7.63 ;
    END
  END chanx_right_out[1]
  PIN chanx_right_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 75.9 26.37 77.28 26.67 ;
    END
  END chanx_right_out[2]
  PIN chanx_right_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 75.9 18.21 77.28 18.51 ;
    END
  END chanx_right_out[3]
  PIN chanx_right_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 75.9 19.57 77.28 19.87 ;
    END
  END chanx_right_out[4]
  PIN chanx_right_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 75.9 14.13 77.28 14.43 ;
    END
  END chanx_right_out[5]
  PIN chanx_right_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 75.9 5.97 77.28 6.27 ;
    END
  END chanx_right_out[6]
  PIN chanx_right_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 75.9 49.49 77.28 49.79 ;
    END
  END chanx_right_out[7]
  PIN chanx_right_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 75.9 53.57 77.28 53.87 ;
    END
  END chanx_right_out[8]
  PIN chanx_right_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 75.9 44.73 77.28 45.03 ;
    END
  END chanx_right_out[9]
  PIN chanx_right_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 75.9 25.01 77.28 25.31 ;
    END
  END chanx_right_out[10]
  PIN chanx_right_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 75.9 42.01 77.28 42.31 ;
    END
  END chanx_right_out[11]
  PIN chanx_right_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 75.9 48.13 77.28 48.43 ;
    END
  END chanx_right_out[12]
  PIN chanx_right_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 75.9 39.29 77.28 39.59 ;
    END
  END chanx_right_out[13]
  PIN chanx_right_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 75.9 61.05 77.28 61.35 ;
    END
  END chanx_right_out[14]
  PIN chanx_right_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 75.9 36.57 77.28 36.87 ;
    END
  END chanx_right_out[15]
  PIN chanx_right_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 75.9 56.97 77.28 57.27 ;
    END
  END chanx_right_out[16]
  PIN chanx_right_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 75.9 58.33 77.28 58.63 ;
    END
  END chanx_right_out[17]
  PIN chanx_right_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 75.9 59.69 77.28 59.99 ;
    END
  END chanx_right_out[18]
  PIN chanx_right_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 75.9 12.77 77.28 13.07 ;
    END
  END chanx_right_out[19]
  PIN bottom_grid_pin_0_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.01 0 45.15 1.36 ;
    END
  END bottom_grid_pin_0_[0]
  PIN bottom_grid_pin_1_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.71 0 19.85 1.36 ;
    END
  END bottom_grid_pin_1_[0]
  PIN bottom_grid_pin_2_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.53 0 4.67 1.36 ;
    END
  END bottom_grid_pin_2_[0]
  PIN bottom_grid_pin_3_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.47 0 22.61 1.36 ;
    END
  END bottom_grid_pin_3_[0]
  PIN bottom_grid_pin_4_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.33 0 41.47 1.36 ;
    END
  END bottom_grid_pin_4_[0]
  PIN bottom_grid_pin_5_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.25 0 42.39 1.36 ;
    END
  END bottom_grid_pin_5_[0]
  PIN bottom_grid_pin_6_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.41 0 40.55 1.36 ;
    END
  END bottom_grid_pin_6_[0]
  PIN bottom_grid_pin_7_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.31 0 24.45 1.36 ;
    END
  END bottom_grid_pin_7_[0]
  PIN bottom_grid_pin_8_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.17 0 43.31 1.36 ;
    END
  END bottom_grid_pin_8_[0]
  PIN bottom_grid_pin_9_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.89 0 58.03 1.36 ;
    END
  END bottom_grid_pin_9_[0]
  PIN bottom_grid_pin_10_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.09 0 44.23 1.36 ;
    END
  END bottom_grid_pin_10_[0]
  PIN bottom_grid_pin_11_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.81 0 58.95 1.36 ;
    END
  END bottom_grid_pin_11_[0]
  PIN bottom_grid_pin_12_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.39 0 23.53 1.36 ;
    END
  END bottom_grid_pin_12_[0]
  PIN bottom_grid_pin_13_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.87 0 18.01 1.36 ;
    END
  END bottom_grid_pin_13_[0]
  PIN bottom_grid_pin_14_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.79 0 18.93 1.36 ;
    END
  END bottom_grid_pin_14_[0]
  PIN bottom_grid_pin_15_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.95 0 17.09 1.36 ;
    END
  END bottom_grid_pin_15_[0]
  PIN ccff_tail[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 57.65 1.38 57.95 ;
    END
  END ccff_tail[0]
  PIN CLB_SC_IN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.81 63.92 58.95 65.28 ;
    END
  END CLB_SC_IN
  PIN CLB_SC_OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.55 0 21.69 1.36 ;
    END
  END CLB_SC_OUT
  PIN SC_IN_TOP
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.31 63.92 70.45 65.28 ;
    END
  END SC_IN_TOP
  PIN SC_IN_BOT
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.31 0 70.45 1.36 ;
    END
  END SC_IN_BOT
  PIN SC_OUT_TOP
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.55 63.92 21.69 65.28 ;
    END
  END SC_OUT_TOP
  PIN SC_OUT_BOT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.63 0 20.77 1.36 ;
    END
  END SC_OUT_BOT
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 23.62 0 24.22 0.6 ;
        RECT 53.06 0 53.66 0.6 ;
        RECT 23.62 64.68 24.22 65.28 ;
        RECT 53.06 64.68 53.66 65.28 ;
      LAYER met5 ;
        RECT 0 10.64 3.2 13.84 ;
        RECT 74.08 10.64 77.28 13.84 ;
        RECT 0 51.44 3.2 54.64 ;
        RECT 74.08 51.44 77.28 54.64 ;
      LAYER met1 ;
        RECT 0 2.48 0.48 2.96 ;
        RECT 76.8 2.48 77.28 2.96 ;
        RECT 0 7.92 0.48 8.4 ;
        RECT 76.8 7.92 77.28 8.4 ;
        RECT 0 13.36 0.48 13.84 ;
        RECT 76.8 13.36 77.28 13.84 ;
        RECT 0 18.8 0.48 19.28 ;
        RECT 76.8 18.8 77.28 19.28 ;
        RECT 0 24.24 0.48 24.72 ;
        RECT 76.8 24.24 77.28 24.72 ;
        RECT 0 29.68 0.48 30.16 ;
        RECT 76.8 29.68 77.28 30.16 ;
        RECT 0 35.12 0.48 35.6 ;
        RECT 76.8 35.12 77.28 35.6 ;
        RECT 0 40.56 0.48 41.04 ;
        RECT 76.8 40.56 77.28 41.04 ;
        RECT 0 46 0.48 46.48 ;
        RECT 76.8 46 77.28 46.48 ;
        RECT 0 51.44 0.48 51.92 ;
        RECT 76.8 51.44 77.28 51.92 ;
        RECT 0 56.88 0.48 57.36 ;
        RECT 76.8 56.88 77.28 57.36 ;
        RECT 0 62.32 0.48 62.8 ;
        RECT 76.8 62.32 77.28 62.8 ;
    END
  END VDD
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 8.9 0 9.5 0.6 ;
        RECT 38.34 0 38.94 0.6 ;
        RECT 67.78 0 68.38 0.6 ;
        RECT 8.9 64.68 9.5 65.28 ;
        RECT 38.34 64.68 38.94 65.28 ;
        RECT 67.78 64.68 68.38 65.28 ;
      LAYER met5 ;
        RECT 0 31.04 3.2 34.24 ;
        RECT 74.08 31.04 77.28 34.24 ;
      LAYER met1 ;
        RECT 0 0 77.28 0.24 ;
        RECT 0 5.2 0.48 5.68 ;
        RECT 76.8 5.2 77.28 5.68 ;
        RECT 0 10.64 0.48 11.12 ;
        RECT 76.8 10.64 77.28 11.12 ;
        RECT 0 16.08 0.48 16.56 ;
        RECT 76.8 16.08 77.28 16.56 ;
        RECT 0 21.52 0.48 22 ;
        RECT 76.8 21.52 77.28 22 ;
        RECT 0 26.96 0.48 27.44 ;
        RECT 76.8 26.96 77.28 27.44 ;
        RECT 0 32.4 0.48 32.88 ;
        RECT 76.8 32.4 77.28 32.88 ;
        RECT 0 37.84 0.48 38.32 ;
        RECT 76.8 37.84 77.28 38.32 ;
        RECT 0 43.28 0.48 43.76 ;
        RECT 76.8 43.28 77.28 43.76 ;
        RECT 0 48.72 0.48 49.2 ;
        RECT 76.8 48.72 77.28 49.2 ;
        RECT 0 54.16 0.48 54.64 ;
        RECT 76.8 54.16 77.28 54.64 ;
        RECT 0 59.6 0.48 60.08 ;
        RECT 76.8 59.6 77.28 60.08 ;
        RECT 0 65.04 77.28 65.28 ;
    END
  END VSS
  OBS
    LAYER li1 ;
      RECT 0 65.195 77.28 65.365 ;
      RECT 76.36 62.475 77.28 62.645 ;
      RECT 0 62.475 3.68 62.645 ;
      RECT 76.36 59.755 77.28 59.925 ;
      RECT 0 59.755 3.68 59.925 ;
      RECT 76.36 57.035 77.28 57.205 ;
      RECT 0 57.035 3.68 57.205 ;
      RECT 76.36 54.315 77.28 54.485 ;
      RECT 0 54.315 1.84 54.485 ;
      RECT 76.36 51.595 77.28 51.765 ;
      RECT 0 51.595 1.84 51.765 ;
      RECT 76.36 48.875 77.28 49.045 ;
      RECT 0 48.875 1.84 49.045 ;
      RECT 76.36 46.155 77.28 46.325 ;
      RECT 0 46.155 1.84 46.325 ;
      RECT 76.36 43.435 77.28 43.605 ;
      RECT 0 43.435 1.84 43.605 ;
      RECT 76.36 40.715 77.28 40.885 ;
      RECT 0 40.715 1.84 40.885 ;
      RECT 76.36 37.995 77.28 38.165 ;
      RECT 0 37.995 3.68 38.165 ;
      RECT 76.36 35.275 77.28 35.445 ;
      RECT 0 35.275 3.68 35.445 ;
      RECT 76.36 32.555 77.28 32.725 ;
      RECT 0 32.555 1.84 32.725 ;
      RECT 76.36 29.835 77.28 30.005 ;
      RECT 0 29.835 1.84 30.005 ;
      RECT 76.36 27.115 77.28 27.285 ;
      RECT 0 27.115 1.84 27.285 ;
      RECT 73.6 24.395 77.28 24.565 ;
      RECT 0 24.395 1.84 24.565 ;
      RECT 73.6 21.675 77.28 21.845 ;
      RECT 0 21.675 1.84 21.845 ;
      RECT 76.36 18.955 77.28 19.125 ;
      RECT 0 18.955 1.84 19.125 ;
      RECT 76.36 16.235 77.28 16.405 ;
      RECT 0 16.235 1.84 16.405 ;
      RECT 76.36 13.515 77.28 13.685 ;
      RECT 0 13.515 1.84 13.685 ;
      RECT 76.36 10.795 77.28 10.965 ;
      RECT 0 10.795 1.84 10.965 ;
      RECT 76.36 8.075 77.28 8.245 ;
      RECT 0 8.075 1.84 8.245 ;
      RECT 76.36 5.355 77.28 5.525 ;
      RECT 0 5.355 1.84 5.525 ;
      RECT 76.36 2.635 77.28 2.805 ;
      RECT 0 2.635 3.68 2.805 ;
      RECT 0 -0.085 77.28 0.085 ;
    LAYER met2 ;
      RECT 67.94 65.095 68.22 65.465 ;
      RECT 38.5 65.095 38.78 65.465 ;
      RECT 9.06 65.095 9.34 65.465 ;
      RECT 20.11 1.54 20.37 1.86 ;
      RECT 67.94 -0.185 68.22 0.185 ;
      RECT 38.5 -0.185 38.78 0.185 ;
      RECT 9.06 -0.185 9.34 0.185 ;
      POLYGON 77 65 77 0.28 70.73 0.28 70.73 1.64 70.03 1.64 70.03 0.28 59.23 0.28 59.23 1.64 58.53 1.64 58.53 0.28 58.31 0.28 58.31 1.64 57.61 1.64 57.61 0.28 45.43 0.28 45.43 1.64 44.73 1.64 44.73 0.28 44.51 0.28 44.51 1.64 43.81 1.64 43.81 0.28 43.59 0.28 43.59 1.64 42.89 1.64 42.89 0.28 42.67 0.28 42.67 1.64 41.97 1.64 41.97 0.28 41.75 0.28 41.75 1.64 41.05 1.64 41.05 0.28 40.83 0.28 40.83 1.64 40.13 1.64 40.13 0.28 24.73 0.28 24.73 1.64 24.03 1.64 24.03 0.28 23.81 0.28 23.81 1.64 23.11 1.64 23.11 0.28 22.89 0.28 22.89 1.64 22.19 1.64 22.19 0.28 21.97 0.28 21.97 1.64 21.27 1.64 21.27 0.28 21.05 0.28 21.05 1.64 20.35 1.64 20.35 0.28 20.13 0.28 20.13 1.64 19.43 1.64 19.43 0.28 19.21 0.28 19.21 1.64 18.51 1.64 18.51 0.28 18.29 0.28 18.29 1.64 17.59 1.64 17.59 0.28 17.37 0.28 17.37 1.64 16.67 1.64 16.67 0.28 4.95 0.28 4.95 1.64 4.25 1.64 4.25 0.28 0.28 0.28 0.28 65 1.95 65 1.95 63.64 2.65 63.64 2.65 65 21.27 65 21.27 63.64 21.97 63.64 21.97 65 58.53 65 58.53 63.64 59.23 63.64 59.23 65 70.03 65 70.03 63.64 70.73 63.64 70.73 65 ;
    LAYER met3 ;
      POLYGON 68.245 65.445 68.245 65.44 68.46 65.44 68.46 65.12 68.245 65.12 68.245 65.115 67.915 65.115 67.915 65.12 67.7 65.12 67.7 65.44 67.915 65.44 67.915 65.445 ;
      POLYGON 38.805 65.445 38.805 65.44 39.02 65.44 39.02 65.12 38.805 65.12 38.805 65.115 38.475 65.115 38.475 65.12 38.26 65.12 38.26 65.44 38.475 65.44 38.475 65.445 ;
      POLYGON 9.365 65.445 9.365 65.44 9.58 65.44 9.58 65.12 9.365 65.12 9.365 65.115 9.035 65.115 9.035 65.12 8.82 65.12 8.82 65.44 9.035 65.44 9.035 65.445 ;
      POLYGON 76.065 53.205 76.065 52.875 75.735 52.875 75.735 52.89 44.93 52.89 44.93 53.19 75.735 53.19 75.735 53.205 ;
      POLYGON 75.59 44.35 75.59 44.07 75.5 44.07 75.5 43.355 75.275 43.355 75.275 43.685 75.29 43.685 75.29 44.05 61.49 44.05 61.49 44.35 ;
      POLYGON 31.43 41.63 31.43 41.33 1.23 41.33 1.23 41.61 1.78 41.61 1.78 41.63 ;
      POLYGON 75.63 40.28 75.63 39.96 75.25 39.96 75.25 39.97 62.87 39.97 62.87 40.27 75.25 40.27 75.25 40.28 ;
      POLYGON 17.63 38.91 17.63 38.61 1.78 38.61 1.78 38.63 1.23 38.63 1.23 38.91 ;
      POLYGON 68.245 0.165 68.245 0.16 68.46 0.16 68.46 -0.16 68.245 -0.16 68.245 -0.165 67.915 -0.165 67.915 -0.16 67.7 -0.16 67.7 0.16 67.915 0.16 67.915 0.165 ;
      POLYGON 38.805 0.165 38.805 0.16 39.02 0.16 39.02 -0.16 38.805 -0.16 38.805 -0.165 38.475 -0.165 38.475 -0.16 38.26 -0.16 38.26 0.16 38.475 0.16 38.475 0.165 ;
      POLYGON 9.365 0.165 9.365 0.16 9.58 0.16 9.58 -0.16 9.365 -0.16 9.365 -0.165 9.035 -0.165 9.035 -0.16 8.82 -0.16 8.82 0.16 9.035 0.16 9.035 0.165 ;
      POLYGON 76.88 64.88 76.88 61.75 75.5 61.75 75.5 60.65 76.88 60.65 76.88 60.39 75.5 60.39 75.5 59.29 76.88 59.29 76.88 59.03 75.5 59.03 75.5 57.93 76.88 57.93 76.88 57.67 75.5 57.67 75.5 56.57 76.88 56.57 76.88 55.63 75.5 55.63 75.5 54.53 76.88 54.53 76.88 54.27 75.5 54.27 75.5 53.17 76.88 53.17 76.88 52.91 75.5 52.91 75.5 51.81 76.88 51.81 76.88 51.55 75.5 51.55 75.5 50.45 76.88 50.45 76.88 50.19 75.5 50.19 75.5 49.09 76.88 49.09 76.88 48.83 75.5 48.83 75.5 47.73 76.88 47.73 76.88 47.47 75.5 47.47 75.5 46.37 76.88 46.37 76.88 45.43 75.5 45.43 75.5 44.33 76.88 44.33 76.88 44.07 75.5 44.07 75.5 42.97 76.88 42.97 76.88 42.71 75.5 42.71 75.5 41.61 76.88 41.61 76.88 41.35 75.5 41.35 75.5 40.25 76.88 40.25 76.88 39.99 75.5 39.99 75.5 38.89 76.88 38.89 76.88 38.63 75.5 38.63 75.5 37.53 76.88 37.53 76.88 37.27 75.5 37.27 75.5 36.17 76.88 36.17 76.88 35.91 75.5 35.91 75.5 34.81 76.88 34.81 76.88 34.55 75.5 34.55 75.5 33.45 76.88 33.45 76.88 33.19 75.5 33.19 75.5 32.09 76.88 32.09 76.88 31.15 75.5 31.15 75.5 30.05 76.88 30.05 76.88 29.79 75.5 29.79 75.5 28.69 76.88 28.69 76.88 28.43 75.5 28.43 75.5 27.33 76.88 27.33 76.88 27.07 75.5 27.07 75.5 25.97 76.88 25.97 76.88 25.71 75.5 25.71 75.5 24.61 76.88 24.61 76.88 24.35 75.5 24.35 75.5 23.25 76.88 23.25 76.88 22.99 75.5 22.99 75.5 21.89 76.88 21.89 76.88 21.63 75.5 21.63 75.5 20.53 76.88 20.53 76.88 20.27 75.5 20.27 75.5 19.17 76.88 19.17 76.88 18.91 75.5 18.91 75.5 17.81 76.88 17.81 76.88 17.55 75.5 17.55 75.5 16.45 76.88 16.45 76.88 16.19 75.5 16.19 75.5 15.09 76.88 15.09 76.88 14.83 75.5 14.83 75.5 13.73 76.88 13.73 76.88 13.47 75.5 13.47 75.5 12.37 76.88 12.37 76.88 12.11 75.5 12.11 75.5 11.01 76.88 11.01 76.88 10.75 75.5 10.75 75.5 9.65 76.88 9.65 76.88 9.39 75.5 9.39 75.5 8.29 76.88 8.29 76.88 8.03 75.5 8.03 75.5 6.93 76.88 6.93 76.88 6.67 75.5 6.67 75.5 5.57 76.88 5.57 76.88 5.31 75.5 5.31 75.5 4.21 76.88 4.21 76.88 0.4 0.4 0.4 0.4 3.53 1.78 3.53 1.78 4.63 0.4 4.63 0.4 4.89 1.78 4.89 1.78 5.99 0.4 5.99 0.4 6.25 1.78 6.25 1.78 7.35 0.4 7.35 0.4 7.61 1.78 7.61 1.78 8.71 0.4 8.71 0.4 8.97 1.78 8.97 1.78 10.07 0.4 10.07 0.4 10.33 1.78 10.33 1.78 11.43 0.4 11.43 0.4 11.69 1.78 11.69 1.78 12.79 0.4 12.79 0.4 13.05 1.78 13.05 1.78 14.15 0.4 14.15 0.4 15.09 1.78 15.09 1.78 16.19 0.4 16.19 0.4 16.45 1.78 16.45 1.78 17.55 0.4 17.55 0.4 17.81 1.78 17.81 1.78 18.91 0.4 18.91 0.4 19.17 1.78 19.17 1.78 20.27 0.4 20.27 0.4 20.53 1.78 20.53 1.78 21.63 0.4 21.63 0.4 21.89 1.78 21.89 1.78 22.99 0.4 22.99 0.4 23.25 1.78 23.25 1.78 24.35 0.4 24.35 0.4 24.61 1.78 24.61 1.78 25.71 0.4 25.71 0.4 25.97 1.78 25.97 1.78 27.07 0.4 27.07 0.4 28.01 1.78 28.01 1.78 29.11 0.4 29.11 0.4 29.37 1.78 29.37 1.78 30.47 0.4 30.47 0.4 30.73 1.78 30.73 1.78 31.83 0.4 31.83 0.4 32.77 1.78 32.77 1.78 33.87 0.4 33.87 0.4 34.13 1.78 34.13 1.78 35.23 0.4 35.23 0.4 36.17 1.78 36.17 1.78 37.27 0.4 37.27 0.4 37.53 1.78 37.53 1.78 38.63 0.4 38.63 0.4 38.89 1.78 38.89 1.78 39.99 0.4 39.99 0.4 40.25 1.78 40.25 1.78 41.35 0.4 41.35 0.4 41.61 1.78 41.61 1.78 42.71 0.4 42.71 0.4 42.97 1.78 42.97 1.78 44.07 0.4 44.07 0.4 44.33 1.78 44.33 1.78 45.43 0.4 45.43 0.4 45.69 1.78 45.69 1.78 46.79 0.4 46.79 0.4 47.73 1.78 47.73 1.78 48.83 0.4 48.83 0.4 49.09 1.78 49.09 1.78 50.19 0.4 50.19 0.4 50.45 1.78 50.45 1.78 51.55 0.4 51.55 0.4 51.81 1.78 51.81 1.78 52.91 0.4 52.91 0.4 53.17 1.78 53.17 1.78 54.27 0.4 54.27 0.4 54.53 1.78 54.53 1.78 55.63 0.4 55.63 0.4 55.89 1.78 55.89 1.78 56.99 0.4 56.99 0.4 57.25 1.78 57.25 1.78 58.35 0.4 58.35 0.4 58.61 1.78 58.61 1.78 59.71 0.4 59.71 0.4 59.97 1.78 59.97 1.78 61.07 0.4 61.07 0.4 61.33 1.78 61.33 1.78 62.43 0.4 62.43 0.4 64.88 ;
    LAYER met1 ;
      POLYGON 77 64.76 77 63.08 76.52 63.08 76.52 62.04 77 62.04 77 60.36 76.52 60.36 76.52 59.32 77 59.32 77 57.64 76.52 57.64 76.52 56.6 77 56.6 77 54.92 76.52 54.92 76.52 53.88 77 53.88 77 52.2 76.52 52.2 76.52 51.16 77 51.16 77 49.48 76.52 49.48 76.52 48.44 77 48.44 77 46.76 76.52 46.76 76.52 45.72 77 45.72 77 44.04 76.52 44.04 76.52 43 77 43 77 41.32 76.52 41.32 76.52 40.28 77 40.28 77 38.6 76.52 38.6 76.52 37.56 77 37.56 77 35.88 76.52 35.88 76.52 34.84 77 34.84 77 33.16 76.52 33.16 76.52 32.12 77 32.12 77 30.44 76.52 30.44 76.52 29.4 77 29.4 77 27.72 76.52 27.72 76.52 26.68 77 26.68 77 25 76.52 25 76.52 23.96 77 23.96 77 22.28 76.52 22.28 76.52 21.24 77 21.24 77 19.56 76.52 19.56 76.52 18.52 77 18.52 77 16.84 76.52 16.84 76.52 15.8 77 15.8 77 14.12 76.52 14.12 76.52 13.08 77 13.08 77 11.4 76.52 11.4 76.52 10.36 77 10.36 77 8.68 76.52 8.68 76.52 7.64 77 7.64 77 5.96 76.52 5.96 76.52 4.92 77 4.92 77 3.24 76.52 3.24 76.52 2.2 77 2.2 77 0.52 0.28 0.52 0.28 2.2 0.76 2.2 0.76 3.24 0.28 3.24 0.28 4.92 0.76 4.92 0.76 5.96 0.28 5.96 0.28 7.64 0.76 7.64 0.76 8.68 0.28 8.68 0.28 10.36 0.76 10.36 0.76 11.4 0.28 11.4 0.28 13.08 0.76 13.08 0.76 14.12 0.28 14.12 0.28 15.8 0.76 15.8 0.76 16.84 0.28 16.84 0.28 18.52 0.76 18.52 0.76 19.56 0.28 19.56 0.28 21.24 0.76 21.24 0.76 22.28 0.28 22.28 0.28 23.96 0.76 23.96 0.76 25 0.28 25 0.28 26.68 0.76 26.68 0.76 27.72 0.28 27.72 0.28 29.4 0.76 29.4 0.76 30.44 0.28 30.44 0.28 32.12 0.76 32.12 0.76 33.16 0.28 33.16 0.28 34.84 0.76 34.84 0.76 35.88 0.28 35.88 0.28 37.56 0.76 37.56 0.76 38.6 0.28 38.6 0.28 40.28 0.76 40.28 0.76 41.32 0.28 41.32 0.28 43 0.76 43 0.76 44.04 0.28 44.04 0.28 45.72 0.76 45.72 0.76 46.76 0.28 46.76 0.28 48.44 0.76 48.44 0.76 49.48 0.28 49.48 0.28 51.16 0.76 51.16 0.76 52.2 0.28 52.2 0.28 53.88 0.76 53.88 0.76 54.92 0.28 54.92 0.28 56.6 0.76 56.6 0.76 57.64 0.28 57.64 0.28 59.32 0.76 59.32 0.76 60.36 0.28 60.36 0.28 62.04 0.76 62.04 0.76 63.08 0.28 63.08 0.28 64.76 ;
    LAYER met5 ;
      POLYGON 75.68 63.68 75.68 56.24 72.48 56.24 72.48 49.84 75.68 49.84 75.68 35.84 72.48 35.84 72.48 29.44 75.68 29.44 75.68 15.44 72.48 15.44 72.48 9.04 75.68 9.04 75.68 1.6 1.6 1.6 1.6 9.04 4.8 9.04 4.8 15.44 1.6 15.44 1.6 29.44 4.8 29.44 4.8 35.84 1.6 35.84 1.6 49.84 4.8 49.84 4.8 56.24 1.6 56.24 1.6 63.68 ;
    LAYER met4 ;
      POLYGON 76.88 64.88 76.88 0.4 68.78 0.4 68.78 1 67.38 1 67.38 0.4 54.06 0.4 54.06 1 52.66 1 52.66 0.4 39.34 0.4 39.34 1 37.94 1 37.94 0.4 24.62 0.4 24.62 1 23.22 1 23.22 0.4 9.9 0.4 9.9 1 8.5 1 8.5 0.4 0.4 0.4 0.4 64.88 8.5 64.88 8.5 64.28 9.9 64.28 9.9 64.88 23.22 64.88 23.22 64.28 24.62 64.28 24.62 64.88 37.94 64.88 37.94 64.28 39.34 64.28 39.34 64.88 52.66 64.88 52.66 64.28 54.06 64.28 54.06 64.88 67.38 64.88 67.38 64.28 68.78 64.28 68.78 64.88 ;
    LAYER li1 ;
      RECT 0.17 0.17 77.11 65.11 ;
    LAYER mcon ;
      RECT 76.965 65.195 77.135 65.365 ;
      RECT 76.505 65.195 76.675 65.365 ;
      RECT 76.045 65.195 76.215 65.365 ;
      RECT 75.585 65.195 75.755 65.365 ;
      RECT 75.125 65.195 75.295 65.365 ;
      RECT 74.665 65.195 74.835 65.365 ;
      RECT 74.205 65.195 74.375 65.365 ;
      RECT 73.745 65.195 73.915 65.365 ;
      RECT 73.285 65.195 73.455 65.365 ;
      RECT 72.825 65.195 72.995 65.365 ;
      RECT 72.365 65.195 72.535 65.365 ;
      RECT 71.905 65.195 72.075 65.365 ;
      RECT 71.445 65.195 71.615 65.365 ;
      RECT 70.985 65.195 71.155 65.365 ;
      RECT 70.525 65.195 70.695 65.365 ;
      RECT 70.065 65.195 70.235 65.365 ;
      RECT 69.605 65.195 69.775 65.365 ;
      RECT 69.145 65.195 69.315 65.365 ;
      RECT 68.685 65.195 68.855 65.365 ;
      RECT 68.225 65.195 68.395 65.365 ;
      RECT 67.765 65.195 67.935 65.365 ;
      RECT 67.305 65.195 67.475 65.365 ;
      RECT 66.845 65.195 67.015 65.365 ;
      RECT 66.385 65.195 66.555 65.365 ;
      RECT 65.925 65.195 66.095 65.365 ;
      RECT 65.465 65.195 65.635 65.365 ;
      RECT 65.005 65.195 65.175 65.365 ;
      RECT 64.545 65.195 64.715 65.365 ;
      RECT 64.085 65.195 64.255 65.365 ;
      RECT 63.625 65.195 63.795 65.365 ;
      RECT 63.165 65.195 63.335 65.365 ;
      RECT 62.705 65.195 62.875 65.365 ;
      RECT 62.245 65.195 62.415 65.365 ;
      RECT 61.785 65.195 61.955 65.365 ;
      RECT 61.325 65.195 61.495 65.365 ;
      RECT 60.865 65.195 61.035 65.365 ;
      RECT 60.405 65.195 60.575 65.365 ;
      RECT 59.945 65.195 60.115 65.365 ;
      RECT 59.485 65.195 59.655 65.365 ;
      RECT 59.025 65.195 59.195 65.365 ;
      RECT 58.565 65.195 58.735 65.365 ;
      RECT 58.105 65.195 58.275 65.365 ;
      RECT 57.645 65.195 57.815 65.365 ;
      RECT 57.185 65.195 57.355 65.365 ;
      RECT 56.725 65.195 56.895 65.365 ;
      RECT 56.265 65.195 56.435 65.365 ;
      RECT 55.805 65.195 55.975 65.365 ;
      RECT 55.345 65.195 55.515 65.365 ;
      RECT 54.885 65.195 55.055 65.365 ;
      RECT 54.425 65.195 54.595 65.365 ;
      RECT 53.965 65.195 54.135 65.365 ;
      RECT 53.505 65.195 53.675 65.365 ;
      RECT 53.045 65.195 53.215 65.365 ;
      RECT 52.585 65.195 52.755 65.365 ;
      RECT 52.125 65.195 52.295 65.365 ;
      RECT 51.665 65.195 51.835 65.365 ;
      RECT 51.205 65.195 51.375 65.365 ;
      RECT 50.745 65.195 50.915 65.365 ;
      RECT 50.285 65.195 50.455 65.365 ;
      RECT 49.825 65.195 49.995 65.365 ;
      RECT 49.365 65.195 49.535 65.365 ;
      RECT 48.905 65.195 49.075 65.365 ;
      RECT 48.445 65.195 48.615 65.365 ;
      RECT 47.985 65.195 48.155 65.365 ;
      RECT 47.525 65.195 47.695 65.365 ;
      RECT 47.065 65.195 47.235 65.365 ;
      RECT 46.605 65.195 46.775 65.365 ;
      RECT 46.145 65.195 46.315 65.365 ;
      RECT 45.685 65.195 45.855 65.365 ;
      RECT 45.225 65.195 45.395 65.365 ;
      RECT 44.765 65.195 44.935 65.365 ;
      RECT 44.305 65.195 44.475 65.365 ;
      RECT 43.845 65.195 44.015 65.365 ;
      RECT 43.385 65.195 43.555 65.365 ;
      RECT 42.925 65.195 43.095 65.365 ;
      RECT 42.465 65.195 42.635 65.365 ;
      RECT 42.005 65.195 42.175 65.365 ;
      RECT 41.545 65.195 41.715 65.365 ;
      RECT 41.085 65.195 41.255 65.365 ;
      RECT 40.625 65.195 40.795 65.365 ;
      RECT 40.165 65.195 40.335 65.365 ;
      RECT 39.705 65.195 39.875 65.365 ;
      RECT 39.245 65.195 39.415 65.365 ;
      RECT 38.785 65.195 38.955 65.365 ;
      RECT 38.325 65.195 38.495 65.365 ;
      RECT 37.865 65.195 38.035 65.365 ;
      RECT 37.405 65.195 37.575 65.365 ;
      RECT 36.945 65.195 37.115 65.365 ;
      RECT 36.485 65.195 36.655 65.365 ;
      RECT 36.025 65.195 36.195 65.365 ;
      RECT 35.565 65.195 35.735 65.365 ;
      RECT 35.105 65.195 35.275 65.365 ;
      RECT 34.645 65.195 34.815 65.365 ;
      RECT 34.185 65.195 34.355 65.365 ;
      RECT 33.725 65.195 33.895 65.365 ;
      RECT 33.265 65.195 33.435 65.365 ;
      RECT 32.805 65.195 32.975 65.365 ;
      RECT 32.345 65.195 32.515 65.365 ;
      RECT 31.885 65.195 32.055 65.365 ;
      RECT 31.425 65.195 31.595 65.365 ;
      RECT 30.965 65.195 31.135 65.365 ;
      RECT 30.505 65.195 30.675 65.365 ;
      RECT 30.045 65.195 30.215 65.365 ;
      RECT 29.585 65.195 29.755 65.365 ;
      RECT 29.125 65.195 29.295 65.365 ;
      RECT 28.665 65.195 28.835 65.365 ;
      RECT 28.205 65.195 28.375 65.365 ;
      RECT 27.745 65.195 27.915 65.365 ;
      RECT 27.285 65.195 27.455 65.365 ;
      RECT 26.825 65.195 26.995 65.365 ;
      RECT 26.365 65.195 26.535 65.365 ;
      RECT 25.905 65.195 26.075 65.365 ;
      RECT 25.445 65.195 25.615 65.365 ;
      RECT 24.985 65.195 25.155 65.365 ;
      RECT 24.525 65.195 24.695 65.365 ;
      RECT 24.065 65.195 24.235 65.365 ;
      RECT 23.605 65.195 23.775 65.365 ;
      RECT 23.145 65.195 23.315 65.365 ;
      RECT 22.685 65.195 22.855 65.365 ;
      RECT 22.225 65.195 22.395 65.365 ;
      RECT 21.765 65.195 21.935 65.365 ;
      RECT 21.305 65.195 21.475 65.365 ;
      RECT 20.845 65.195 21.015 65.365 ;
      RECT 20.385 65.195 20.555 65.365 ;
      RECT 19.925 65.195 20.095 65.365 ;
      RECT 19.465 65.195 19.635 65.365 ;
      RECT 19.005 65.195 19.175 65.365 ;
      RECT 18.545 65.195 18.715 65.365 ;
      RECT 18.085 65.195 18.255 65.365 ;
      RECT 17.625 65.195 17.795 65.365 ;
      RECT 17.165 65.195 17.335 65.365 ;
      RECT 16.705 65.195 16.875 65.365 ;
      RECT 16.245 65.195 16.415 65.365 ;
      RECT 15.785 65.195 15.955 65.365 ;
      RECT 15.325 65.195 15.495 65.365 ;
      RECT 14.865 65.195 15.035 65.365 ;
      RECT 14.405 65.195 14.575 65.365 ;
      RECT 13.945 65.195 14.115 65.365 ;
      RECT 13.485 65.195 13.655 65.365 ;
      RECT 13.025 65.195 13.195 65.365 ;
      RECT 12.565 65.195 12.735 65.365 ;
      RECT 12.105 65.195 12.275 65.365 ;
      RECT 11.645 65.195 11.815 65.365 ;
      RECT 11.185 65.195 11.355 65.365 ;
      RECT 10.725 65.195 10.895 65.365 ;
      RECT 10.265 65.195 10.435 65.365 ;
      RECT 9.805 65.195 9.975 65.365 ;
      RECT 9.345 65.195 9.515 65.365 ;
      RECT 8.885 65.195 9.055 65.365 ;
      RECT 8.425 65.195 8.595 65.365 ;
      RECT 7.965 65.195 8.135 65.365 ;
      RECT 7.505 65.195 7.675 65.365 ;
      RECT 7.045 65.195 7.215 65.365 ;
      RECT 6.585 65.195 6.755 65.365 ;
      RECT 6.125 65.195 6.295 65.365 ;
      RECT 5.665 65.195 5.835 65.365 ;
      RECT 5.205 65.195 5.375 65.365 ;
      RECT 4.745 65.195 4.915 65.365 ;
      RECT 4.285 65.195 4.455 65.365 ;
      RECT 3.825 65.195 3.995 65.365 ;
      RECT 3.365 65.195 3.535 65.365 ;
      RECT 2.905 65.195 3.075 65.365 ;
      RECT 2.445 65.195 2.615 65.365 ;
      RECT 1.985 65.195 2.155 65.365 ;
      RECT 1.525 65.195 1.695 65.365 ;
      RECT 1.065 65.195 1.235 65.365 ;
      RECT 0.605 65.195 0.775 65.365 ;
      RECT 0.145 65.195 0.315 65.365 ;
      RECT 76.965 62.475 77.135 62.645 ;
      RECT 76.505 62.475 76.675 62.645 ;
      RECT 0.605 62.475 0.775 62.645 ;
      RECT 0.145 62.475 0.315 62.645 ;
      RECT 76.965 59.755 77.135 59.925 ;
      RECT 76.505 59.755 76.675 59.925 ;
      RECT 0.605 59.755 0.775 59.925 ;
      RECT 0.145 59.755 0.315 59.925 ;
      RECT 76.965 57.035 77.135 57.205 ;
      RECT 76.505 57.035 76.675 57.205 ;
      RECT 0.605 57.035 0.775 57.205 ;
      RECT 0.145 57.035 0.315 57.205 ;
      RECT 76.965 54.315 77.135 54.485 ;
      RECT 76.505 54.315 76.675 54.485 ;
      RECT 0.605 54.315 0.775 54.485 ;
      RECT 0.145 54.315 0.315 54.485 ;
      RECT 76.965 51.595 77.135 51.765 ;
      RECT 76.505 51.595 76.675 51.765 ;
      RECT 0.605 51.595 0.775 51.765 ;
      RECT 0.145 51.595 0.315 51.765 ;
      RECT 76.965 48.875 77.135 49.045 ;
      RECT 76.505 48.875 76.675 49.045 ;
      RECT 0.605 48.875 0.775 49.045 ;
      RECT 0.145 48.875 0.315 49.045 ;
      RECT 76.965 46.155 77.135 46.325 ;
      RECT 76.505 46.155 76.675 46.325 ;
      RECT 0.605 46.155 0.775 46.325 ;
      RECT 0.145 46.155 0.315 46.325 ;
      RECT 76.965 43.435 77.135 43.605 ;
      RECT 76.505 43.435 76.675 43.605 ;
      RECT 0.605 43.435 0.775 43.605 ;
      RECT 0.145 43.435 0.315 43.605 ;
      RECT 76.965 40.715 77.135 40.885 ;
      RECT 76.505 40.715 76.675 40.885 ;
      RECT 0.605 40.715 0.775 40.885 ;
      RECT 0.145 40.715 0.315 40.885 ;
      RECT 76.965 37.995 77.135 38.165 ;
      RECT 76.505 37.995 76.675 38.165 ;
      RECT 0.605 37.995 0.775 38.165 ;
      RECT 0.145 37.995 0.315 38.165 ;
      RECT 76.965 35.275 77.135 35.445 ;
      RECT 76.505 35.275 76.675 35.445 ;
      RECT 0.605 35.275 0.775 35.445 ;
      RECT 0.145 35.275 0.315 35.445 ;
      RECT 76.965 32.555 77.135 32.725 ;
      RECT 76.505 32.555 76.675 32.725 ;
      RECT 0.605 32.555 0.775 32.725 ;
      RECT 0.145 32.555 0.315 32.725 ;
      RECT 76.965 29.835 77.135 30.005 ;
      RECT 76.505 29.835 76.675 30.005 ;
      RECT 0.605 29.835 0.775 30.005 ;
      RECT 0.145 29.835 0.315 30.005 ;
      RECT 76.965 27.115 77.135 27.285 ;
      RECT 76.505 27.115 76.675 27.285 ;
      RECT 0.605 27.115 0.775 27.285 ;
      RECT 0.145 27.115 0.315 27.285 ;
      RECT 76.965 24.395 77.135 24.565 ;
      RECT 76.505 24.395 76.675 24.565 ;
      RECT 0.605 24.395 0.775 24.565 ;
      RECT 0.145 24.395 0.315 24.565 ;
      RECT 76.965 21.675 77.135 21.845 ;
      RECT 76.505 21.675 76.675 21.845 ;
      RECT 0.605 21.675 0.775 21.845 ;
      RECT 0.145 21.675 0.315 21.845 ;
      RECT 76.965 18.955 77.135 19.125 ;
      RECT 76.505 18.955 76.675 19.125 ;
      RECT 0.605 18.955 0.775 19.125 ;
      RECT 0.145 18.955 0.315 19.125 ;
      RECT 76.965 16.235 77.135 16.405 ;
      RECT 76.505 16.235 76.675 16.405 ;
      RECT 0.605 16.235 0.775 16.405 ;
      RECT 0.145 16.235 0.315 16.405 ;
      RECT 76.965 13.515 77.135 13.685 ;
      RECT 76.505 13.515 76.675 13.685 ;
      RECT 0.605 13.515 0.775 13.685 ;
      RECT 0.145 13.515 0.315 13.685 ;
      RECT 76.965 10.795 77.135 10.965 ;
      RECT 76.505 10.795 76.675 10.965 ;
      RECT 0.605 10.795 0.775 10.965 ;
      RECT 0.145 10.795 0.315 10.965 ;
      RECT 76.965 8.075 77.135 8.245 ;
      RECT 76.505 8.075 76.675 8.245 ;
      RECT 0.605 8.075 0.775 8.245 ;
      RECT 0.145 8.075 0.315 8.245 ;
      RECT 76.965 5.355 77.135 5.525 ;
      RECT 76.505 5.355 76.675 5.525 ;
      RECT 0.605 5.355 0.775 5.525 ;
      RECT 0.145 5.355 0.315 5.525 ;
      RECT 76.965 2.635 77.135 2.805 ;
      RECT 76.505 2.635 76.675 2.805 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 76.965 -0.085 77.135 0.085 ;
      RECT 76.505 -0.085 76.675 0.085 ;
      RECT 76.045 -0.085 76.215 0.085 ;
      RECT 75.585 -0.085 75.755 0.085 ;
      RECT 75.125 -0.085 75.295 0.085 ;
      RECT 74.665 -0.085 74.835 0.085 ;
      RECT 74.205 -0.085 74.375 0.085 ;
      RECT 73.745 -0.085 73.915 0.085 ;
      RECT 73.285 -0.085 73.455 0.085 ;
      RECT 72.825 -0.085 72.995 0.085 ;
      RECT 72.365 -0.085 72.535 0.085 ;
      RECT 71.905 -0.085 72.075 0.085 ;
      RECT 71.445 -0.085 71.615 0.085 ;
      RECT 70.985 -0.085 71.155 0.085 ;
      RECT 70.525 -0.085 70.695 0.085 ;
      RECT 70.065 -0.085 70.235 0.085 ;
      RECT 69.605 -0.085 69.775 0.085 ;
      RECT 69.145 -0.085 69.315 0.085 ;
      RECT 68.685 -0.085 68.855 0.085 ;
      RECT 68.225 -0.085 68.395 0.085 ;
      RECT 67.765 -0.085 67.935 0.085 ;
      RECT 67.305 -0.085 67.475 0.085 ;
      RECT 66.845 -0.085 67.015 0.085 ;
      RECT 66.385 -0.085 66.555 0.085 ;
      RECT 65.925 -0.085 66.095 0.085 ;
      RECT 65.465 -0.085 65.635 0.085 ;
      RECT 65.005 -0.085 65.175 0.085 ;
      RECT 64.545 -0.085 64.715 0.085 ;
      RECT 64.085 -0.085 64.255 0.085 ;
      RECT 63.625 -0.085 63.795 0.085 ;
      RECT 63.165 -0.085 63.335 0.085 ;
      RECT 62.705 -0.085 62.875 0.085 ;
      RECT 62.245 -0.085 62.415 0.085 ;
      RECT 61.785 -0.085 61.955 0.085 ;
      RECT 61.325 -0.085 61.495 0.085 ;
      RECT 60.865 -0.085 61.035 0.085 ;
      RECT 60.405 -0.085 60.575 0.085 ;
      RECT 59.945 -0.085 60.115 0.085 ;
      RECT 59.485 -0.085 59.655 0.085 ;
      RECT 59.025 -0.085 59.195 0.085 ;
      RECT 58.565 -0.085 58.735 0.085 ;
      RECT 58.105 -0.085 58.275 0.085 ;
      RECT 57.645 -0.085 57.815 0.085 ;
      RECT 57.185 -0.085 57.355 0.085 ;
      RECT 56.725 -0.085 56.895 0.085 ;
      RECT 56.265 -0.085 56.435 0.085 ;
      RECT 55.805 -0.085 55.975 0.085 ;
      RECT 55.345 -0.085 55.515 0.085 ;
      RECT 54.885 -0.085 55.055 0.085 ;
      RECT 54.425 -0.085 54.595 0.085 ;
      RECT 53.965 -0.085 54.135 0.085 ;
      RECT 53.505 -0.085 53.675 0.085 ;
      RECT 53.045 -0.085 53.215 0.085 ;
      RECT 52.585 -0.085 52.755 0.085 ;
      RECT 52.125 -0.085 52.295 0.085 ;
      RECT 51.665 -0.085 51.835 0.085 ;
      RECT 51.205 -0.085 51.375 0.085 ;
      RECT 50.745 -0.085 50.915 0.085 ;
      RECT 50.285 -0.085 50.455 0.085 ;
      RECT 49.825 -0.085 49.995 0.085 ;
      RECT 49.365 -0.085 49.535 0.085 ;
      RECT 48.905 -0.085 49.075 0.085 ;
      RECT 48.445 -0.085 48.615 0.085 ;
      RECT 47.985 -0.085 48.155 0.085 ;
      RECT 47.525 -0.085 47.695 0.085 ;
      RECT 47.065 -0.085 47.235 0.085 ;
      RECT 46.605 -0.085 46.775 0.085 ;
      RECT 46.145 -0.085 46.315 0.085 ;
      RECT 45.685 -0.085 45.855 0.085 ;
      RECT 45.225 -0.085 45.395 0.085 ;
      RECT 44.765 -0.085 44.935 0.085 ;
      RECT 44.305 -0.085 44.475 0.085 ;
      RECT 43.845 -0.085 44.015 0.085 ;
      RECT 43.385 -0.085 43.555 0.085 ;
      RECT 42.925 -0.085 43.095 0.085 ;
      RECT 42.465 -0.085 42.635 0.085 ;
      RECT 42.005 -0.085 42.175 0.085 ;
      RECT 41.545 -0.085 41.715 0.085 ;
      RECT 41.085 -0.085 41.255 0.085 ;
      RECT 40.625 -0.085 40.795 0.085 ;
      RECT 40.165 -0.085 40.335 0.085 ;
      RECT 39.705 -0.085 39.875 0.085 ;
      RECT 39.245 -0.085 39.415 0.085 ;
      RECT 38.785 -0.085 38.955 0.085 ;
      RECT 38.325 -0.085 38.495 0.085 ;
      RECT 37.865 -0.085 38.035 0.085 ;
      RECT 37.405 -0.085 37.575 0.085 ;
      RECT 36.945 -0.085 37.115 0.085 ;
      RECT 36.485 -0.085 36.655 0.085 ;
      RECT 36.025 -0.085 36.195 0.085 ;
      RECT 35.565 -0.085 35.735 0.085 ;
      RECT 35.105 -0.085 35.275 0.085 ;
      RECT 34.645 -0.085 34.815 0.085 ;
      RECT 34.185 -0.085 34.355 0.085 ;
      RECT 33.725 -0.085 33.895 0.085 ;
      RECT 33.265 -0.085 33.435 0.085 ;
      RECT 32.805 -0.085 32.975 0.085 ;
      RECT 32.345 -0.085 32.515 0.085 ;
      RECT 31.885 -0.085 32.055 0.085 ;
      RECT 31.425 -0.085 31.595 0.085 ;
      RECT 30.965 -0.085 31.135 0.085 ;
      RECT 30.505 -0.085 30.675 0.085 ;
      RECT 30.045 -0.085 30.215 0.085 ;
      RECT 29.585 -0.085 29.755 0.085 ;
      RECT 29.125 -0.085 29.295 0.085 ;
      RECT 28.665 -0.085 28.835 0.085 ;
      RECT 28.205 -0.085 28.375 0.085 ;
      RECT 27.745 -0.085 27.915 0.085 ;
      RECT 27.285 -0.085 27.455 0.085 ;
      RECT 26.825 -0.085 26.995 0.085 ;
      RECT 26.365 -0.085 26.535 0.085 ;
      RECT 25.905 -0.085 26.075 0.085 ;
      RECT 25.445 -0.085 25.615 0.085 ;
      RECT 24.985 -0.085 25.155 0.085 ;
      RECT 24.525 -0.085 24.695 0.085 ;
      RECT 24.065 -0.085 24.235 0.085 ;
      RECT 23.605 -0.085 23.775 0.085 ;
      RECT 23.145 -0.085 23.315 0.085 ;
      RECT 22.685 -0.085 22.855 0.085 ;
      RECT 22.225 -0.085 22.395 0.085 ;
      RECT 21.765 -0.085 21.935 0.085 ;
      RECT 21.305 -0.085 21.475 0.085 ;
      RECT 20.845 -0.085 21.015 0.085 ;
      RECT 20.385 -0.085 20.555 0.085 ;
      RECT 19.925 -0.085 20.095 0.085 ;
      RECT 19.465 -0.085 19.635 0.085 ;
      RECT 19.005 -0.085 19.175 0.085 ;
      RECT 18.545 -0.085 18.715 0.085 ;
      RECT 18.085 -0.085 18.255 0.085 ;
      RECT 17.625 -0.085 17.795 0.085 ;
      RECT 17.165 -0.085 17.335 0.085 ;
      RECT 16.705 -0.085 16.875 0.085 ;
      RECT 16.245 -0.085 16.415 0.085 ;
      RECT 15.785 -0.085 15.955 0.085 ;
      RECT 15.325 -0.085 15.495 0.085 ;
      RECT 14.865 -0.085 15.035 0.085 ;
      RECT 14.405 -0.085 14.575 0.085 ;
      RECT 13.945 -0.085 14.115 0.085 ;
      RECT 13.485 -0.085 13.655 0.085 ;
      RECT 13.025 -0.085 13.195 0.085 ;
      RECT 12.565 -0.085 12.735 0.085 ;
      RECT 12.105 -0.085 12.275 0.085 ;
      RECT 11.645 -0.085 11.815 0.085 ;
      RECT 11.185 -0.085 11.355 0.085 ;
      RECT 10.725 -0.085 10.895 0.085 ;
      RECT 10.265 -0.085 10.435 0.085 ;
      RECT 9.805 -0.085 9.975 0.085 ;
      RECT 9.345 -0.085 9.515 0.085 ;
      RECT 8.885 -0.085 9.055 0.085 ;
      RECT 8.425 -0.085 8.595 0.085 ;
      RECT 7.965 -0.085 8.135 0.085 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.145 -0.085 0.315 0.085 ;
    LAYER via ;
      RECT 68.005 65.205 68.155 65.355 ;
      RECT 38.565 65.205 38.715 65.355 ;
      RECT 9.125 65.205 9.275 65.355 ;
      RECT 23.385 1.625 23.535 1.775 ;
      RECT 22.465 1.625 22.615 1.775 ;
      RECT 68.005 -0.075 68.155 0.075 ;
      RECT 38.565 -0.075 38.715 0.075 ;
      RECT 9.125 -0.075 9.275 0.075 ;
    LAYER via2 ;
      RECT 67.98 65.18 68.18 65.38 ;
      RECT 38.54 65.18 38.74 65.38 ;
      RECT 9.1 65.18 9.3 65.38 ;
      RECT 1.74 57.7 1.94 57.9 ;
      RECT 1.74 53.62 1.94 53.82 ;
      RECT 75.34 43.42 75.54 43.62 ;
      RECT 75.8 39.34 76 39.54 ;
      RECT 1.28 39.34 1.48 39.54 ;
      RECT 75.34 36.62 75.54 36.82 ;
      RECT 75.8 33.9 76 34.1 ;
      RECT 1.74 23.7 1.94 23.9 ;
      RECT 75.34 14.18 75.54 14.38 ;
      RECT 1.74 6.7 1.94 6.9 ;
      RECT 75.8 6.02 76 6.22 ;
      RECT 1.28 3.98 1.48 4.18 ;
      RECT 67.98 -0.1 68.18 0.1 ;
      RECT 38.54 -0.1 38.74 0.1 ;
      RECT 9.1 -0.1 9.3 0.1 ;
    LAYER via3 ;
      RECT 67.98 65.18 68.18 65.38 ;
      RECT 38.54 65.18 38.74 65.38 ;
      RECT 9.1 65.18 9.3 65.38 ;
      RECT 75.34 10.1 75.54 10.3 ;
      RECT 67.98 -0.1 68.18 0.1 ;
      RECT 38.54 -0.1 38.74 0.1 ;
      RECT 9.1 -0.1 9.3 0.1 ;
    LAYER OVERLAP ;
      POLYGON 0 0 0 65.28 77.28 65.28 77.28 0 ;
  END
END cbx_1__1_

END LIBRARY
