VERSION 5.7 ;
BUSBITCHARS "[]" ;

UNITS
  DATABASE MICRONS 1000 ;
END UNITS

MANUFACTURINGGRID 0.005 ;

LAYER li1
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.46 ;
  WIDTH 0.17 ;
END li1

LAYER mcon
  TYPE CUT ;
END mcon

LAYER met1
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.34 ;
  WIDTH 0.14 ;
END met1

LAYER via
  TYPE CUT ;
END via

LAYER met2
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.46 ;
  WIDTH 0.14 ;
END met2

LAYER via2
  TYPE CUT ;
END via2

LAYER met3
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.68 ;
  WIDTH 0.3 ;
END met3

LAYER via3
  TYPE CUT ;
END via3

LAYER met4
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.92 ;
  WIDTH 0.3 ;
END met4

LAYER via4
  TYPE CUT ;
END via4

LAYER met5
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 3.4 ;
  WIDTH 1.6 ;
END met5

LAYER nwell
  TYPE MASTERSLICE ;
END nwell

LAYER pwell
  TYPE MASTERSLICE ;
END pwell

LAYER OVERLAP
  TYPE OVERLAP ;
END OVERLAP

VIA L1M1_PR
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.145 -0.115 0.145 0.115 ;
END L1M1_PR

VIA L1M1_PR_R
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.115 -0.145 0.115 0.145 ;
END L1M1_PR_R

VIA L1M1_PR_M
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.115 -0.145 0.115 0.145 ;
END L1M1_PR_M

VIA L1M1_PR_MR
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.145 -0.115 0.145 0.115 ;
END L1M1_PR_MR

VIA L1M1_PR_C
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.145 -0.145 0.145 0.145 ;
END L1M1_PR_C

VIA M1M2_PR
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR

VIA M1M2_PR_Enc
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_Enc

VIA M1M2_PR_R
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_R

VIA M1M2_PR_R_Enc
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR_R_Enc

VIA M1M2_PR_M
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_M

VIA M1M2_PR_M_Enc
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR_M_Enc

VIA M1M2_PR_MR
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR_MR

VIA M1M2_PR_MR_Enc
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_MR_Enc

VIA M1M2_PR_C
  LAYER met1 ;
    RECT -0.16 -0.16 0.16 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.16 0.16 0.16 ;
END M1M2_PR_C

VIA M2M3_PR
  LAYER met2 ;
    RECT -0.14 -0.185 0.14 0.185 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR

VIA M2M3_PR_R
  LAYER met2 ;
    RECT -0.185 -0.14 0.185 0.14 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_R

VIA M2M3_PR_M
  LAYER met2 ;
    RECT -0.14 -0.185 0.14 0.185 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_M

VIA M2M3_PR_MR
  LAYER met2 ;
    RECT -0.185 -0.14 0.185 0.14 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_MR

VIA M2M3_PR_C
  LAYER met2 ;
    RECT -0.185 -0.185 0.185 0.185 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_C

VIA M3M4_PR
  LAYER met3 ;
    RECT -0.19 -0.16 0.19 0.16 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR

VIA M3M4_PR_R
  LAYER met3 ;
    RECT -0.16 -0.19 0.16 0.19 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_R

VIA M3M4_PR_M
  LAYER met3 ;
    RECT -0.19 -0.16 0.19 0.16 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_M

VIA M3M4_PR_MR
  LAYER met3 ;
    RECT -0.16 -0.19 0.16 0.19 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_MR

VIA M3M4_PR_C
  LAYER met3 ;
    RECT -0.19 -0.19 0.19 0.19 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_C

VIA M4M5_PR
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR

VIA M4M5_PR_R
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_R

VIA M4M5_PR_M
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_M

VIA M4M5_PR_MR
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_MR

VIA M4M5_PR_C
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_C

SITE unit
  CLASS CORE ;
  SYMMETRY Y ;
  SIZE 0.46 BY 2.72 ;
END unit

SITE unithddbl
  CLASS CORE ;
  SIZE 0.46 BY 5.44 ;
END unithddbl

MACRO sb_2__0_
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  SIZE 103.96 BY 125.12 ;
  SYMMETRY X Y ;
  PIN pReset[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 74.22 0.595 74.36 ;
    END
  END pReset[0]
  PIN chany_top_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.38 124.635 72.52 125.12 ;
    END
  END chany_top_in[0]
  PIN chany_top_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 61.03 124.32 61.33 125.12 ;
    END
  END chany_top_in[1]
  PIN chany_top_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.28 124.635 33.42 125.12 ;
    END
  END chany_top_in[2]
  PIN chany_top_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.2 124.635 57.34 125.12 ;
    END
  END chany_top_in[3]
  PIN chany_top_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.22 124.635 51.36 125.12 ;
    END
  END chany_top_in[4]
  PIN chany_top_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.34 124.635 61.48 125.12 ;
    END
  END chany_top_in[5]
  PIN chany_top_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.36 124.635 55.5 125.12 ;
    END
  END chany_top_in[6]
  PIN chany_top_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.62 124.635 69.76 125.12 ;
    END
  END chany_top_in[7]
  PIN chany_top_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.3 124.635 73.44 125.12 ;
    END
  END chany_top_in[8]
  PIN chany_top_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.7 124.635 68.84 125.12 ;
    END
  END chany_top_in[9]
  PIN chany_top_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.78 124.635 90.92 125.12 ;
    END
  END chany_top_in[10]
  PIN chany_top_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.36 124.635 78.5 125.12 ;
    END
  END chany_top_in[11]
  PIN chany_top_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.46 124.635 71.6 125.12 ;
    END
  END chany_top_in[12]
  PIN chany_top_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.78 124.635 67.92 125.12 ;
    END
  END chany_top_in[13]
  PIN chany_top_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.52 124.635 76.66 125.12 ;
    END
  END chany_top_in[14]
  PIN chany_top_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.46 124.635 94.6 125.12 ;
    END
  END chany_top_in[15]
  PIN chany_top_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.54 124.635 70.68 125.12 ;
    END
  END chany_top_in[16]
  PIN chany_top_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.86 124.635 90 125.12 ;
    END
  END chany_top_in[17]
  PIN chany_top_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.02 124.635 88.16 125.12 ;
    END
  END chany_top_in[18]
  PIN chany_top_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.54 124.635 93.68 125.12 ;
    END
  END chany_top_in[19]
  PIN chany_top_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.14 124.635 75.28 125.12 ;
    END
  END chany_top_in[20]
  PIN chany_top_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.28 124.635 56.42 125.12 ;
    END
  END chany_top_in[21]
  PIN chany_top_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.88 124.635 38.02 125.12 ;
    END
  END chany_top_in[22]
  PIN chany_top_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.86 124.635 44 125.12 ;
    END
  END chany_top_in[23]
  PIN chany_top_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.2 124.635 34.34 125.12 ;
    END
  END chany_top_in[24]
  PIN chany_top_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.94 124.635 43.08 125.12 ;
    END
  END chany_top_in[25]
  PIN chany_top_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.7 124.635 91.84 125.12 ;
    END
  END chany_top_in[26]
  PIN chany_top_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.12 124.635 81.26 125.12 ;
    END
  END chany_top_in[27]
  PIN chany_top_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.2 124.635 80.34 125.12 ;
    END
  END chany_top_in[28]
  PIN chany_top_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.28 124.635 79.42 125.12 ;
    END
  END chany_top_in[29]
  PIN top_left_grid_pin_44_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.18 119.195 17.32 119.68 ;
    END
  END top_left_grid_pin_44_[0]
  PIN top_left_grid_pin_45_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.12 119.195 12.26 119.68 ;
    END
  END top_left_grid_pin_45_[0]
  PIN top_left_grid_pin_46_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.02 119.195 19.16 119.68 ;
    END
  END top_left_grid_pin_46_[0]
  PIN top_left_grid_pin_47_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.4 119.195 20.54 119.68 ;
    END
  END top_left_grid_pin_47_[0]
  PIN top_left_grid_pin_48_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.84 119.195 3.98 119.68 ;
    END
  END top_left_grid_pin_48_[0]
  PIN top_left_grid_pin_49_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.42 119.195 14.56 119.68 ;
    END
  END top_left_grid_pin_49_[0]
  PIN top_left_grid_pin_50_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.2 119.195 11.34 119.68 ;
    END
  END top_left_grid_pin_50_[0]
  PIN top_left_grid_pin_51_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.1 119.195 18.24 119.68 ;
    END
  END top_left_grid_pin_51_[0]
  PIN top_right_grid_pin_1_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.18 124.635 63.32 125.12 ;
    END
  END top_right_grid_pin_1_[0]
  PIN chanx_left_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 69.8 0.595 69.94 ;
    END
  END chanx_left_in[0]
  PIN chanx_left_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 106.95 0.8 107.25 ;
    END
  END chanx_left_in[1]
  PIN chanx_left_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 115.02 0.595 115.16 ;
    END
  END chanx_left_in[2]
  PIN chanx_left_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 47.36 0.595 47.5 ;
    END
  END chanx_left_in[3]
  PIN chanx_left_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 72.52 0.595 72.66 ;
    END
  END chanx_left_in[4]
  PIN chanx_left_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 63.34 0.595 63.48 ;
    END
  END chanx_left_in[5]
  PIN chanx_left_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 48.04 0.595 48.18 ;
    END
  END chanx_left_in[6]
  PIN chanx_left_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 71.84 0.595 71.98 ;
    END
  END chanx_left_in[7]
  PIN chanx_left_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 45.32 0.595 45.46 ;
    END
  END chanx_left_in[8]
  PIN chanx_left_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 101.51 0.8 101.81 ;
    END
  END chanx_left_in[9]
  PIN chanx_left_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 50.08 0.595 50.22 ;
    END
  END chanx_left_in[10]
  PIN chanx_left_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 58.92 0.595 59.06 ;
    END
  END chanx_left_in[11]
  PIN chanx_left_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 85.1 0.595 85.24 ;
    END
  END chanx_left_in[12]
  PIN chanx_left_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 105.59 0.8 105.89 ;
    END
  END chanx_left_in[13]
  PIN chanx_left_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 95.39 0.8 95.69 ;
    END
  END chanx_left_in[14]
  PIN chanx_left_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 102.44 0.595 102.58 ;
    END
  END chanx_left_in[15]
  PIN chanx_left_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 104.48 0.595 104.62 ;
    END
  END chanx_left_in[16]
  PIN chanx_left_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 98.79 0.8 99.09 ;
    END
  END chanx_left_in[17]
  PIN chanx_left_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 111.03 0.8 111.33 ;
    END
  END chanx_left_in[18]
  PIN chanx_left_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 87.91 0.8 88.21 ;
    END
  END chanx_left_in[19]
  PIN chanx_left_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 88.5 0.595 88.64 ;
    END
  END chanx_left_in[20]
  PIN chanx_left_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 102.87 0.8 103.17 ;
    END
  END chanx_left_in[21]
  PIN chanx_left_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 81.11 0.8 81.41 ;
    END
  END chanx_left_in[22]
  PIN chanx_left_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 58.24 0.595 58.38 ;
    END
  END chanx_left_in[23]
  PIN chanx_left_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 56.2 0.595 56.34 ;
    END
  END chanx_left_in[24]
  PIN chanx_left_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 108.31 0.8 108.61 ;
    END
  END chanx_left_in[25]
  PIN chanx_left_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 86.55 0.8 86.85 ;
    END
  END chanx_left_in[26]
  PIN chanx_left_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 112.39 0.8 112.69 ;
    END
  END chanx_left_in[27]
  PIN chanx_left_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 100.15 0.8 100.45 ;
    END
  END chanx_left_in[28]
  PIN chanx_left_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 104.23 0.8 104.53 ;
    END
  END chanx_left_in[29]
  PIN left_bottom_grid_pin_1_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 66.06 0.595 66.2 ;
    END
  END left_bottom_grid_pin_1_[0]
  PIN left_bottom_grid_pin_3_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 94.03 0.8 94.33 ;
    END
  END left_bottom_grid_pin_3_[0]
  PIN left_bottom_grid_pin_5_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 113.75 0.8 114.05 ;
    END
  END left_bottom_grid_pin_5_[0]
  PIN left_bottom_grid_pin_7_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 97.43 0.8 97.73 ;
    END
  END left_bottom_grid_pin_7_[0]
  PIN left_bottom_grid_pin_9_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 64.02 0.595 64.16 ;
    END
  END left_bottom_grid_pin_9_[0]
  PIN left_bottom_grid_pin_11_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 92.67 0.8 92.97 ;
    END
  END left_bottom_grid_pin_11_[0]
  PIN left_bottom_grid_pin_13_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 68.78 0.595 68.92 ;
    END
  END left_bottom_grid_pin_13_[0]
  PIN left_bottom_grid_pin_15_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 89.27 0.8 89.57 ;
    END
  END left_bottom_grid_pin_15_[0]
  PIN left_bottom_grid_pin_17_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 67.08 0.595 67.22 ;
    END
  END left_bottom_grid_pin_17_[0]
  PIN ccff_head[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.72 124.635 39.86 125.12 ;
    END
  END ccff_head[0]
  PIN chany_top_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.96 124.635 83.1 125.12 ;
    END
  END chany_top_out[0]
  PIN chany_top_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.88 124.635 84.02 125.12 ;
    END
  END chany_top_out[1]
  PIN chany_top_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.72 124.635 85.86 125.12 ;
    END
  END chany_top_out[2]
  PIN chany_top_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.8 124.635 84.94 125.12 ;
    END
  END chany_top_out[3]
  PIN chany_top_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.62 124.635 46.76 125.12 ;
    END
  END chany_top_out[4]
  PIN chany_top_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 37.11 124.32 37.41 125.12 ;
    END
  END chany_top_out[5]
  PIN chany_top_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.02 124.635 65.16 125.12 ;
    END
  END chany_top_out[6]
  PIN chany_top_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.78 124.635 44.92 125.12 ;
    END
  END chany_top_out[7]
  PIN chany_top_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.04 124.635 59.18 125.12 ;
    END
  END chany_top_out[8]
  PIN chany_top_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.62 124.635 92.76 125.12 ;
    END
  END chany_top_out[9]
  PIN chany_top_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.64 124.635 40.78 125.12 ;
    END
  END chany_top_out[10]
  PIN chany_top_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.94 124.635 66.08 125.12 ;
    END
  END chany_top_out[11]
  PIN chany_top_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.38 124.635 95.52 125.12 ;
    END
  END chany_top_out[12]
  PIN chany_top_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.7 124.635 45.84 125.12 ;
    END
  END chany_top_out[13]
  PIN chany_top_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.1 124.635 64.24 125.12 ;
    END
  END chany_top_out[14]
  PIN chany_top_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.44 124.635 54.58 125.12 ;
    END
  END chany_top_out[15]
  PIN chany_top_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.96 124.635 37.1 125.12 ;
    END
  END chany_top_out[16]
  PIN chany_top_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.22 124.635 74.36 125.12 ;
    END
  END chany_top_out[17]
  PIN chany_top_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.04 124.635 82.18 125.12 ;
    END
  END chany_top_out[18]
  PIN chany_top_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.3 124.635 50.44 125.12 ;
    END
  END chany_top_out[19]
  PIN chany_top_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.06 124.635 53.2 125.12 ;
    END
  END chany_top_out[20]
  PIN chany_top_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.92 124.635 49.06 125.12 ;
    END
  END chany_top_out[21]
  PIN chany_top_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.26 124.635 62.4 125.12 ;
    END
  END chany_top_out[22]
  PIN chany_top_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.86 124.635 67 125.12 ;
    END
  END chany_top_out[23]
  PIN chany_top_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.64 124.635 86.78 125.12 ;
    END
  END chany_top_out[24]
  PIN chany_top_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48 124.635 48.14 125.12 ;
    END
  END chany_top_out[25]
  PIN chany_top_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.12 124.635 58.26 125.12 ;
    END
  END chany_top_out[26]
  PIN chany_top_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.14 124.635 52.28 125.12 ;
    END
  END chany_top_out[27]
  PIN chany_top_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.8 124.635 38.94 125.12 ;
    END
  END chany_top_out[28]
  PIN chany_top_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.44 124.635 77.58 125.12 ;
    END
  END chany_top_out[29]
  PIN chanx_left_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 85.19 0.8 85.49 ;
    END
  END chanx_left_out[0]
  PIN chanx_left_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 55.52 0.595 55.66 ;
    END
  END chanx_left_out[1]
  PIN chanx_left_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 60.96 0.595 61.1 ;
    END
  END chanx_left_out[2]
  PIN chanx_left_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 83.83 0.8 84.13 ;
    END
  END chanx_left_out[3]
  PIN chanx_left_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 115.7 0.595 115.84 ;
    END
  END chanx_left_out[4]
  PIN chanx_left_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 61.64 0.595 61.78 ;
    END
  END chanx_left_out[5]
  PIN chanx_left_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 87.82 0.595 87.96 ;
    END
  END chanx_left_out[6]
  PIN chanx_left_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 94.28 0.595 94.42 ;
    END
  END chanx_left_out[7]
  PIN chanx_left_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 82.72 0.595 82.86 ;
    END
  END chanx_left_out[8]
  PIN chanx_left_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 99.04 0.595 99.18 ;
    END
  END chanx_left_out[9]
  PIN chanx_left_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 117.74 0.595 117.88 ;
    END
  END chanx_left_out[10]
  PIN chanx_left_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 93.6 0.595 93.74 ;
    END
  END chanx_left_out[11]
  PIN chanx_left_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 99.72 0.595 99.86 ;
    END
  END chanx_left_out[12]
  PIN chanx_left_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 91.22 0.595 91.36 ;
    END
  END chanx_left_out[13]
  PIN chanx_left_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 80.68 0.595 80.82 ;
    END
  END chanx_left_out[14]
  PIN chanx_left_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 112.98 0.595 113.12 ;
    END
  END chanx_left_out[15]
  PIN chanx_left_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 101.76 0.595 101.9 ;
    END
  END chanx_left_out[16]
  PIN chanx_left_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 90.54 0.595 90.68 ;
    END
  END chanx_left_out[17]
  PIN chanx_left_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 110.26 0.595 110.4 ;
    END
  END chanx_left_out[18]
  PIN chanx_left_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 109.67 0.8 109.97 ;
    END
  END chanx_left_out[19]
  PIN chanx_left_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 82.47 0.8 82.77 ;
    END
  END chanx_left_out[20]
  PIN chanx_left_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 97 0.595 97.14 ;
    END
  END chanx_left_out[21]
  PIN chanx_left_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 79.75 0.8 80.05 ;
    END
  END chanx_left_out[22]
  PIN chanx_left_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 83.4 0.595 83.54 ;
    END
  END chanx_left_out[23]
  PIN chanx_left_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 107.54 0.595 107.68 ;
    END
  END chanx_left_out[24]
  PIN chanx_left_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 109.58 0.595 109.72 ;
    END
  END chanx_left_out[25]
  PIN chanx_left_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 80 0.595 80.14 ;
    END
  END chanx_left_out[26]
  PIN chanx_left_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 112.3 0.595 112.44 ;
    END
  END chanx_left_out[27]
  PIN chanx_left_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 105.16 0.595 105.3 ;
    END
  END chanx_left_out[28]
  PIN chanx_left_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 106.86 0.595 107 ;
    END
  END chanx_left_out[29]
  PIN ccff_tail[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 85.78 0.595 85.92 ;
    END
  END ccff_tail[0]
  PIN pReset_W_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 95.98 0.595 96.12 ;
    END
  END pReset_W_in
  PIN pReset_N_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.58 124.635 35.72 125.12 ;
    END
  END pReset_N_out
  PIN prog_clk_0_N_in
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER met2 ;
        RECT 42.02 124.635 42.16 125.12 ;
    END
  END prog_clk_0_N_in
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0 17.44 3.2 20.64 ;
        RECT 100.76 17.44 103.96 20.64 ;
        RECT 0 58.24 3.2 61.44 ;
        RECT 100.76 58.24 103.96 61.44 ;
        RECT 0 99.04 3.2 102.24 ;
        RECT 100.76 99.04 103.96 102.24 ;
      LAYER met4 ;
        RECT 13.5 0 14.1 0.6 ;
        RECT 44.78 0 45.38 0.6 ;
        RECT 74.22 0 74.82 0.6 ;
        RECT 13.5 119.08 14.1 119.68 ;
        RECT 44.78 124.52 45.38 125.12 ;
        RECT 74.22 124.52 74.82 125.12 ;
      LAYER met1 ;
        RECT 0 2.48 0.48 2.96 ;
        RECT 103.48 2.48 103.96 2.96 ;
        RECT 0 7.92 0.48 8.4 ;
        RECT 103.48 7.92 103.96 8.4 ;
        RECT 0 13.36 0.48 13.84 ;
        RECT 103.48 13.36 103.96 13.84 ;
        RECT 0 18.8 0.48 19.28 ;
        RECT 103.48 18.8 103.96 19.28 ;
        RECT 0 24.24 0.48 24.72 ;
        RECT 103.48 24.24 103.96 24.72 ;
        RECT 0 29.68 0.48 30.16 ;
        RECT 103.48 29.68 103.96 30.16 ;
        RECT 0 35.12 0.48 35.6 ;
        RECT 103.48 35.12 103.96 35.6 ;
        RECT 0 40.56 0.48 41.04 ;
        RECT 103.48 40.56 103.96 41.04 ;
        RECT 0 46 0.48 46.48 ;
        RECT 103.48 46 103.96 46.48 ;
        RECT 0 51.44 0.48 51.92 ;
        RECT 103.48 51.44 103.96 51.92 ;
        RECT 0 56.88 0.48 57.36 ;
        RECT 103.48 56.88 103.96 57.36 ;
        RECT 0 62.32 0.48 62.8 ;
        RECT 103.48 62.32 103.96 62.8 ;
        RECT 0 67.76 0.48 68.24 ;
        RECT 103.48 67.76 103.96 68.24 ;
        RECT 0 73.2 0.48 73.68 ;
        RECT 103.48 73.2 103.96 73.68 ;
        RECT 0 78.64 0.48 79.12 ;
        RECT 103.48 78.64 103.96 79.12 ;
        RECT 0 84.08 0.48 84.56 ;
        RECT 103.48 84.08 103.96 84.56 ;
        RECT 0 89.52 0.48 90 ;
        RECT 103.48 89.52 103.96 90 ;
        RECT 0 94.96 0.48 95.44 ;
        RECT 103.48 94.96 103.96 95.44 ;
        RECT 0 100.4 0.48 100.88 ;
        RECT 103.48 100.4 103.96 100.88 ;
        RECT 0 105.84 0.48 106.32 ;
        RECT 103.48 105.84 103.96 106.32 ;
        RECT 0 111.28 0.48 111.76 ;
        RECT 103.48 111.28 103.96 111.76 ;
        RECT 0 116.72 0.48 117.2 ;
        RECT 103.48 116.72 103.96 117.2 ;
        RECT 30.36 122.16 30.84 122.64 ;
        RECT 103.48 122.16 103.96 122.64 ;
    END
  END VDD
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0 37.84 3.2 41.04 ;
        RECT 100.76 37.84 103.96 41.04 ;
        RECT 0 78.64 3.2 81.84 ;
        RECT 100.76 78.64 103.96 81.84 ;
      LAYER met4 ;
        RECT 59.5 0 60.1 0.6 ;
        RECT 88.94 0 89.54 0.6 ;
        RECT 59.5 124.52 60.1 125.12 ;
        RECT 88.94 124.52 89.54 125.12 ;
      LAYER met1 ;
        RECT 0 -0.24 0.48 0.24 ;
        RECT 103.48 -0.24 103.96 0.24 ;
        RECT 0 5.2 0.48 5.68 ;
        RECT 103.48 5.2 103.96 5.68 ;
        RECT 0 10.64 0.48 11.12 ;
        RECT 103.48 10.64 103.96 11.12 ;
        RECT 0 16.08 0.48 16.56 ;
        RECT 103.48 16.08 103.96 16.56 ;
        RECT 0 21.52 0.48 22 ;
        RECT 103.48 21.52 103.96 22 ;
        RECT 0 26.96 0.48 27.44 ;
        RECT 103.48 26.96 103.96 27.44 ;
        RECT 0 32.4 0.48 32.88 ;
        RECT 103.48 32.4 103.96 32.88 ;
        RECT 0 37.84 0.48 38.32 ;
        RECT 103.48 37.84 103.96 38.32 ;
        RECT 0 43.28 0.48 43.76 ;
        RECT 103.48 43.28 103.96 43.76 ;
        RECT 0 48.72 0.48 49.2 ;
        RECT 103.48 48.72 103.96 49.2 ;
        RECT 0 54.16 0.48 54.64 ;
        RECT 103.48 54.16 103.96 54.64 ;
        RECT 0 59.6 0.48 60.08 ;
        RECT 103.48 59.6 103.96 60.08 ;
        RECT 0 65.04 0.48 65.52 ;
        RECT 103.48 65.04 103.96 65.52 ;
        RECT 0 70.48 0.48 70.96 ;
        RECT 103.48 70.48 103.96 70.96 ;
        RECT 0 75.92 0.48 76.4 ;
        RECT 103.48 75.92 103.96 76.4 ;
        RECT 0 81.36 0.48 81.84 ;
        RECT 103.48 81.36 103.96 81.84 ;
        RECT 0 86.8 0.48 87.28 ;
        RECT 103.48 86.8 103.96 87.28 ;
        RECT 0 92.24 0.48 92.72 ;
        RECT 103.48 92.24 103.96 92.72 ;
        RECT 0 97.68 0.48 98.16 ;
        RECT 103.48 97.68 103.96 98.16 ;
        RECT 0 103.12 0.48 103.6 ;
        RECT 103.48 103.12 103.96 103.6 ;
        RECT 0 108.56 0.48 109.04 ;
        RECT 103.48 108.56 103.96 109.04 ;
        RECT 0 114 0.48 114.48 ;
        RECT 103.48 114 103.96 114.48 ;
        RECT 0 119.44 0.48 119.92 ;
        RECT 103.48 119.44 103.96 119.92 ;
        RECT 30.36 124.88 30.84 125.36 ;
        RECT 103.48 124.88 103.96 125.36 ;
    END
  END VSS
  OBS
    LAYER met1 ;
      POLYGON 103.2 125.36 103.2 124.88 89.4 124.88 89.4 124.87 89.08 124.87 89.08 124.88 59.96 124.88 59.96 124.87 59.64 124.87 59.64 124.88 31.12 124.88 31.12 125.36 ;
      RECT 0.76 119.44 52.76 119.92 ;
      POLYGON 89.4 0.25 89.4 0.24 103.2 0.24 103.2 -0.24 0.76 -0.24 0.76 0.24 59.64 0.24 59.64 0.25 59.96 0.25 59.96 0.24 89.08 0.24 89.08 0.25 ;
      POLYGON 103.2 124.84 103.2 124.6 103.68 124.6 103.68 122.92 103.2 122.92 103.2 121.88 103.68 121.88 103.68 120.2 103.2 120.2 103.2 119.16 103.68 119.16 103.68 117.48 103.2 117.48 103.2 116.44 103.68 116.44 103.68 114.76 103.2 114.76 103.2 113.72 103.68 113.72 103.68 112.04 103.2 112.04 103.2 111 103.68 111 103.68 109.32 103.2 109.32 103.2 108.28 103.68 108.28 103.68 106.6 103.2 106.6 103.2 105.56 103.68 105.56 103.68 103.88 103.2 103.88 103.2 102.84 103.68 102.84 103.68 101.16 103.2 101.16 103.2 100.12 103.68 100.12 103.68 98.44 103.2 98.44 103.2 97.4 103.68 97.4 103.68 95.72 103.2 95.72 103.2 94.68 103.68 94.68 103.68 93 103.2 93 103.2 91.96 103.68 91.96 103.68 90.28 103.2 90.28 103.2 89.24 103.68 89.24 103.68 87.56 103.2 87.56 103.2 86.52 103.68 86.52 103.68 84.84 103.2 84.84 103.2 83.8 103.68 83.8 103.68 82.12 103.2 82.12 103.2 81.08 103.68 81.08 103.68 79.4 103.2 79.4 103.2 78.36 103.68 78.36 103.68 76.68 103.2 76.68 103.2 75.64 103.68 75.64 103.68 73.96 103.2 73.96 103.2 72.92 103.68 72.92 103.68 71.24 103.2 71.24 103.2 70.2 103.68 70.2 103.68 68.52 103.2 68.52 103.2 67.48 103.68 67.48 103.68 65.8 103.2 65.8 103.2 64.76 103.68 64.76 103.68 63.08 103.2 63.08 103.2 62.04 103.68 62.04 103.68 60.36 103.2 60.36 103.2 59.32 103.68 59.32 103.68 57.64 103.2 57.64 103.2 56.6 103.68 56.6 103.68 54.92 103.2 54.92 103.2 53.88 103.68 53.88 103.68 52.2 103.2 52.2 103.2 51.16 103.68 51.16 103.68 49.48 103.2 49.48 103.2 48.44 103.68 48.44 103.68 46.76 103.2 46.76 103.2 45.72 103.68 45.72 103.68 44.04 103.2 44.04 103.2 43 103.68 43 103.68 41.32 103.2 41.32 103.2 40.28 103.68 40.28 103.68 38.6 103.2 38.6 103.2 37.56 103.68 37.56 103.68 35.88 103.2 35.88 103.2 34.84 103.68 34.84 103.68 33.16 103.2 33.16 103.2 32.12 103.68 32.12 103.68 30.44 103.2 30.44 103.2 29.4 103.68 29.4 103.68 27.72 103.2 27.72 103.2 26.68 103.68 26.68 103.68 25 103.2 25 103.2 23.96 103.68 23.96 103.68 22.28 103.2 22.28 103.2 21.24 103.68 21.24 103.68 19.56 103.2 19.56 103.2 18.52 103.68 18.52 103.68 16.84 103.2 16.84 103.2 15.8 103.68 15.8 103.68 14.12 103.2 14.12 103.2 13.08 103.68 13.08 103.68 11.4 103.2 11.4 103.2 10.36 103.68 10.36 103.68 8.68 103.2 8.68 103.2 7.64 103.68 7.64 103.68 5.96 103.2 5.96 103.2 4.92 103.68 4.92 103.68 3.24 103.2 3.24 103.2 2.2 103.68 2.2 103.68 0.52 103.2 0.52 103.2 0.28 0.76 0.28 0.76 0.52 0.28 0.52 0.28 2.2 0.76 2.2 0.76 3.24 0.28 3.24 0.28 4.92 0.76 4.92 0.76 5.96 0.28 5.96 0.28 7.64 0.76 7.64 0.76 8.68 0.28 8.68 0.28 10.36 0.76 10.36 0.76 11.4 0.28 11.4 0.28 13.08 0.76 13.08 0.76 14.12 0.28 14.12 0.28 15.8 0.76 15.8 0.76 16.84 0.28 16.84 0.28 18.52 0.76 18.52 0.76 19.56 0.28 19.56 0.28 21.24 0.76 21.24 0.76 22.28 0.28 22.28 0.28 23.96 0.76 23.96 0.76 25 0.28 25 0.28 26.68 0.76 26.68 0.76 27.72 0.28 27.72 0.28 29.4 0.76 29.4 0.76 30.44 0.28 30.44 0.28 32.12 0.76 32.12 0.76 33.16 0.28 33.16 0.28 34.84 0.76 34.84 0.76 35.88 0.28 35.88 0.28 37.56 0.76 37.56 0.76 38.6 0.28 38.6 0.28 40.28 0.76 40.28 0.76 41.32 0.28 41.32 0.28 43 0.76 43 0.76 44.04 0.28 44.04 0.28 45.04 0.875 45.04 0.875 45.74 0.76 45.74 0.76 46.76 0.28 46.76 0.28 47.08 0.875 47.08 0.875 48.46 0.76 48.46 0.76 49.48 0.28 49.48 0.28 49.8 0.875 49.8 0.875 50.5 0.28 50.5 0.28 51.16 0.76 51.16 0.76 52.2 0.28 52.2 0.28 53.88 0.76 53.88 0.76 54.92 0.28 54.92 0.28 55.24 0.875 55.24 0.875 56.62 0.76 56.62 0.76 57.64 0.28 57.64 0.28 57.96 0.875 57.96 0.875 59.34 0.76 59.34 0.76 60.36 0.28 60.36 0.28 60.68 0.875 60.68 0.875 62.06 0.76 62.06 0.76 63.06 0.875 63.06 0.875 64.44 0.28 64.44 0.28 64.76 0.76 64.76 0.76 65.78 0.875 65.78 0.875 66.48 0.28 66.48 0.28 66.8 0.875 66.8 0.875 67.5 0.76 67.5 0.76 68.5 0.875 68.5 0.875 69.2 0.28 69.2 0.28 69.52 0.875 69.52 0.875 70.22 0.76 70.22 0.76 71.24 0.28 71.24 0.28 71.56 0.875 71.56 0.875 72.94 0.76 72.94 0.76 73.94 0.875 73.94 0.875 74.64 0.28 74.64 0.28 75.64 0.76 75.64 0.76 76.68 0.28 76.68 0.28 78.36 0.76 78.36 0.76 79.4 0.28 79.4 0.28 79.72 0.875 79.72 0.875 81.1 0.76 81.1 0.76 82.12 0.28 82.12 0.28 82.44 0.875 82.44 0.875 83.82 0.76 83.82 0.76 84.82 0.875 84.82 0.875 86.2 0.28 86.2 0.28 86.52 0.76 86.52 0.76 87.54 0.875 87.54 0.875 88.92 0.28 88.92 0.28 89.24 0.76 89.24 0.76 90.26 0.875 90.26 0.875 91.64 0.28 91.64 0.28 91.96 0.76 91.96 0.76 93 0.28 93 0.28 93.32 0.875 93.32 0.875 94.7 0.76 94.7 0.76 95.7 0.875 95.7 0.875 96.4 0.28 96.4 0.28 96.72 0.875 96.72 0.875 97.42 0.76 97.42 0.76 98.44 0.28 98.44 0.28 98.76 0.875 98.76 0.875 100.14 0.76 100.14 0.76 101.16 0.28 101.16 0.28 101.48 0.875 101.48 0.875 102.86 0.76 102.86 0.76 103.88 0.28 103.88 0.28 104.2 0.875 104.2 0.875 105.58 0.76 105.58 0.76 106.58 0.875 106.58 0.875 107.96 0.28 107.96 0.28 108.28 0.76 108.28 0.76 109.3 0.875 109.3 0.875 110.68 0.28 110.68 0.28 111 0.76 111 0.76 112.02 0.875 112.02 0.875 113.4 0.28 113.4 0.28 113.72 0.76 113.72 0.76 114.74 0.875 114.74 0.875 116.12 0.28 116.12 0.28 116.44 0.76 116.44 0.76 117.46 0.875 117.46 0.875 118.16 0.28 118.16 0.28 119.16 0.76 119.16 0.76 119.4 30.64 119.4 30.64 121.88 31.12 121.88 31.12 122.92 30.64 122.92 30.64 124.6 31.12 124.6 31.12 124.84 ;
    LAYER met2 ;
      RECT 89.1 124.815 89.38 125.185 ;
      RECT 59.66 124.815 59.94 125.185 ;
      POLYGON 55.08 125.02 55.08 124.88 55.04 124.88 55.04 95.98 54.9 95.98 54.9 125.02 ;
      POLYGON 53.66 125.02 53.66 120.12 53.52 120.12 53.52 124.88 53.48 124.88 53.48 125.02 ;
      POLYGON 48.6 125.02 48.6 112.64 48.46 112.64 48.46 124.88 48.42 124.88 48.42 125.02 ;
      POLYGON 44.5 125.02 44.5 124.88 44.46 124.88 44.46 118.76 44.32 118.76 44.32 125.02 ;
      POLYGON 33.88 125.02 33.88 102.1 33.74 102.1 33.74 124.88 33.7 124.88 33.7 125.02 ;
      RECT 75.54 124.11 75.8 124.43 ;
      RECT 18.5 118.67 18.76 118.99 ;
      RECT 89.1 -0.065 89.38 0.305 ;
      RECT 59.66 -0.065 59.94 0.305 ;
      POLYGON 103.68 124.84 103.68 0.28 0.28 0.28 0.28 119.4 3.56 119.4 3.56 118.915 4.26 118.915 4.26 119.4 10.92 119.4 10.92 118.915 11.62 118.915 11.62 119.4 11.84 119.4 11.84 118.915 12.54 118.915 12.54 119.4 14.14 119.4 14.14 118.915 14.84 118.915 14.84 119.4 16.9 119.4 16.9 118.915 17.6 118.915 17.6 119.4 17.82 119.4 17.82 118.915 18.52 118.915 18.52 119.4 18.74 119.4 18.74 118.915 19.44 118.915 19.44 119.4 20.12 119.4 20.12 118.915 20.82 118.915 20.82 119.4 30.64 119.4 30.64 124.84 33 124.84 33 124.355 33.7 124.355 33.7 124.84 33.92 124.84 33.92 124.355 34.62 124.355 34.62 124.84 35.3 124.84 35.3 124.355 36 124.355 36 124.84 36.68 124.84 36.68 124.355 37.38 124.355 37.38 124.84 37.6 124.84 37.6 124.355 38.3 124.355 38.3 124.84 38.52 124.84 38.52 124.355 39.22 124.355 39.22 124.84 39.44 124.84 39.44 124.355 40.14 124.355 40.14 124.84 40.36 124.84 40.36 124.355 41.06 124.355 41.06 124.84 41.74 124.84 41.74 124.355 42.44 124.355 42.44 124.84 42.66 124.84 42.66 124.355 43.36 124.355 43.36 124.84 43.58 124.84 43.58 124.355 44.28 124.355 44.28 124.84 44.5 124.84 44.5 124.355 45.2 124.355 45.2 124.84 45.42 124.84 45.42 124.355 46.12 124.355 46.12 124.84 46.34 124.84 46.34 124.355 47.04 124.355 47.04 124.84 47.72 124.84 47.72 124.355 48.42 124.355 48.42 124.84 48.64 124.84 48.64 124.355 49.34 124.355 49.34 124.84 50.02 124.84 50.02 124.355 50.72 124.355 50.72 124.84 50.94 124.84 50.94 124.355 51.64 124.355 51.64 124.84 51.86 124.84 51.86 124.355 52.56 124.355 52.56 124.84 52.78 124.84 52.78 124.355 53.48 124.355 53.48 124.84 54.16 124.84 54.16 124.355 54.86 124.355 54.86 124.84 55.08 124.84 55.08 124.355 55.78 124.355 55.78 124.84 56 124.84 56 124.355 56.7 124.355 56.7 124.84 56.92 124.84 56.92 124.355 57.62 124.355 57.62 124.84 57.84 124.84 57.84 124.355 58.54 124.355 58.54 124.84 58.76 124.84 58.76 124.355 59.46 124.355 59.46 124.84 61.06 124.84 61.06 124.355 61.76 124.355 61.76 124.84 61.98 124.84 61.98 124.355 62.68 124.355 62.68 124.84 62.9 124.84 62.9 124.355 63.6 124.355 63.6 124.84 63.82 124.84 63.82 124.355 64.52 124.355 64.52 124.84 64.74 124.84 64.74 124.355 65.44 124.355 65.44 124.84 65.66 124.84 65.66 124.355 66.36 124.355 66.36 124.84 66.58 124.84 66.58 124.355 67.28 124.355 67.28 124.84 67.5 124.84 67.5 124.355 68.2 124.355 68.2 124.84 68.42 124.84 68.42 124.355 69.12 124.355 69.12 124.84 69.34 124.84 69.34 124.355 70.04 124.355 70.04 124.84 70.26 124.84 70.26 124.355 70.96 124.355 70.96 124.84 71.18 124.84 71.18 124.355 71.88 124.355 71.88 124.84 72.1 124.84 72.1 124.355 72.8 124.355 72.8 124.84 73.02 124.84 73.02 124.355 73.72 124.355 73.72 124.84 73.94 124.84 73.94 124.355 74.64 124.355 74.64 124.84 74.86 124.84 74.86 124.355 75.56 124.355 75.56 124.84 76.24 124.84 76.24 124.355 76.94 124.355 76.94 124.84 77.16 124.84 77.16 124.355 77.86 124.355 77.86 124.84 78.08 124.84 78.08 124.355 78.78 124.355 78.78 124.84 79 124.84 79 124.355 79.7 124.355 79.7 124.84 79.92 124.84 79.92 124.355 80.62 124.355 80.62 124.84 80.84 124.84 80.84 124.355 81.54 124.355 81.54 124.84 81.76 124.84 81.76 124.355 82.46 124.355 82.46 124.84 82.68 124.84 82.68 124.355 83.38 124.355 83.38 124.84 83.6 124.84 83.6 124.355 84.3 124.355 84.3 124.84 84.52 124.84 84.52 124.355 85.22 124.355 85.22 124.84 85.44 124.84 85.44 124.355 86.14 124.355 86.14 124.84 86.36 124.84 86.36 124.355 87.06 124.355 87.06 124.84 87.74 124.84 87.74 124.355 88.44 124.355 88.44 124.84 89.58 124.84 89.58 124.355 90.28 124.355 90.28 124.84 90.5 124.84 90.5 124.355 91.2 124.355 91.2 124.84 91.42 124.84 91.42 124.355 92.12 124.355 92.12 124.84 92.34 124.84 92.34 124.355 93.04 124.355 93.04 124.84 93.26 124.84 93.26 124.355 93.96 124.355 93.96 124.84 94.18 124.84 94.18 124.355 94.88 124.355 94.88 124.84 95.1 124.84 95.1 124.355 95.8 124.355 95.8 124.84 ;
    LAYER met4 ;
      POLYGON 57.665 124.945 57.665 124.615 57.65 124.615 57.65 69.55 57.35 69.55 57.35 124.615 57.335 124.615 57.335 124.945 ;
      POLYGON 49.385 124.945 49.385 124.615 49.37 124.615 49.37 59.35 49.07 59.35 49.07 124.615 49.055 124.615 49.055 124.945 ;
      POLYGON 32.825 124.945 32.825 124.615 32.81 124.615 32.81 106.95 32.51 106.95 32.51 124.615 32.495 124.615 32.495 124.945 ;
      POLYGON 103.56 124.72 103.56 0.4 89.94 0.4 89.94 1 88.54 1 88.54 0.4 75.22 0.4 75.22 1 73.82 1 73.82 0.4 60.5 0.4 60.5 1 59.1 1 59.1 0.4 45.78 0.4 45.78 1 44.38 1 44.38 0.4 14.5 0.4 14.5 1 13.1 1 13.1 0.4 0.4 0.4 0.4 119.28 13.1 119.28 13.1 118.68 14.5 118.68 14.5 119.28 30.76 119.28 30.76 124.72 36.71 124.72 36.71 123.92 37.81 123.92 37.81 124.72 44.38 124.72 44.38 124.12 45.78 124.12 45.78 124.72 59.1 124.72 59.1 124.12 60.5 124.12 60.5 124.72 60.63 124.72 60.63 123.92 61.73 123.92 61.73 124.72 73.82 124.72 73.82 124.12 75.22 124.12 75.22 124.72 88.54 124.72 88.54 124.12 89.94 124.12 89.94 124.72 ;
    LAYER met3 ;
      POLYGON 89.405 125.165 89.405 125.16 89.62 125.16 89.62 124.84 89.405 124.84 89.405 124.835 89.075 124.835 89.075 124.84 88.86 124.84 88.86 125.16 89.075 125.16 89.075 125.165 ;
      POLYGON 59.965 125.165 59.965 125.16 60.18 125.16 60.18 124.84 59.965 124.84 59.965 124.835 59.635 124.835 59.635 124.84 59.42 124.84 59.42 125.16 59.635 125.16 59.635 125.165 ;
      POLYGON 58.355 124.945 58.355 124.615 58.025 124.615 58.025 124.63 57.69 124.63 57.69 124.62 57.31 124.62 57.31 124.94 57.69 124.94 57.69 124.93 58.025 124.93 58.025 124.945 ;
      POLYGON 43.175 124.945 43.175 124.93 49.03 124.93 49.03 124.94 49.41 124.94 49.41 124.62 49.03 124.62 49.03 124.63 43.175 124.63 43.175 124.615 42.845 124.615 42.845 124.945 ;
      POLYGON 37.195 124.945 37.195 124.615 36.865 124.615 36.865 124.63 32.85 124.63 32.85 124.62 32.47 124.62 32.47 124.94 32.85 124.94 32.85 124.93 36.865 124.93 36.865 124.945 ;
      POLYGON 89.405 0.285 89.405 0.28 89.62 0.28 89.62 -0.04 89.405 -0.04 89.405 -0.045 89.075 -0.045 89.075 -0.04 88.86 -0.04 88.86 0.28 89.075 0.28 89.075 0.285 ;
      POLYGON 59.965 0.285 59.965 0.28 60.18 0.28 60.18 -0.04 59.965 -0.04 59.965 -0.045 59.635 -0.045 59.635 -0.04 59.42 -0.04 59.42 0.28 59.635 0.28 59.635 0.285 ;
      POLYGON 103.56 124.72 103.56 0.4 0.4 0.4 0.4 79.35 1.2 79.35 1.2 80.45 0.4 80.45 0.4 80.71 1.2 80.71 1.2 81.81 0.4 81.81 0.4 82.07 1.2 82.07 1.2 83.17 0.4 83.17 0.4 83.43 1.2 83.43 1.2 84.53 0.4 84.53 0.4 84.79 1.2 84.79 1.2 85.89 0.4 85.89 0.4 86.15 1.2 86.15 1.2 87.25 0.4 87.25 0.4 87.51 1.2 87.51 1.2 88.61 0.4 88.61 0.4 88.87 1.2 88.87 1.2 89.97 0.4 89.97 0.4 92.27 1.2 92.27 1.2 93.37 0.4 93.37 0.4 93.63 1.2 93.63 1.2 94.73 0.4 94.73 0.4 94.99 1.2 94.99 1.2 96.09 0.4 96.09 0.4 97.03 1.2 97.03 1.2 98.13 0.4 98.13 0.4 98.39 1.2 98.39 1.2 99.49 0.4 99.49 0.4 99.75 1.2 99.75 1.2 100.85 0.4 100.85 0.4 101.11 1.2 101.11 1.2 102.21 0.4 102.21 0.4 102.47 1.2 102.47 1.2 103.57 0.4 103.57 0.4 103.83 1.2 103.83 1.2 104.93 0.4 104.93 0.4 105.19 1.2 105.19 1.2 106.29 0.4 106.29 0.4 106.55 1.2 106.55 1.2 107.65 0.4 107.65 0.4 107.91 1.2 107.91 1.2 109.01 0.4 109.01 0.4 109.27 1.2 109.27 1.2 110.37 0.4 110.37 0.4 110.63 1.2 110.63 1.2 111.73 0.4 111.73 0.4 111.99 1.2 111.99 1.2 113.09 0.4 113.09 0.4 113.35 1.2 113.35 1.2 114.45 0.4 114.45 0.4 119.28 30.76 119.28 30.76 124.72 ;
    LAYER met5 ;
      POLYGON 102.36 123.52 102.36 103.84 99.16 103.84 99.16 97.44 102.36 97.44 102.36 83.44 99.16 83.44 99.16 77.04 102.36 77.04 102.36 63.04 99.16 63.04 99.16 56.64 102.36 56.64 102.36 42.64 99.16 42.64 99.16 36.24 102.36 36.24 102.36 22.24 99.16 22.24 99.16 15.84 102.36 15.84 102.36 1.6 1.6 1.6 1.6 15.84 4.8 15.84 4.8 22.24 1.6 22.24 1.6 36.24 4.8 36.24 4.8 42.64 1.6 42.64 1.6 56.64 4.8 56.64 4.8 63.04 1.6 63.04 1.6 77.04 4.8 77.04 4.8 83.44 1.6 83.44 1.6 97.44 4.8 97.44 4.8 103.84 1.6 103.84 1.6 118.08 31.96 118.08 31.96 123.52 ;
    LAYER li1 ;
      POLYGON 103.96 125.205 103.96 125.035 99.265 125.035 99.265 124.235 98.935 124.235 98.935 125.035 98.425 125.035 98.425 124.555 98.095 124.555 98.095 125.035 97.585 125.035 97.585 124.555 97.255 124.555 97.255 125.035 96.665 125.035 96.665 124.555 96.495 124.555 96.495 125.035 95.825 125.035 95.825 124.555 95.655 124.555 95.655 125.035 92.825 125.035 92.825 124.235 92.495 124.235 92.495 125.035 91.985 125.035 91.985 124.555 91.655 124.555 91.655 125.035 91.145 125.035 91.145 124.555 90.815 124.555 90.815 125.035 90.225 125.035 90.225 124.555 90.055 124.555 90.055 125.035 89.385 125.035 89.385 124.555 89.215 124.555 89.215 125.035 87.605 125.035 87.605 124.575 87.35 124.575 87.35 125.035 86.68 125.035 86.68 124.575 86.51 124.575 86.51 125.035 85.84 125.035 85.84 124.575 85.67 124.575 85.67 125.035 85 125.035 85 124.575 84.83 124.575 84.83 125.035 84.16 125.035 84.16 124.575 83.855 124.575 83.855 125.035 82.085 125.035 82.085 124.575 81.83 124.575 81.83 125.035 81.16 125.035 81.16 124.575 80.99 124.575 80.99 125.035 80.32 125.035 80.32 124.575 80.15 124.575 80.15 125.035 79.48 125.035 79.48 124.575 79.31 124.575 79.31 125.035 78.64 125.035 78.64 124.575 78.335 124.575 78.335 125.035 77.025 125.035 77.025 124.575 76.77 124.575 76.77 125.035 76.1 125.035 76.1 124.575 75.93 124.575 75.93 125.035 75.26 125.035 75.26 124.575 75.09 124.575 75.09 125.035 74.42 125.035 74.42 124.575 74.25 124.575 74.25 125.035 73.58 125.035 73.58 124.575 73.275 124.575 73.275 125.035 69.205 125.035 69.205 124.575 68.95 124.575 68.95 125.035 68.28 125.035 68.28 124.575 68.11 124.575 68.11 125.035 67.44 125.035 67.44 124.575 67.27 124.575 67.27 125.035 66.6 125.035 66.6 124.575 66.43 124.575 66.43 125.035 65.76 125.035 65.76 124.575 65.455 124.575 65.455 125.035 62.925 125.035 62.925 124.235 62.595 124.235 62.595 125.035 62.085 125.035 62.085 124.555 61.755 124.555 61.755 125.035 61.245 125.035 61.245 124.555 60.915 124.555 60.915 125.035 60.325 125.035 60.325 124.555 60.155 124.555 60.155 125.035 59.485 125.035 59.485 124.555 59.315 124.555 59.315 125.035 56.525 125.035 56.525 124.575 56.22 124.575 56.22 125.035 54.735 125.035 54.735 124.595 54.545 124.595 54.545 125.035 52.645 125.035 52.645 124.575 52.315 124.575 52.315 125.035 49.715 125.035 49.715 124.675 49.385 124.675 49.385 125.035 48.685 125.035 48.685 124.655 48.355 124.655 48.355 125.035 44.485 125.035 44.485 124.575 44.18 124.575 44.18 125.035 43.51 125.035 43.51 124.575 43.34 124.575 43.34 125.035 42.67 125.035 42.67 124.575 42.5 124.575 42.5 125.035 41.83 125.035 41.83 124.575 41.66 124.575 41.66 125.035 40.99 125.035 40.99 124.575 40.735 124.575 40.735 125.035 38.085 125.035 38.085 124.235 37.755 124.235 37.755 125.035 37.245 125.035 37.245 124.555 36.915 124.555 36.915 125.035 36.405 125.035 36.405 124.555 36.075 124.555 36.075 125.035 35.485 125.035 35.485 124.555 35.315 124.555 35.315 125.035 34.645 125.035 34.645 124.555 34.475 124.555 34.475 125.035 30.36 125.035 30.36 125.205 ;
      RECT 103.04 122.315 103.96 122.485 ;
      RECT 30.36 122.315 34.04 122.485 ;
      RECT 103.5 119.595 103.96 119.765 ;
      POLYGON 34.04 119.765 34.04 119.595 26.085 119.595 26.085 119.135 25.78 119.135 25.78 119.595 25.11 119.595 25.11 119.135 24.94 119.135 24.94 119.595 24.27 119.595 24.27 119.135 24.1 119.135 24.1 119.595 23.43 119.595 23.43 119.135 23.26 119.135 23.26 119.595 22.59 119.595 22.59 119.135 22.335 119.135 22.335 119.595 20.645 119.595 20.645 119.195 20.315 119.195 20.315 119.595 18.355 119.595 18.355 119.06 17.845 119.06 17.845 119.595 13.205 119.595 13.205 119.135 12.9 119.135 12.9 119.595 12.23 119.595 12.23 119.135 12.06 119.135 12.06 119.595 11.39 119.595 11.39 119.135 11.22 119.135 11.22 119.595 10.55 119.595 10.55 119.135 10.38 119.135 10.38 119.595 9.71 119.595 9.71 119.135 9.455 119.135 9.455 119.595 7.265 119.595 7.265 118.795 6.935 118.795 6.935 119.595 6.425 119.595 6.425 119.115 6.095 119.115 6.095 119.595 5.585 119.595 5.585 119.115 5.255 119.115 5.255 119.595 4.665 119.595 4.665 119.115 4.495 119.115 4.495 119.595 3.825 119.595 3.825 119.115 3.655 119.115 3.655 119.595 0 119.595 0 119.765 ;
      RECT 103.04 116.875 103.96 117.045 ;
      RECT 0 116.875 1.84 117.045 ;
      RECT 103.04 114.155 103.96 114.325 ;
      RECT 0 114.155 3.68 114.325 ;
      RECT 103.04 111.435 103.96 111.605 ;
      RECT 0 111.435 3.68 111.605 ;
      RECT 103.04 108.715 103.96 108.885 ;
      RECT 0 108.715 1.84 108.885 ;
      RECT 103.04 105.995 103.96 106.165 ;
      RECT 0 105.995 3.68 106.165 ;
      RECT 103.04 103.275 103.96 103.445 ;
      RECT 0 103.275 3.68 103.445 ;
      RECT 103.04 100.555 103.96 100.725 ;
      RECT 0 100.555 3.68 100.725 ;
      RECT 102.12 97.835 103.96 98.005 ;
      RECT 0 97.835 3.68 98.005 ;
      RECT 102.12 95.115 103.96 95.285 ;
      RECT 0 95.115 3.68 95.285 ;
      RECT 103.04 92.395 103.96 92.565 ;
      RECT 0 92.395 3.68 92.565 ;
      RECT 103.5 89.675 103.96 89.845 ;
      RECT 0 89.675 3.68 89.845 ;
      RECT 103.5 86.955 103.96 87.125 ;
      RECT 0 86.955 3.68 87.125 ;
      RECT 103.04 84.235 103.96 84.405 ;
      RECT 0 84.235 3.68 84.405 ;
      RECT 103.04 81.515 103.96 81.685 ;
      RECT 0 81.515 3.68 81.685 ;
      RECT 103.04 78.795 103.96 78.965 ;
      RECT 0 78.795 1.84 78.965 ;
      RECT 103.04 76.075 103.96 76.245 ;
      RECT 0 76.075 3.68 76.245 ;
      RECT 103.04 73.355 103.96 73.525 ;
      RECT 0 73.355 3.68 73.525 ;
      RECT 103.04 70.635 103.96 70.805 ;
      RECT 0 70.635 1.84 70.805 ;
      RECT 100.28 67.915 103.96 68.085 ;
      RECT 0 67.915 3.68 68.085 ;
      RECT 100.28 65.195 103.96 65.365 ;
      RECT 0 65.195 3.68 65.365 ;
      RECT 103.04 62.475 103.96 62.645 ;
      RECT 0 62.475 3.68 62.645 ;
      RECT 102.12 59.755 103.96 59.925 ;
      RECT 0 59.755 1.84 59.925 ;
      RECT 102.12 57.035 103.96 57.205 ;
      RECT 0 57.035 3.68 57.205 ;
      RECT 103.04 54.315 103.96 54.485 ;
      RECT 0 54.315 3.68 54.485 ;
      RECT 103.5 51.595 103.96 51.765 ;
      RECT 0 51.595 3.68 51.765 ;
      RECT 103.04 48.875 103.96 49.045 ;
      RECT 0 48.875 3.68 49.045 ;
      RECT 103.04 46.155 103.96 46.325 ;
      RECT 0 46.155 1.84 46.325 ;
      RECT 100.28 43.435 103.96 43.605 ;
      RECT 0 43.435 3.68 43.605 ;
      RECT 100.28 40.715 103.96 40.885 ;
      RECT 0 40.715 3.68 40.885 ;
      RECT 103.5 37.995 103.96 38.165 ;
      RECT 0 37.995 1.84 38.165 ;
      RECT 103.5 35.275 103.96 35.445 ;
      RECT 0 35.275 3.68 35.445 ;
      RECT 103.5 32.555 103.96 32.725 ;
      RECT 0 32.555 3.68 32.725 ;
      RECT 103.04 29.835 103.96 30.005 ;
      RECT 0 29.835 3.68 30.005 ;
      RECT 103.04 27.115 103.96 27.285 ;
      RECT 0 27.115 3.68 27.285 ;
      RECT 103.5 24.395 103.96 24.565 ;
      RECT 0 24.395 3.68 24.565 ;
      RECT 103.5 21.675 103.96 21.845 ;
      RECT 0 21.675 3.68 21.845 ;
      RECT 103.5 18.955 103.96 19.125 ;
      RECT 0 18.955 3.68 19.125 ;
      RECT 103.5 16.235 103.96 16.405 ;
      RECT 0 16.235 3.68 16.405 ;
      RECT 103.04 13.515 103.96 13.685 ;
      RECT 0 13.515 3.68 13.685 ;
      RECT 103.04 10.795 103.96 10.965 ;
      RECT 0 10.795 3.68 10.965 ;
      RECT 103.04 8.075 103.96 8.245 ;
      RECT 0 8.075 3.68 8.245 ;
      RECT 103.04 5.355 103.96 5.525 ;
      RECT 0 5.355 3.68 5.525 ;
      RECT 103.04 2.635 103.96 2.805 ;
      RECT 0 2.635 3.68 2.805 ;
      RECT 0 -0.085 103.96 0.085 ;
      POLYGON 103.79 124.95 103.79 0.17 0.17 0.17 0.17 119.51 30.53 119.51 30.53 124.95 ;
    LAYER via ;
      RECT 89.165 124.925 89.315 125.075 ;
      RECT 59.725 124.925 59.875 125.075 ;
      RECT 95.375 124.535 95.525 124.685 ;
      RECT 86.635 124.535 86.785 124.685 ;
      RECT 83.875 124.535 84.025 124.685 ;
      RECT 50.295 124.535 50.445 124.685 ;
      RECT 89.165 0.045 89.315 0.195 ;
      RECT 59.725 0.045 59.875 0.195 ;
    LAYER via2 ;
      RECT 89.14 124.9 89.34 125.1 ;
      RECT 59.7 124.9 59.9 125.1 ;
      RECT 58.09 124.68 58.29 124.88 ;
      RECT 42.91 124.68 43.11 124.88 ;
      RECT 36.93 124.68 37.13 124.88 ;
      RECT 89.14 0.02 89.34 0.22 ;
      RECT 59.7 0.02 59.9 0.22 ;
    LAYER via3 ;
      RECT 89.14 124.9 89.34 125.1 ;
      RECT 59.7 124.9 59.9 125.1 ;
      RECT 57.4 124.68 57.6 124.88 ;
      RECT 49.12 124.68 49.32 124.88 ;
      RECT 32.56 124.68 32.76 124.88 ;
      RECT 89.14 0.02 89.34 0.22 ;
      RECT 59.7 0.02 59.9 0.22 ;
    LAYER OVERLAP ;
      POLYGON 0 0 0 119.68 30.36 119.68 30.36 125.12 103.96 125.12 103.96 0 ;
  END
END sb_2__0_

END LIBRARY
