VERSION 5.7 ;
BUSBITCHARS "[]" ;

UNITS
  DATABASE MICRONS 1000 ;
END UNITS

MANUFACTURINGGRID 0.005 ;

LAYER nwell
  TYPE MASTERSLICE ;
END nwell

LAYER pwell
  TYPE MASTERSLICE ;
END pwell

LAYER fieldpoly
  TYPE MASTERSLICE ;
END fieldpoly

LAYER li1
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.46 ;
  WIDTH 0.17 ;
END li1

LAYER mcon
  TYPE CUT ;
END mcon

LAYER met1
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.34 ;
  WIDTH 0.14 ;
END met1

LAYER via
  TYPE CUT ;
END via

LAYER met2
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.46 ;
  WIDTH 0.14 ;
END met2

LAYER via2
  TYPE CUT ;
END via2

LAYER met3
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.68 ;
  WIDTH 0.3 ;
END met3

LAYER via3
  TYPE CUT ;
END via3

LAYER met4
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.92 ;
  WIDTH 0.3 ;
END met4

LAYER via4
  TYPE CUT ;
END via4

LAYER met5
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 3.4 ;
  WIDTH 1.6 ;
END met5

LAYER diff
  TYPE MASTERSLICE ;
END diff

LAYER licon1
  TYPE MASTERSLICE ;
END licon1

LAYER OVERLAP
  TYPE OVERLAP ;
END OVERLAP

VIA L1M1_PR
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.145 -0.115 0.145 0.115 ;
END L1M1_PR

VIA L1M1_PR_R
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.115 -0.145 0.115 0.145 ;
END L1M1_PR_R

VIA L1M1_PR_M
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.115 -0.145 0.115 0.145 ;
END L1M1_PR_M

VIA L1M1_PR_MR
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.145 -0.115 0.145 0.115 ;
END L1M1_PR_MR

VIA L1M1_PR_C
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.145 -0.145 0.145 0.145 ;
END L1M1_PR_C

VIA M1M2_PR
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR

VIA M1M2_PR_Enc
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_Enc

VIA M1M2_PR_R
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_R

VIA M1M2_PR_R_Enc
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR_R_Enc

VIA M1M2_PR_M
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_M

VIA M1M2_PR_M_Enc
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR_M_Enc

VIA M1M2_PR_MR
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR_MR

VIA M1M2_PR_MR_Enc
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_MR_Enc

VIA M1M2_PR_C
  LAYER met1 ;
    RECT -0.16 -0.16 0.16 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.16 0.16 0.16 ;
END M1M2_PR_C

VIA M2M3_PR
  LAYER met2 ;
    RECT -0.14 -0.185 0.14 0.185 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR

VIA M2M3_PR_R
  LAYER met2 ;
    RECT -0.185 -0.14 0.185 0.14 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_R

VIA M2M3_PR_M
  LAYER met2 ;
    RECT -0.14 -0.185 0.14 0.185 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_M

VIA M2M3_PR_MR
  LAYER met2 ;
    RECT -0.185 -0.14 0.185 0.14 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_MR

VIA M2M3_PR_C
  LAYER met2 ;
    RECT -0.185 -0.185 0.185 0.185 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_C

VIA M3M4_PR
  LAYER met3 ;
    RECT -0.19 -0.16 0.19 0.16 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR

VIA M3M4_PR_R
  LAYER met3 ;
    RECT -0.16 -0.19 0.16 0.19 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_R

VIA M3M4_PR_M
  LAYER met3 ;
    RECT -0.19 -0.16 0.19 0.16 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_M

VIA M3M4_PR_MR
  LAYER met3 ;
    RECT -0.16 -0.19 0.16 0.19 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_MR

VIA M3M4_PR_C
  LAYER met3 ;
    RECT -0.19 -0.19 0.19 0.19 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_C

VIA M4M5_PR
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR

VIA M4M5_PR_R
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_R

VIA M4M5_PR_M
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_M

VIA M4M5_PR_MR
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_MR

VIA M4M5_PR_C
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_C

SITE unit
  CLASS CORE ;
  SYMMETRY Y ;
  SIZE 0.46 BY 2.72 ;
END unit

SITE unithddbl
  CLASS CORE ;
  SIZE 0.46 BY 5.44 ;
END unithddbl

MACRO sb_0__2_
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  SIZE 84.64 BY 81.6 ;
  SYMMETRY X Y ;
  PIN prog_clk[0]
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER met3 ;
        RECT 83.26 19.57 84.64 19.87 ;
    END
  END prog_clk[0]
  PIN chanx_right_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 83.26 61.05 84.64 61.35 ;
    END
  END chanx_right_in[0]
  PIN chanx_right_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 83.26 39.29 84.64 39.59 ;
    END
  END chanx_right_in[1]
  PIN chanx_right_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 83.26 74.65 84.64 74.95 ;
    END
  END chanx_right_in[2]
  PIN chanx_right_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 83.26 56.97 84.64 57.27 ;
    END
  END chanx_right_in[3]
  PIN chanx_right_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 83.26 63.77 84.64 64.07 ;
    END
  END chanx_right_in[4]
  PIN chanx_right_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 83.26 69.21 84.64 69.51 ;
    END
  END chanx_right_in[5]
  PIN chanx_right_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 83.26 22.97 84.64 23.27 ;
    END
  END chanx_right_in[6]
  PIN chanx_right_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 83.26 73.29 84.64 73.59 ;
    END
  END chanx_right_in[7]
  PIN chanx_right_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 83.26 66.49 84.64 66.79 ;
    END
  END chanx_right_in[8]
  PIN chanx_right_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 83.26 21.61 84.64 21.91 ;
    END
  END chanx_right_in[9]
  PIN chanx_right_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 83.26 62.41 84.64 62.71 ;
    END
  END chanx_right_in[10]
  PIN chanx_right_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 83.26 36.57 84.64 36.87 ;
    END
  END chanx_right_in[11]
  PIN chanx_right_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 83.26 59.69 84.64 59.99 ;
    END
  END chanx_right_in[12]
  PIN chanx_right_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 83.26 43.37 84.64 43.67 ;
    END
  END chanx_right_in[13]
  PIN chanx_right_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 83.26 35.21 84.64 35.51 ;
    END
  END chanx_right_in[14]
  PIN chanx_right_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 83.26 55.61 84.64 55.91 ;
    END
  END chanx_right_in[15]
  PIN chanx_right_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 83.26 67.85 84.64 68.15 ;
    END
  END chanx_right_in[16]
  PIN chanx_right_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 83.26 44.73 84.64 45.03 ;
    END
  END chanx_right_in[17]
  PIN chanx_right_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 83.26 33.85 84.64 34.15 ;
    END
  END chanx_right_in[18]
  PIN chanx_right_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 83.26 40.65 84.64 40.95 ;
    END
  END chanx_right_in[19]
  PIN right_top_grid_pin_1_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.35 80.24 81.49 81.6 ;
    END
  END right_top_grid_pin_1_[0]
  PIN chany_bottom_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.89 0 35.03 1.36 ;
    END
  END chany_bottom_in[0]
  PIN chany_bottom_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.77 0 24.91 1.36 ;
    END
  END chany_bottom_in[1]
  PIN chany_bottom_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.75 0 53.89 1.36 ;
    END
  END chany_bottom_in[2]
  PIN chany_bottom_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.73 0 36.87 1.36 ;
    END
  END chany_bottom_in[3]
  PIN chany_bottom_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 56.89 0 57.19 1.36 ;
    END
  END chany_bottom_in[4]
  PIN chany_bottom_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.83 0 52.97 1.36 ;
    END
  END chany_bottom_in[5]
  PIN chany_bottom_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.17 0 43.31 1.36 ;
    END
  END chany_bottom_in[6]
  PIN chany_bottom_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.05 0 10.19 1.36 ;
    END
  END chany_bottom_in[7]
  PIN chany_bottom_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.25 0 42.39 1.36 ;
    END
  END chany_bottom_in[8]
  PIN chany_bottom_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.21 0 8.35 1.36 ;
    END
  END chany_bottom_in[9]
  PIN chany_bottom_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.09 0 21.23 1.36 ;
    END
  END chany_bottom_in[10]
  PIN chany_bottom_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.65 0 37.79 1.36 ;
    END
  END chany_bottom_in[11]
  PIN chany_bottom_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.35 0 58.49 1.36 ;
    END
  END chany_bottom_in[12]
  PIN chany_bottom_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.49 0 39.63 1.36 ;
    END
  END chany_bottom_in[13]
  PIN chany_bottom_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.43 0 57.57 1.36 ;
    END
  END chany_bottom_in[14]
  PIN chany_bottom_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.13 0 9.27 1.36 ;
    END
  END chany_bottom_in[15]
  PIN chany_bottom_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.45 0 28.59 1.36 ;
    END
  END chany_bottom_in[16]
  PIN chany_bottom_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.17 0 20.31 1.36 ;
    END
  END chany_bottom_in[17]
  PIN chany_bottom_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.25 0 19.39 1.36 ;
    END
  END chany_bottom_in[18]
  PIN chany_bottom_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.29 0 30.43 1.36 ;
    END
  END chany_bottom_in[19]
  PIN bottom_left_grid_pin_1_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.15 0 3.29 1.36 ;
    END
  END bottom_left_grid_pin_1_[0]
  PIN ccff_head[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.27 80.24 82.41 81.6 ;
    END
  END ccff_head[0]
  PIN chanx_right_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 83.26 58.33 84.64 58.63 ;
    END
  END chanx_right_out[0]
  PIN chanx_right_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 83.26 70.57 84.64 70.87 ;
    END
  END chanx_right_out[1]
  PIN chanx_right_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 83.26 65.13 84.64 65.43 ;
    END
  END chanx_right_out[2]
  PIN chanx_right_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 83.26 47.45 84.64 47.75 ;
    END
  END chanx_right_out[3]
  PIN chanx_right_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 83.26 42.01 84.64 42.31 ;
    END
  END chanx_right_out[4]
  PIN chanx_right_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 83.26 25.69 84.64 25.99 ;
    END
  END chanx_right_out[5]
  PIN chanx_right_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 83.26 32.49 84.64 32.79 ;
    END
  END chanx_right_out[6]
  PIN chanx_right_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 83.26 54.25 84.64 54.55 ;
    END
  END chanx_right_out[7]
  PIN chanx_right_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 83.26 71.93 84.64 72.23 ;
    END
  END chanx_right_out[8]
  PIN chanx_right_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 83.26 48.81 84.64 49.11 ;
    END
  END chanx_right_out[9]
  PIN chanx_right_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 83.26 24.33 84.64 24.63 ;
    END
  END chanx_right_out[10]
  PIN chanx_right_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 83.26 52.89 84.64 53.19 ;
    END
  END chanx_right_out[11]
  PIN chanx_right_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 83.26 37.93 84.64 38.23 ;
    END
  END chanx_right_out[12]
  PIN chanx_right_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 83.26 27.05 84.64 27.35 ;
    END
  END chanx_right_out[13]
  PIN chanx_right_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 83.26 31.13 84.64 31.43 ;
    END
  END chanx_right_out[14]
  PIN chanx_right_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 83.26 50.17 84.64 50.47 ;
    END
  END chanx_right_out[15]
  PIN chanx_right_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 83.26 46.09 84.64 46.39 ;
    END
  END chanx_right_out[16]
  PIN chanx_right_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 83.26 51.53 84.64 51.83 ;
    END
  END chanx_right_out[17]
  PIN chanx_right_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 83.26 28.41 84.64 28.71 ;
    END
  END chanx_right_out[18]
  PIN chanx_right_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 83.26 29.77 84.64 30.07 ;
    END
  END chanx_right_out[19]
  PIN chany_bottom_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.41 0 40.55 1.36 ;
    END
  END chany_bottom_out[0]
  PIN chany_bottom_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.67 0 54.81 1.36 ;
    END
  END chany_bottom_out[1]
  PIN chany_bottom_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.37 0 29.51 1.36 ;
    END
  END chany_bottom_out[2]
  PIN chany_bottom_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.97 0 34.11 1.36 ;
    END
  END chany_bottom_out[3]
  PIN chany_bottom_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.21 0 31.35 1.36 ;
    END
  END chany_bottom_out[4]
  PIN chany_bottom_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.57 0 38.71 1.36 ;
    END
  END chany_bottom_out[5]
  PIN chany_bottom_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.97 0 11.11 1.36 ;
    END
  END chany_bottom_out[6]
  PIN chany_bottom_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.49 0 16.63 1.36 ;
    END
  END chany_bottom_out[7]
  PIN chany_bottom_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.81 0 35.95 1.36 ;
    END
  END chany_bottom_out[8]
  PIN chany_bottom_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.89 0 12.03 1.36 ;
    END
  END chany_bottom_out[9]
  PIN chany_bottom_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.59 0 55.73 1.36 ;
    END
  END chany_bottom_out[10]
  PIN chany_bottom_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.05 0 33.19 1.36 ;
    END
  END chany_bottom_out[11]
  PIN chany_bottom_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.41 0 17.55 1.36 ;
    END
  END chany_bottom_out[12]
  PIN chany_bottom_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.51 0 56.65 1.36 ;
    END
  END chany_bottom_out[13]
  PIN chany_bottom_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.57 0 15.71 1.36 ;
    END
  END chany_bottom_out[14]
  PIN chany_bottom_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.81 0 12.95 1.36 ;
    END
  END chany_bottom_out[15]
  PIN chany_bottom_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.33 0 41.47 1.36 ;
    END
  END chany_bottom_out[16]
  PIN chany_bottom_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.13 0 32.27 1.36 ;
    END
  END chany_bottom_out[17]
  PIN chany_bottom_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.65 0 14.79 1.36 ;
    END
  END chany_bottom_out[18]
  PIN chany_bottom_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.73 0 13.87 1.36 ;
    END
  END chany_bottom_out[19]
  PIN ccff_tail[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.33 0 18.47 1.36 ;
    END
  END ccff_tail[0]
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
  END VDD
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
  END VSS
  OBS
    LAYER li1 ;
      RECT 0 81.515 84.64 81.685 ;
      RECT 84.18 78.795 84.64 78.965 ;
      RECT 0 78.795 3.68 78.965 ;
      RECT 83.72 76.075 84.64 76.245 ;
      RECT 0 76.075 3.68 76.245 ;
      RECT 83.72 73.355 84.64 73.525 ;
      RECT 0 73.355 3.68 73.525 ;
      RECT 83.72 70.635 84.64 70.805 ;
      RECT 0 70.635 3.68 70.805 ;
      RECT 83.72 67.915 84.64 68.085 ;
      RECT 0 67.915 3.68 68.085 ;
      RECT 80.96 65.195 84.64 65.365 ;
      RECT 0 65.195 3.68 65.365 ;
      RECT 80.96 62.475 84.64 62.645 ;
      RECT 0 62.475 3.68 62.645 ;
      RECT 80.96 59.755 84.64 59.925 ;
      RECT 0 59.755 3.68 59.925 ;
      RECT 83.72 57.035 84.64 57.205 ;
      RECT 0 57.035 3.68 57.205 ;
      RECT 83.72 54.315 84.64 54.485 ;
      RECT 0 54.315 3.68 54.485 ;
      RECT 83.72 51.595 84.64 51.765 ;
      RECT 0 51.595 3.68 51.765 ;
      RECT 83.72 48.875 84.64 49.045 ;
      RECT 0 48.875 3.68 49.045 ;
      RECT 83.72 46.155 84.64 46.325 ;
      RECT 0 46.155 3.68 46.325 ;
      RECT 83.72 43.435 84.64 43.605 ;
      RECT 0 43.435 3.68 43.605 ;
      RECT 83.72 40.715 84.64 40.885 ;
      RECT 0 40.715 3.68 40.885 ;
      RECT 83.72 37.995 84.64 38.165 ;
      RECT 0 37.995 3.68 38.165 ;
      RECT 83.72 35.275 84.64 35.445 ;
      RECT 0 35.275 3.68 35.445 ;
      RECT 83.72 32.555 84.64 32.725 ;
      RECT 0 32.555 3.68 32.725 ;
      RECT 83.72 29.835 84.64 30.005 ;
      RECT 0 29.835 3.68 30.005 ;
      RECT 83.72 27.115 84.64 27.285 ;
      RECT 0 27.115 3.68 27.285 ;
      RECT 83.72 24.395 84.64 24.565 ;
      RECT 0 24.395 3.68 24.565 ;
      RECT 83.72 21.675 84.64 21.845 ;
      RECT 0 21.675 3.68 21.845 ;
      RECT 83.72 18.955 84.64 19.125 ;
      RECT 0 18.955 3.68 19.125 ;
      RECT 65.78 16.235 84.64 16.405 ;
      RECT 0 16.235 3.68 16.405 ;
      RECT 65.78 13.515 66.24 13.685 ;
      RECT 0 13.515 3.68 13.685 ;
      RECT 65.32 10.795 66.24 10.965 ;
      RECT 0 10.795 3.68 10.965 ;
      RECT 65.32 8.075 66.24 8.245 ;
      RECT 0 8.075 3.68 8.245 ;
      RECT 62.56 5.355 66.24 5.525 ;
      RECT 0 5.355 3.68 5.525 ;
      RECT 62.56 2.635 66.24 2.805 ;
      RECT 0 2.635 3.68 2.805 ;
      RECT 0 -0.085 66.24 0.085 ;
    LAYER met3 ;
      POLYGON 83.425 72.925 83.425 72.595 83.095 72.595 83.095 72.61 79.89 72.61 79.89 72.91 83.095 72.91 83.095 72.925 ;
      POLYGON 82.86 55.23 82.86 55.21 83.41 55.21 83.41 54.93 58.27 54.93 58.27 55.23 ;
      POLYGON 82.95 32.11 82.95 31.83 82.86 31.83 82.86 31.13 82.65 31.13 82.65 31.81 80.35 31.81 80.35 32.11 ;
      POLYGON 84.24 81.2 84.24 75.35 82.86 75.35 82.86 74.25 84.24 74.25 84.24 73.99 82.86 73.99 82.86 72.89 84.24 72.89 84.24 72.63 82.86 72.63 82.86 71.53 84.24 71.53 84.24 71.27 82.86 71.27 82.86 70.17 84.24 70.17 84.24 69.91 82.86 69.91 82.86 68.81 84.24 68.81 84.24 68.55 82.86 68.55 82.86 67.45 84.24 67.45 84.24 67.19 82.86 67.19 82.86 66.09 84.24 66.09 84.24 65.83 82.86 65.83 82.86 64.73 84.24 64.73 84.24 64.47 82.86 64.47 82.86 63.37 84.24 63.37 84.24 63.11 82.86 63.11 82.86 62.01 84.24 62.01 84.24 61.75 82.86 61.75 82.86 60.65 84.24 60.65 84.24 60.39 82.86 60.39 82.86 59.29 84.24 59.29 84.24 59.03 82.86 59.03 82.86 57.93 84.24 57.93 84.24 57.67 82.86 57.67 82.86 56.57 84.24 56.57 84.24 56.31 82.86 56.31 82.86 55.21 84.24 55.21 84.24 54.95 82.86 54.95 82.86 53.85 84.24 53.85 84.24 53.59 82.86 53.59 82.86 52.49 84.24 52.49 84.24 52.23 82.86 52.23 82.86 51.13 84.24 51.13 84.24 50.87 82.86 50.87 82.86 49.77 84.24 49.77 84.24 49.51 82.86 49.51 82.86 48.41 84.24 48.41 84.24 48.15 82.86 48.15 82.86 47.05 84.24 47.05 84.24 46.79 82.86 46.79 82.86 45.69 84.24 45.69 84.24 45.43 82.86 45.43 82.86 44.33 84.24 44.33 84.24 44.07 82.86 44.07 82.86 42.97 84.24 42.97 84.24 42.71 82.86 42.71 82.86 41.61 84.24 41.61 84.24 41.35 82.86 41.35 82.86 40.25 84.24 40.25 84.24 39.99 82.86 39.99 82.86 38.89 84.24 38.89 84.24 38.63 82.86 38.63 82.86 37.53 84.24 37.53 84.24 37.27 82.86 37.27 82.86 36.17 84.24 36.17 84.24 35.91 82.86 35.91 82.86 34.81 84.24 34.81 84.24 34.55 82.86 34.55 82.86 33.45 84.24 33.45 84.24 33.19 82.86 33.19 82.86 32.09 84.24 32.09 84.24 31.83 82.86 31.83 82.86 30.73 84.24 30.73 84.24 30.47 82.86 30.47 82.86 29.37 84.24 29.37 84.24 29.11 82.86 29.11 82.86 28.01 84.24 28.01 84.24 27.75 82.86 27.75 82.86 26.65 84.24 26.65 84.24 26.39 82.86 26.39 82.86 25.29 84.24 25.29 84.24 25.03 82.86 25.03 82.86 23.93 84.24 23.93 84.24 23.67 82.86 23.67 82.86 22.57 84.24 22.57 84.24 22.31 82.86 22.31 82.86 21.21 84.24 21.21 84.24 20.27 82.86 20.27 82.86 19.17 84.24 19.17 84.24 16.72 65.84 16.72 65.84 0.4 0.4 0.4 0.4 81.2 ;
    LAYER met2 ;
      RECT 38.05 1.54 38.31 1.86 ;
      RECT 19.65 1.54 19.91 1.86 ;
      POLYGON 84.36 81.32 84.36 16.6 65.96 16.6 65.96 0.28 58.77 0.28 58.77 1.64 58.07 1.64 58.07 0.28 57.85 0.28 57.85 1.64 57.15 1.64 57.15 0.28 56.93 0.28 56.93 1.64 56.23 1.64 56.23 0.28 56.01 0.28 56.01 1.64 55.31 1.64 55.31 0.28 55.09 0.28 55.09 1.64 54.39 1.64 54.39 0.28 54.17 0.28 54.17 1.64 53.47 1.64 53.47 0.28 53.25 0.28 53.25 1.64 52.55 1.64 52.55 0.28 43.59 0.28 43.59 1.64 42.89 1.64 42.89 0.28 42.67 0.28 42.67 1.64 41.97 1.64 41.97 0.28 41.75 0.28 41.75 1.64 41.05 1.64 41.05 0.28 40.83 0.28 40.83 1.64 40.13 1.64 40.13 0.28 39.91 0.28 39.91 1.64 39.21 1.64 39.21 0.28 38.99 0.28 38.99 1.64 38.29 1.64 38.29 0.28 38.07 0.28 38.07 1.64 37.37 1.64 37.37 0.28 37.15 0.28 37.15 1.64 36.45 1.64 36.45 0.28 36.23 0.28 36.23 1.64 35.53 1.64 35.53 0.28 35.31 0.28 35.31 1.64 34.61 1.64 34.61 0.28 34.39 0.28 34.39 1.64 33.69 1.64 33.69 0.28 33.47 0.28 33.47 1.64 32.77 1.64 32.77 0.28 32.55 0.28 32.55 1.64 31.85 1.64 31.85 0.28 31.63 0.28 31.63 1.64 30.93 1.64 30.93 0.28 30.71 0.28 30.71 1.64 30.01 1.64 30.01 0.28 29.79 0.28 29.79 1.64 29.09 1.64 29.09 0.28 28.87 0.28 28.87 1.64 28.17 1.64 28.17 0.28 25.19 0.28 25.19 1.64 24.49 1.64 24.49 0.28 21.51 0.28 21.51 1.64 20.81 1.64 20.81 0.28 20.59 0.28 20.59 1.64 19.89 1.64 19.89 0.28 19.67 0.28 19.67 1.64 18.97 1.64 18.97 0.28 18.75 0.28 18.75 1.64 18.05 1.64 18.05 0.28 17.83 0.28 17.83 1.64 17.13 1.64 17.13 0.28 16.91 0.28 16.91 1.64 16.21 1.64 16.21 0.28 15.99 0.28 15.99 1.64 15.29 1.64 15.29 0.28 15.07 0.28 15.07 1.64 14.37 1.64 14.37 0.28 14.15 0.28 14.15 1.64 13.45 1.64 13.45 0.28 13.23 0.28 13.23 1.64 12.53 1.64 12.53 0.28 12.31 0.28 12.31 1.64 11.61 1.64 11.61 0.28 11.39 0.28 11.39 1.64 10.69 1.64 10.69 0.28 10.47 0.28 10.47 1.64 9.77 1.64 9.77 0.28 9.55 0.28 9.55 1.64 8.85 1.64 8.85 0.28 8.63 0.28 8.63 1.64 7.93 1.64 7.93 0.28 3.57 0.28 3.57 1.64 2.87 1.64 2.87 0.28 0.28 0.28 0.28 81.32 81.07 81.32 81.07 79.96 81.77 79.96 81.77 81.32 81.99 81.32 81.99 79.96 82.69 79.96 82.69 81.32 ;
    LAYER met4 ;
      POLYGON 84.24 81.2 84.24 16.72 65.84 16.72 65.84 0.4 57.59 0.4 57.59 1.76 56.49 1.76 56.49 0.4 0.4 0.4 0.4 81.2 ;
    LAYER li1 ;
      RECT 65.865 80.79 66.615 81.335 ;
      RECT 17.105 80.79 17.855 81.335 ;
      RECT 65.865 16.585 66.615 17.13 ;
      RECT 17.105 0.265 17.855 0.81 ;
      POLYGON 84.3 81.26 84.3 16.66 65.9 16.66 65.9 0.34 0.34 0.34 0.34 81.26 ;
    LAYER met1 ;
      RECT 0 81.36 84.64 81.84 ;
      RECT 84.18 78.64 84.64 79.12 ;
      RECT 0 78.64 3.68 79.12 ;
      RECT 83.72 75.92 84.64 76.4 ;
      RECT 0 75.92 3.68 76.4 ;
      RECT 83.72 73.2 84.64 73.68 ;
      RECT 0 73.2 3.68 73.68 ;
      RECT 83.72 70.48 84.64 70.96 ;
      RECT 0 70.48 3.68 70.96 ;
      RECT 83.72 67.76 84.64 68.24 ;
      RECT 0 67.76 3.68 68.24 ;
      RECT 80.96 65.04 84.64 65.52 ;
      RECT 0 65.04 3.68 65.52 ;
      RECT 80.96 62.32 84.64 62.8 ;
      RECT 0 62.32 3.68 62.8 ;
      RECT 80.96 59.6 84.64 60.08 ;
      RECT 0 59.6 3.68 60.08 ;
      RECT 83.72 56.88 84.64 57.36 ;
      RECT 0 56.88 3.68 57.36 ;
      RECT 83.72 54.16 84.64 54.64 ;
      RECT 0 54.16 3.68 54.64 ;
      RECT 83.72 51.44 84.64 51.92 ;
      RECT 0 51.44 3.68 51.92 ;
      RECT 83.72 48.72 84.64 49.2 ;
      RECT 0 48.72 3.68 49.2 ;
      RECT 83.72 46 84.64 46.48 ;
      RECT 0 46 3.68 46.48 ;
      RECT 83.72 43.28 84.64 43.76 ;
      RECT 0 43.28 3.68 43.76 ;
      RECT 83.72 40.56 84.64 41.04 ;
      RECT 0 40.56 3.68 41.04 ;
      RECT 83.72 37.84 84.64 38.32 ;
      RECT 0 37.84 3.68 38.32 ;
      RECT 83.72 35.12 84.64 35.6 ;
      RECT 0 35.12 3.68 35.6 ;
      RECT 83.72 32.4 84.64 32.88 ;
      RECT 0 32.4 3.68 32.88 ;
      RECT 83.72 29.68 84.64 30.16 ;
      RECT 0 29.68 3.68 30.16 ;
      RECT 83.72 26.96 84.64 27.44 ;
      RECT 0 26.96 3.68 27.44 ;
      RECT 83.72 24.24 84.64 24.72 ;
      RECT 0 24.24 3.68 24.72 ;
      RECT 83.72 21.52 84.64 22 ;
      RECT 0 21.52 3.68 22 ;
      RECT 83.72 18.8 84.64 19.28 ;
      RECT 0 18.8 3.68 19.28 ;
      RECT 65.78 16.08 84.64 16.56 ;
      RECT 0 16.08 3.68 16.56 ;
      RECT 65.78 13.36 66.24 13.84 ;
      RECT 0 13.36 3.68 13.84 ;
      RECT 65.32 10.64 66.24 11.12 ;
      RECT 0 10.64 3.68 11.12 ;
      RECT 65.32 7.92 66.24 8.4 ;
      RECT 0 7.92 3.68 8.4 ;
      RECT 62.56 5.2 66.24 5.68 ;
      RECT 0 5.2 3.68 5.68 ;
      RECT 62.56 2.48 66.24 2.96 ;
      RECT 0 2.48 3.68 2.96 ;
      RECT 0 -0.24 66.24 0.24 ;
      POLYGON 84.36 81.32 84.36 16.6 65.96 16.6 65.96 0.28 0.28 0.28 0.28 81.32 ;
    LAYER met5 ;
      POLYGON 81.44 78.4 81.44 19.52 63.04 19.52 63.04 3.2 3.2 3.2 3.2 78.4 ;
    LAYER mcon ;
      RECT 84.325 81.515 84.495 81.685 ;
      RECT 83.865 81.515 84.035 81.685 ;
      RECT 83.405 81.515 83.575 81.685 ;
      RECT 82.945 81.515 83.115 81.685 ;
      RECT 82.485 81.515 82.655 81.685 ;
      RECT 82.025 81.515 82.195 81.685 ;
      RECT 81.565 81.515 81.735 81.685 ;
      RECT 81.105 81.515 81.275 81.685 ;
      RECT 80.645 81.515 80.815 81.685 ;
      RECT 80.185 81.515 80.355 81.685 ;
      RECT 79.725 81.515 79.895 81.685 ;
      RECT 79.265 81.515 79.435 81.685 ;
      RECT 78.805 81.515 78.975 81.685 ;
      RECT 78.345 81.515 78.515 81.685 ;
      RECT 77.885 81.515 78.055 81.685 ;
      RECT 77.425 81.515 77.595 81.685 ;
      RECT 76.965 81.515 77.135 81.685 ;
      RECT 76.505 81.515 76.675 81.685 ;
      RECT 76.045 81.515 76.215 81.685 ;
      RECT 75.585 81.515 75.755 81.685 ;
      RECT 75.125 81.515 75.295 81.685 ;
      RECT 74.665 81.515 74.835 81.685 ;
      RECT 74.205 81.515 74.375 81.685 ;
      RECT 73.745 81.515 73.915 81.685 ;
      RECT 73.285 81.515 73.455 81.685 ;
      RECT 72.825 81.515 72.995 81.685 ;
      RECT 72.365 81.515 72.535 81.685 ;
      RECT 71.905 81.515 72.075 81.685 ;
      RECT 71.445 81.515 71.615 81.685 ;
      RECT 70.985 81.515 71.155 81.685 ;
      RECT 70.525 81.515 70.695 81.685 ;
      RECT 70.065 81.515 70.235 81.685 ;
      RECT 69.605 81.515 69.775 81.685 ;
      RECT 69.145 81.515 69.315 81.685 ;
      RECT 68.685 81.515 68.855 81.685 ;
      RECT 68.225 81.515 68.395 81.685 ;
      RECT 67.765 81.515 67.935 81.685 ;
      RECT 67.305 81.515 67.475 81.685 ;
      RECT 66.845 81.515 67.015 81.685 ;
      RECT 66.385 81.515 66.555 81.685 ;
      RECT 65.925 81.515 66.095 81.685 ;
      RECT 65.465 81.515 65.635 81.685 ;
      RECT 65.005 81.515 65.175 81.685 ;
      RECT 64.545 81.515 64.715 81.685 ;
      RECT 64.085 81.515 64.255 81.685 ;
      RECT 63.625 81.515 63.795 81.685 ;
      RECT 63.165 81.515 63.335 81.685 ;
      RECT 62.705 81.515 62.875 81.685 ;
      RECT 62.245 81.515 62.415 81.685 ;
      RECT 61.785 81.515 61.955 81.685 ;
      RECT 61.325 81.515 61.495 81.685 ;
      RECT 60.865 81.515 61.035 81.685 ;
      RECT 60.405 81.515 60.575 81.685 ;
      RECT 59.945 81.515 60.115 81.685 ;
      RECT 59.485 81.515 59.655 81.685 ;
      RECT 59.025 81.515 59.195 81.685 ;
      RECT 58.565 81.515 58.735 81.685 ;
      RECT 58.105 81.515 58.275 81.685 ;
      RECT 57.645 81.515 57.815 81.685 ;
      RECT 57.185 81.515 57.355 81.685 ;
      RECT 56.725 81.515 56.895 81.685 ;
      RECT 56.265 81.515 56.435 81.685 ;
      RECT 55.805 81.515 55.975 81.685 ;
      RECT 55.345 81.515 55.515 81.685 ;
      RECT 54.885 81.515 55.055 81.685 ;
      RECT 54.425 81.515 54.595 81.685 ;
      RECT 53.965 81.515 54.135 81.685 ;
      RECT 53.505 81.515 53.675 81.685 ;
      RECT 53.045 81.515 53.215 81.685 ;
      RECT 52.585 81.515 52.755 81.685 ;
      RECT 52.125 81.515 52.295 81.685 ;
      RECT 51.665 81.515 51.835 81.685 ;
      RECT 51.205 81.515 51.375 81.685 ;
      RECT 50.745 81.515 50.915 81.685 ;
      RECT 50.285 81.515 50.455 81.685 ;
      RECT 49.825 81.515 49.995 81.685 ;
      RECT 49.365 81.515 49.535 81.685 ;
      RECT 48.905 81.515 49.075 81.685 ;
      RECT 48.445 81.515 48.615 81.685 ;
      RECT 47.985 81.515 48.155 81.685 ;
      RECT 47.525 81.515 47.695 81.685 ;
      RECT 47.065 81.515 47.235 81.685 ;
      RECT 46.605 81.515 46.775 81.685 ;
      RECT 46.145 81.515 46.315 81.685 ;
      RECT 45.685 81.515 45.855 81.685 ;
      RECT 45.225 81.515 45.395 81.685 ;
      RECT 44.765 81.515 44.935 81.685 ;
      RECT 44.305 81.515 44.475 81.685 ;
      RECT 43.845 81.515 44.015 81.685 ;
      RECT 43.385 81.515 43.555 81.685 ;
      RECT 42.925 81.515 43.095 81.685 ;
      RECT 42.465 81.515 42.635 81.685 ;
      RECT 42.005 81.515 42.175 81.685 ;
      RECT 41.545 81.515 41.715 81.685 ;
      RECT 41.085 81.515 41.255 81.685 ;
      RECT 40.625 81.515 40.795 81.685 ;
      RECT 40.165 81.515 40.335 81.685 ;
      RECT 39.705 81.515 39.875 81.685 ;
      RECT 39.245 81.515 39.415 81.685 ;
      RECT 38.785 81.515 38.955 81.685 ;
      RECT 38.325 81.515 38.495 81.685 ;
      RECT 37.865 81.515 38.035 81.685 ;
      RECT 37.405 81.515 37.575 81.685 ;
      RECT 36.945 81.515 37.115 81.685 ;
      RECT 36.485 81.515 36.655 81.685 ;
      RECT 36.025 81.515 36.195 81.685 ;
      RECT 35.565 81.515 35.735 81.685 ;
      RECT 35.105 81.515 35.275 81.685 ;
      RECT 34.645 81.515 34.815 81.685 ;
      RECT 34.185 81.515 34.355 81.685 ;
      RECT 33.725 81.515 33.895 81.685 ;
      RECT 33.265 81.515 33.435 81.685 ;
      RECT 32.805 81.515 32.975 81.685 ;
      RECT 32.345 81.515 32.515 81.685 ;
      RECT 31.885 81.515 32.055 81.685 ;
      RECT 31.425 81.515 31.595 81.685 ;
      RECT 30.965 81.515 31.135 81.685 ;
      RECT 30.505 81.515 30.675 81.685 ;
      RECT 30.045 81.515 30.215 81.685 ;
      RECT 29.585 81.515 29.755 81.685 ;
      RECT 29.125 81.515 29.295 81.685 ;
      RECT 28.665 81.515 28.835 81.685 ;
      RECT 28.205 81.515 28.375 81.685 ;
      RECT 27.745 81.515 27.915 81.685 ;
      RECT 27.285 81.515 27.455 81.685 ;
      RECT 26.825 81.515 26.995 81.685 ;
      RECT 26.365 81.515 26.535 81.685 ;
      RECT 25.905 81.515 26.075 81.685 ;
      RECT 25.445 81.515 25.615 81.685 ;
      RECT 24.985 81.515 25.155 81.685 ;
      RECT 24.525 81.515 24.695 81.685 ;
      RECT 24.065 81.515 24.235 81.685 ;
      RECT 23.605 81.515 23.775 81.685 ;
      RECT 23.145 81.515 23.315 81.685 ;
      RECT 22.685 81.515 22.855 81.685 ;
      RECT 22.225 81.515 22.395 81.685 ;
      RECT 21.765 81.515 21.935 81.685 ;
      RECT 21.305 81.515 21.475 81.685 ;
      RECT 20.845 81.515 21.015 81.685 ;
      RECT 20.385 81.515 20.555 81.685 ;
      RECT 19.925 81.515 20.095 81.685 ;
      RECT 19.465 81.515 19.635 81.685 ;
      RECT 19.005 81.515 19.175 81.685 ;
      RECT 18.545 81.515 18.715 81.685 ;
      RECT 18.085 81.515 18.255 81.685 ;
      RECT 17.625 81.515 17.795 81.685 ;
      RECT 17.165 81.515 17.335 81.685 ;
      RECT 16.705 81.515 16.875 81.685 ;
      RECT 16.245 81.515 16.415 81.685 ;
      RECT 15.785 81.515 15.955 81.685 ;
      RECT 15.325 81.515 15.495 81.685 ;
      RECT 14.865 81.515 15.035 81.685 ;
      RECT 14.405 81.515 14.575 81.685 ;
      RECT 13.945 81.515 14.115 81.685 ;
      RECT 13.485 81.515 13.655 81.685 ;
      RECT 13.025 81.515 13.195 81.685 ;
      RECT 12.565 81.515 12.735 81.685 ;
      RECT 12.105 81.515 12.275 81.685 ;
      RECT 11.645 81.515 11.815 81.685 ;
      RECT 11.185 81.515 11.355 81.685 ;
      RECT 10.725 81.515 10.895 81.685 ;
      RECT 10.265 81.515 10.435 81.685 ;
      RECT 9.805 81.515 9.975 81.685 ;
      RECT 9.345 81.515 9.515 81.685 ;
      RECT 8.885 81.515 9.055 81.685 ;
      RECT 8.425 81.515 8.595 81.685 ;
      RECT 7.965 81.515 8.135 81.685 ;
      RECT 7.505 81.515 7.675 81.685 ;
      RECT 7.045 81.515 7.215 81.685 ;
      RECT 6.585 81.515 6.755 81.685 ;
      RECT 6.125 81.515 6.295 81.685 ;
      RECT 5.665 81.515 5.835 81.685 ;
      RECT 5.205 81.515 5.375 81.685 ;
      RECT 4.745 81.515 4.915 81.685 ;
      RECT 4.285 81.515 4.455 81.685 ;
      RECT 3.825 81.515 3.995 81.685 ;
      RECT 3.365 81.515 3.535 81.685 ;
      RECT 2.905 81.515 3.075 81.685 ;
      RECT 2.445 81.515 2.615 81.685 ;
      RECT 1.985 81.515 2.155 81.685 ;
      RECT 1.525 81.515 1.695 81.685 ;
      RECT 1.065 81.515 1.235 81.685 ;
      RECT 0.605 81.515 0.775 81.685 ;
      RECT 0.145 81.515 0.315 81.685 ;
      RECT 84.325 78.795 84.495 78.965 ;
      RECT 0.145 78.795 0.315 78.965 ;
      RECT 84.325 76.075 84.495 76.245 ;
      RECT 0.145 76.075 0.315 76.245 ;
      RECT 84.325 73.355 84.495 73.525 ;
      RECT 0.145 73.355 0.315 73.525 ;
      RECT 84.325 70.635 84.495 70.805 ;
      RECT 0.145 70.635 0.315 70.805 ;
      RECT 84.325 67.915 84.495 68.085 ;
      RECT 0.145 67.915 0.315 68.085 ;
      RECT 84.325 65.195 84.495 65.365 ;
      RECT 0.145 65.195 0.315 65.365 ;
      RECT 84.325 62.475 84.495 62.645 ;
      RECT 0.145 62.475 0.315 62.645 ;
      RECT 84.325 59.755 84.495 59.925 ;
      RECT 0.145 59.755 0.315 59.925 ;
      RECT 84.325 57.035 84.495 57.205 ;
      RECT 0.145 57.035 0.315 57.205 ;
      RECT 84.325 54.315 84.495 54.485 ;
      RECT 0.145 54.315 0.315 54.485 ;
      RECT 84.325 51.595 84.495 51.765 ;
      RECT 0.145 51.595 0.315 51.765 ;
      RECT 84.325 48.875 84.495 49.045 ;
      RECT 0.145 48.875 0.315 49.045 ;
      RECT 84.325 46.155 84.495 46.325 ;
      RECT 0.145 46.155 0.315 46.325 ;
      RECT 84.325 43.435 84.495 43.605 ;
      RECT 0.145 43.435 0.315 43.605 ;
      RECT 84.325 40.715 84.495 40.885 ;
      RECT 0.145 40.715 0.315 40.885 ;
      RECT 84.325 37.995 84.495 38.165 ;
      RECT 0.145 37.995 0.315 38.165 ;
      RECT 84.325 35.275 84.495 35.445 ;
      RECT 0.145 35.275 0.315 35.445 ;
      RECT 84.325 32.555 84.495 32.725 ;
      RECT 0.145 32.555 0.315 32.725 ;
      RECT 84.325 29.835 84.495 30.005 ;
      RECT 0.145 29.835 0.315 30.005 ;
      RECT 84.325 27.115 84.495 27.285 ;
      RECT 0.145 27.115 0.315 27.285 ;
      RECT 84.325 24.395 84.495 24.565 ;
      RECT 0.145 24.395 0.315 24.565 ;
      RECT 84.325 21.675 84.495 21.845 ;
      RECT 0.145 21.675 0.315 21.845 ;
      RECT 84.325 18.955 84.495 19.125 ;
      RECT 0.145 18.955 0.315 19.125 ;
      RECT 84.325 16.235 84.495 16.405 ;
      RECT 83.865 16.235 84.035 16.405 ;
      RECT 83.405 16.235 83.575 16.405 ;
      RECT 82.945 16.235 83.115 16.405 ;
      RECT 82.485 16.235 82.655 16.405 ;
      RECT 82.025 16.235 82.195 16.405 ;
      RECT 81.565 16.235 81.735 16.405 ;
      RECT 81.105 16.235 81.275 16.405 ;
      RECT 80.645 16.235 80.815 16.405 ;
      RECT 80.185 16.235 80.355 16.405 ;
      RECT 79.725 16.235 79.895 16.405 ;
      RECT 79.265 16.235 79.435 16.405 ;
      RECT 78.805 16.235 78.975 16.405 ;
      RECT 78.345 16.235 78.515 16.405 ;
      RECT 77.885 16.235 78.055 16.405 ;
      RECT 77.425 16.235 77.595 16.405 ;
      RECT 76.965 16.235 77.135 16.405 ;
      RECT 76.505 16.235 76.675 16.405 ;
      RECT 76.045 16.235 76.215 16.405 ;
      RECT 75.585 16.235 75.755 16.405 ;
      RECT 75.125 16.235 75.295 16.405 ;
      RECT 74.665 16.235 74.835 16.405 ;
      RECT 74.205 16.235 74.375 16.405 ;
      RECT 73.745 16.235 73.915 16.405 ;
      RECT 73.285 16.235 73.455 16.405 ;
      RECT 72.825 16.235 72.995 16.405 ;
      RECT 72.365 16.235 72.535 16.405 ;
      RECT 71.905 16.235 72.075 16.405 ;
      RECT 71.445 16.235 71.615 16.405 ;
      RECT 70.985 16.235 71.155 16.405 ;
      RECT 70.525 16.235 70.695 16.405 ;
      RECT 70.065 16.235 70.235 16.405 ;
      RECT 69.605 16.235 69.775 16.405 ;
      RECT 69.145 16.235 69.315 16.405 ;
      RECT 68.685 16.235 68.855 16.405 ;
      RECT 68.225 16.235 68.395 16.405 ;
      RECT 67.765 16.235 67.935 16.405 ;
      RECT 67.305 16.235 67.475 16.405 ;
      RECT 66.845 16.235 67.015 16.405 ;
      RECT 66.385 16.235 66.555 16.405 ;
      RECT 65.925 16.235 66.095 16.405 ;
      RECT 0.145 16.235 0.315 16.405 ;
      RECT 65.925 13.515 66.095 13.685 ;
      RECT 0.145 13.515 0.315 13.685 ;
      RECT 65.925 10.795 66.095 10.965 ;
      RECT 0.145 10.795 0.315 10.965 ;
      RECT 65.925 8.075 66.095 8.245 ;
      RECT 0.145 8.075 0.315 8.245 ;
      RECT 65.925 5.355 66.095 5.525 ;
      RECT 0.145 5.355 0.315 5.525 ;
      RECT 65.925 2.635 66.095 2.805 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 65.925 -0.085 66.095 0.085 ;
      RECT 65.465 -0.085 65.635 0.085 ;
      RECT 65.005 -0.085 65.175 0.085 ;
      RECT 64.545 -0.085 64.715 0.085 ;
      RECT 64.085 -0.085 64.255 0.085 ;
      RECT 63.625 -0.085 63.795 0.085 ;
      RECT 63.165 -0.085 63.335 0.085 ;
      RECT 62.705 -0.085 62.875 0.085 ;
      RECT 62.245 -0.085 62.415 0.085 ;
      RECT 61.785 -0.085 61.955 0.085 ;
      RECT 61.325 -0.085 61.495 0.085 ;
      RECT 60.865 -0.085 61.035 0.085 ;
      RECT 60.405 -0.085 60.575 0.085 ;
      RECT 59.945 -0.085 60.115 0.085 ;
      RECT 59.485 -0.085 59.655 0.085 ;
      RECT 59.025 -0.085 59.195 0.085 ;
      RECT 58.565 -0.085 58.735 0.085 ;
      RECT 58.105 -0.085 58.275 0.085 ;
      RECT 57.645 -0.085 57.815 0.085 ;
      RECT 57.185 -0.085 57.355 0.085 ;
      RECT 56.725 -0.085 56.895 0.085 ;
      RECT 56.265 -0.085 56.435 0.085 ;
      RECT 55.805 -0.085 55.975 0.085 ;
      RECT 55.345 -0.085 55.515 0.085 ;
      RECT 54.885 -0.085 55.055 0.085 ;
      RECT 54.425 -0.085 54.595 0.085 ;
      RECT 53.965 -0.085 54.135 0.085 ;
      RECT 53.505 -0.085 53.675 0.085 ;
      RECT 53.045 -0.085 53.215 0.085 ;
      RECT 52.585 -0.085 52.755 0.085 ;
      RECT 52.125 -0.085 52.295 0.085 ;
      RECT 51.665 -0.085 51.835 0.085 ;
      RECT 51.205 -0.085 51.375 0.085 ;
      RECT 50.745 -0.085 50.915 0.085 ;
      RECT 50.285 -0.085 50.455 0.085 ;
      RECT 49.825 -0.085 49.995 0.085 ;
      RECT 49.365 -0.085 49.535 0.085 ;
      RECT 48.905 -0.085 49.075 0.085 ;
      RECT 48.445 -0.085 48.615 0.085 ;
      RECT 47.985 -0.085 48.155 0.085 ;
      RECT 47.525 -0.085 47.695 0.085 ;
      RECT 47.065 -0.085 47.235 0.085 ;
      RECT 46.605 -0.085 46.775 0.085 ;
      RECT 46.145 -0.085 46.315 0.085 ;
      RECT 45.685 -0.085 45.855 0.085 ;
      RECT 45.225 -0.085 45.395 0.085 ;
      RECT 44.765 -0.085 44.935 0.085 ;
      RECT 44.305 -0.085 44.475 0.085 ;
      RECT 43.845 -0.085 44.015 0.085 ;
      RECT 43.385 -0.085 43.555 0.085 ;
      RECT 42.925 -0.085 43.095 0.085 ;
      RECT 42.465 -0.085 42.635 0.085 ;
      RECT 42.005 -0.085 42.175 0.085 ;
      RECT 41.545 -0.085 41.715 0.085 ;
      RECT 41.085 -0.085 41.255 0.085 ;
      RECT 40.625 -0.085 40.795 0.085 ;
      RECT 40.165 -0.085 40.335 0.085 ;
      RECT 39.705 -0.085 39.875 0.085 ;
      RECT 39.245 -0.085 39.415 0.085 ;
      RECT 38.785 -0.085 38.955 0.085 ;
      RECT 38.325 -0.085 38.495 0.085 ;
      RECT 37.865 -0.085 38.035 0.085 ;
      RECT 37.405 -0.085 37.575 0.085 ;
      RECT 36.945 -0.085 37.115 0.085 ;
      RECT 36.485 -0.085 36.655 0.085 ;
      RECT 36.025 -0.085 36.195 0.085 ;
      RECT 35.565 -0.085 35.735 0.085 ;
      RECT 35.105 -0.085 35.275 0.085 ;
      RECT 34.645 -0.085 34.815 0.085 ;
      RECT 34.185 -0.085 34.355 0.085 ;
      RECT 33.725 -0.085 33.895 0.085 ;
      RECT 33.265 -0.085 33.435 0.085 ;
      RECT 32.805 -0.085 32.975 0.085 ;
      RECT 32.345 -0.085 32.515 0.085 ;
      RECT 31.885 -0.085 32.055 0.085 ;
      RECT 31.425 -0.085 31.595 0.085 ;
      RECT 30.965 -0.085 31.135 0.085 ;
      RECT 30.505 -0.085 30.675 0.085 ;
      RECT 30.045 -0.085 30.215 0.085 ;
      RECT 29.585 -0.085 29.755 0.085 ;
      RECT 29.125 -0.085 29.295 0.085 ;
      RECT 28.665 -0.085 28.835 0.085 ;
      RECT 28.205 -0.085 28.375 0.085 ;
      RECT 27.745 -0.085 27.915 0.085 ;
      RECT 27.285 -0.085 27.455 0.085 ;
      RECT 26.825 -0.085 26.995 0.085 ;
      RECT 26.365 -0.085 26.535 0.085 ;
      RECT 25.905 -0.085 26.075 0.085 ;
      RECT 25.445 -0.085 25.615 0.085 ;
      RECT 24.985 -0.085 25.155 0.085 ;
      RECT 24.525 -0.085 24.695 0.085 ;
      RECT 24.065 -0.085 24.235 0.085 ;
      RECT 23.605 -0.085 23.775 0.085 ;
      RECT 23.145 -0.085 23.315 0.085 ;
      RECT 22.685 -0.085 22.855 0.085 ;
      RECT 22.225 -0.085 22.395 0.085 ;
      RECT 21.765 -0.085 21.935 0.085 ;
      RECT 21.305 -0.085 21.475 0.085 ;
      RECT 20.845 -0.085 21.015 0.085 ;
      RECT 20.385 -0.085 20.555 0.085 ;
      RECT 19.925 -0.085 20.095 0.085 ;
      RECT 19.465 -0.085 19.635 0.085 ;
      RECT 19.005 -0.085 19.175 0.085 ;
      RECT 18.545 -0.085 18.715 0.085 ;
      RECT 18.085 -0.085 18.255 0.085 ;
      RECT 17.625 -0.085 17.795 0.085 ;
      RECT 17.165 -0.085 17.335 0.085 ;
      RECT 16.705 -0.085 16.875 0.085 ;
      RECT 16.245 -0.085 16.415 0.085 ;
      RECT 15.785 -0.085 15.955 0.085 ;
      RECT 15.325 -0.085 15.495 0.085 ;
      RECT 14.865 -0.085 15.035 0.085 ;
      RECT 14.405 -0.085 14.575 0.085 ;
      RECT 13.945 -0.085 14.115 0.085 ;
      RECT 13.485 -0.085 13.655 0.085 ;
      RECT 13.025 -0.085 13.195 0.085 ;
      RECT 12.565 -0.085 12.735 0.085 ;
      RECT 12.105 -0.085 12.275 0.085 ;
      RECT 11.645 -0.085 11.815 0.085 ;
      RECT 11.185 -0.085 11.355 0.085 ;
      RECT 10.725 -0.085 10.895 0.085 ;
      RECT 10.265 -0.085 10.435 0.085 ;
      RECT 9.805 -0.085 9.975 0.085 ;
      RECT 9.345 -0.085 9.515 0.085 ;
      RECT 8.885 -0.085 9.055 0.085 ;
      RECT 8.425 -0.085 8.595 0.085 ;
      RECT 7.965 -0.085 8.135 0.085 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.145 -0.085 0.315 0.085 ;
    LAYER via ;
      RECT 18.325 1.625 18.475 1.775 ;
    LAYER via2 ;
      RECT 82.7 71.98 82.9 72.18 ;
      RECT 83.16 59.74 83.36 59.94 ;
      RECT 82.7 54.3 82.9 54.5 ;
      RECT 83.16 51.58 83.36 51.78 ;
      RECT 82.7 48.86 82.9 49.06 ;
      RECT 83.16 29.82 83.36 30.02 ;
      RECT 82.7 28.46 82.9 28.66 ;
      RECT 83.16 24.38 83.36 24.58 ;
    LAYER fieldpoly ;
      POLYGON 84.5 81.46 84.5 16.46 66.1 16.46 66.1 0.14 0.14 0.14 0.14 81.46 ;
    LAYER diff ;
      POLYGON 84.64 81.6 84.64 16.32 66.24 16.32 66.24 0 0 0 0 81.6 ;
    LAYER nwell ;
      RECT 83.99 77.465 84.83 80.295 ;
      RECT -0.19 77.465 3.87 80.295 ;
      RECT 83.53 72.025 84.83 74.855 ;
      RECT -0.19 72.025 3.87 74.855 ;
      POLYGON 84.83 69.415 84.83 66.585 83.99 66.585 83.99 67.81 83.53 67.81 83.53 69.415 ;
      RECT -0.19 66.585 3.87 69.415 ;
      RECT 80.77 61.145 84.83 63.975 ;
      RECT -0.19 61.145 3.87 63.975 ;
      RECT 83.53 55.705 84.83 58.535 ;
      RECT -0.19 55.705 3.87 58.535 ;
      RECT 83.53 50.265 84.83 53.095 ;
      RECT -0.19 50.265 3.87 53.095 ;
      RECT 83.53 44.825 84.83 47.655 ;
      RECT -0.19 44.825 3.87 47.655 ;
      RECT 83.53 39.385 84.83 42.215 ;
      RECT -0.19 39.385 3.87 42.215 ;
      RECT 83.53 33.945 84.83 36.775 ;
      RECT -0.19 33.945 3.87 36.775 ;
      RECT 83.53 28.505 84.83 31.335 ;
      RECT -0.19 28.505 3.87 31.335 ;
      RECT 83.53 23.065 84.83 25.895 ;
      RECT -0.19 23.065 3.87 25.895 ;
      POLYGON 84.83 20.455 84.83 17.625 83.99 17.625 83.99 18.85 83.53 18.85 83.53 20.455 ;
      RECT -0.19 17.625 3.87 20.455 ;
      RECT 65.59 12.185 66.43 15.015 ;
      RECT -0.19 12.185 3.87 15.015 ;
      RECT 65.13 6.745 66.43 9.575 ;
      POLYGON 3.87 9.575 3.87 7.97 2.03 7.97 2.03 6.745 -0.19 6.745 -0.19 9.575 ;
      POLYGON 66.43 4.135 66.43 1.305 65.59 1.305 65.59 2.53 62.37 2.53 62.37 4.135 ;
      RECT -0.19 1.305 3.87 4.135 ;
      POLYGON 84.64 81.6 84.64 16.32 66.24 16.32 66.24 0 0 0 0 81.6 ;
    LAYER pwell ;
      RECT 77.87 81.55 78.09 81.72 ;
      RECT 74.19 81.55 74.41 81.72 ;
      RECT 70.51 81.55 70.73 81.72 ;
      RECT 66.83 81.55 67.05 81.72 ;
      RECT 62.23 81.55 62.45 81.72 ;
      RECT 58.55 81.55 58.77 81.72 ;
      RECT 54.87 81.55 55.09 81.72 ;
      RECT 51.19 81.55 51.41 81.72 ;
      RECT 47.51 81.55 47.73 81.72 ;
      RECT 43.83 81.55 44.05 81.72 ;
      RECT 40.15 81.55 40.37 81.72 ;
      RECT 36.47 81.55 36.69 81.72 ;
      RECT 32.79 81.55 33.01 81.72 ;
      RECT 29.11 81.55 29.33 81.72 ;
      RECT 25.43 81.55 25.65 81.72 ;
      RECT 21.75 81.55 21.97 81.72 ;
      RECT 18.07 81.55 18.29 81.72 ;
      RECT 11.17 81.55 11.39 81.72 ;
      RECT 7.49 81.55 7.71 81.72 ;
      RECT 3.81 81.55 4.03 81.72 ;
      RECT 0.13 81.55 0.35 81.72 ;
      RECT 81.595 81.54 81.705 81.66 ;
      RECT 14.895 81.54 15.005 81.66 ;
      RECT 84.32 81.545 84.44 81.655 ;
      RECT 16.7 81.545 16.82 81.655 ;
      RECT 83.415 81.54 83.575 81.65 ;
      RECT 83.415 16.27 83.575 16.38 ;
      RECT 81.595 16.26 81.705 16.38 ;
      RECT 84.32 16.265 84.44 16.375 ;
      RECT 77.87 16.2 78.09 16.37 ;
      RECT 74.19 16.2 74.41 16.37 ;
      RECT 70.51 16.2 70.73 16.37 ;
      RECT 66.83 16.2 67.05 16.37 ;
      RECT 14.895 -0.06 15.005 0.06 ;
      RECT 65.92 -0.055 66.04 0.055 ;
      RECT 16.7 -0.055 16.82 0.055 ;
      RECT 62.23 -0.12 62.45 0.05 ;
      RECT 58.55 -0.12 58.77 0.05 ;
      RECT 54.87 -0.12 55.09 0.05 ;
      RECT 51.19 -0.12 51.41 0.05 ;
      RECT 47.51 -0.12 47.73 0.05 ;
      RECT 43.83 -0.12 44.05 0.05 ;
      RECT 40.15 -0.12 40.37 0.05 ;
      RECT 36.47 -0.12 36.69 0.05 ;
      RECT 32.79 -0.12 33.01 0.05 ;
      RECT 29.11 -0.12 29.33 0.05 ;
      RECT 25.43 -0.12 25.65 0.05 ;
      RECT 21.75 -0.12 21.97 0.05 ;
      RECT 18.07 -0.12 18.29 0.05 ;
      RECT 11.17 -0.12 11.39 0.05 ;
      RECT 7.49 -0.12 7.71 0.05 ;
      RECT 3.81 -0.12 4.03 0.05 ;
      RECT 0.13 -0.12 0.35 0.05 ;
      POLYGON 84.64 81.6 84.64 16.32 66.24 16.32 66.24 0 0 0 0 81.6 ;
    LAYER OVERLAP ;
      POLYGON 0 0 0 81.6 84.64 81.6 84.64 16.32 66.24 16.32 66.24 0 ;
  END
END sb_0__2_

END LIBRARY
