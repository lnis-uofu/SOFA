//
//
//
//
//
//
//
//
`timescale 1ns / 1ps

//
module fpga_core(prog_clk,
                Test_en,
                clk,
                gfpga_pad_GPIO_A,
                gfpga_pad_GPIO_IE,
                gfpga_pad_GPIO_OE,
                gfpga_pad_GPIO_Y,
                ccff_head,
                ccff_tail);
//
input [0:0] prog_clk;
//
input [0:0] Test_en;
//
input [0:0] clk;
//
output [0:47] gfpga_pad_GPIO_A;
//
output [0:47] gfpga_pad_GPIO_IE;
//
output [0:47] gfpga_pad_GPIO_OE;
//
inout [0:47] gfpga_pad_GPIO_Y;
//
input [0:0] ccff_head;
//
output [0:0] ccff_tail;

//
//


//
//


wire [0:0] cbx_1__0__0_bottom_grid_pin_0_;
wire [0:0] cbx_1__0__0_ccff_tail;
wire [0:19] cbx_1__0__0_chanx_left_out;
wire [0:19] cbx_1__0__0_chanx_right_out;
wire [0:0] cbx_1__0__0_top_grid_pin_16_;
wire [0:0] cbx_1__0__0_top_grid_pin_17_;
wire [0:0] cbx_1__0__0_top_grid_pin_18_;
wire [0:0] cbx_1__0__0_top_grid_pin_19_;
wire [0:0] cbx_1__0__0_top_grid_pin_20_;
wire [0:0] cbx_1__0__0_top_grid_pin_21_;
wire [0:0] cbx_1__0__0_top_grid_pin_22_;
wire [0:0] cbx_1__0__0_top_grid_pin_23_;
wire [0:0] cbx_1__0__0_top_grid_pin_24_;
wire [0:0] cbx_1__0__0_top_grid_pin_25_;
wire [0:0] cbx_1__0__0_top_grid_pin_26_;
wire [0:0] cbx_1__0__0_top_grid_pin_27_;
wire [0:0] cbx_1__0__0_top_grid_pin_28_;
wire [0:0] cbx_1__0__0_top_grid_pin_29_;
wire [0:0] cbx_1__0__0_top_grid_pin_30_;
wire [0:0] cbx_1__0__0_top_grid_pin_31_;
wire [0:0] cbx_1__0__10_bottom_grid_pin_0_;
wire [0:0] cbx_1__0__10_ccff_tail;
wire [0:19] cbx_1__0__10_chanx_left_out;
wire [0:19] cbx_1__0__10_chanx_right_out;
wire [0:0] cbx_1__0__10_top_grid_pin_16_;
wire [0:0] cbx_1__0__10_top_grid_pin_17_;
wire [0:0] cbx_1__0__10_top_grid_pin_18_;
wire [0:0] cbx_1__0__10_top_grid_pin_19_;
wire [0:0] cbx_1__0__10_top_grid_pin_20_;
wire [0:0] cbx_1__0__10_top_grid_pin_21_;
wire [0:0] cbx_1__0__10_top_grid_pin_22_;
wire [0:0] cbx_1__0__10_top_grid_pin_23_;
wire [0:0] cbx_1__0__10_top_grid_pin_24_;
wire [0:0] cbx_1__0__10_top_grid_pin_25_;
wire [0:0] cbx_1__0__10_top_grid_pin_26_;
wire [0:0] cbx_1__0__10_top_grid_pin_27_;
wire [0:0] cbx_1__0__10_top_grid_pin_28_;
wire [0:0] cbx_1__0__10_top_grid_pin_29_;
wire [0:0] cbx_1__0__10_top_grid_pin_30_;
wire [0:0] cbx_1__0__10_top_grid_pin_31_;
wire [0:0] cbx_1__0__11_bottom_grid_pin_0_;
wire [0:0] cbx_1__0__11_ccff_tail;
wire [0:19] cbx_1__0__11_chanx_left_out;
wire [0:19] cbx_1__0__11_chanx_right_out;
wire [0:0] cbx_1__0__11_top_grid_pin_16_;
wire [0:0] cbx_1__0__11_top_grid_pin_17_;
wire [0:0] cbx_1__0__11_top_grid_pin_18_;
wire [0:0] cbx_1__0__11_top_grid_pin_19_;
wire [0:0] cbx_1__0__11_top_grid_pin_20_;
wire [0:0] cbx_1__0__11_top_grid_pin_21_;
wire [0:0] cbx_1__0__11_top_grid_pin_22_;
wire [0:0] cbx_1__0__11_top_grid_pin_23_;
wire [0:0] cbx_1__0__11_top_grid_pin_24_;
wire [0:0] cbx_1__0__11_top_grid_pin_25_;
wire [0:0] cbx_1__0__11_top_grid_pin_26_;
wire [0:0] cbx_1__0__11_top_grid_pin_27_;
wire [0:0] cbx_1__0__11_top_grid_pin_28_;
wire [0:0] cbx_1__0__11_top_grid_pin_29_;
wire [0:0] cbx_1__0__11_top_grid_pin_30_;
wire [0:0] cbx_1__0__11_top_grid_pin_31_;
wire [0:0] cbx_1__0__1_bottom_grid_pin_0_;
wire [0:0] cbx_1__0__1_ccff_tail;
wire [0:19] cbx_1__0__1_chanx_left_out;
wire [0:19] cbx_1__0__1_chanx_right_out;
wire [0:0] cbx_1__0__1_top_grid_pin_16_;
wire [0:0] cbx_1__0__1_top_grid_pin_17_;
wire [0:0] cbx_1__0__1_top_grid_pin_18_;
wire [0:0] cbx_1__0__1_top_grid_pin_19_;
wire [0:0] cbx_1__0__1_top_grid_pin_20_;
wire [0:0] cbx_1__0__1_top_grid_pin_21_;
wire [0:0] cbx_1__0__1_top_grid_pin_22_;
wire [0:0] cbx_1__0__1_top_grid_pin_23_;
wire [0:0] cbx_1__0__1_top_grid_pin_24_;
wire [0:0] cbx_1__0__1_top_grid_pin_25_;
wire [0:0] cbx_1__0__1_top_grid_pin_26_;
wire [0:0] cbx_1__0__1_top_grid_pin_27_;
wire [0:0] cbx_1__0__1_top_grid_pin_28_;
wire [0:0] cbx_1__0__1_top_grid_pin_29_;
wire [0:0] cbx_1__0__1_top_grid_pin_30_;
wire [0:0] cbx_1__0__1_top_grid_pin_31_;
wire [0:0] cbx_1__0__2_bottom_grid_pin_0_;
wire [0:0] cbx_1__0__2_ccff_tail;
wire [0:19] cbx_1__0__2_chanx_left_out;
wire [0:19] cbx_1__0__2_chanx_right_out;
wire [0:0] cbx_1__0__2_top_grid_pin_16_;
wire [0:0] cbx_1__0__2_top_grid_pin_17_;
wire [0:0] cbx_1__0__2_top_grid_pin_18_;
wire [0:0] cbx_1__0__2_top_grid_pin_19_;
wire [0:0] cbx_1__0__2_top_grid_pin_20_;
wire [0:0] cbx_1__0__2_top_grid_pin_21_;
wire [0:0] cbx_1__0__2_top_grid_pin_22_;
wire [0:0] cbx_1__0__2_top_grid_pin_23_;
wire [0:0] cbx_1__0__2_top_grid_pin_24_;
wire [0:0] cbx_1__0__2_top_grid_pin_25_;
wire [0:0] cbx_1__0__2_top_grid_pin_26_;
wire [0:0] cbx_1__0__2_top_grid_pin_27_;
wire [0:0] cbx_1__0__2_top_grid_pin_28_;
wire [0:0] cbx_1__0__2_top_grid_pin_29_;
wire [0:0] cbx_1__0__2_top_grid_pin_30_;
wire [0:0] cbx_1__0__2_top_grid_pin_31_;
wire [0:0] cbx_1__0__3_bottom_grid_pin_0_;
wire [0:0] cbx_1__0__3_ccff_tail;
wire [0:19] cbx_1__0__3_chanx_left_out;
wire [0:19] cbx_1__0__3_chanx_right_out;
wire [0:0] cbx_1__0__3_top_grid_pin_16_;
wire [0:0] cbx_1__0__3_top_grid_pin_17_;
wire [0:0] cbx_1__0__3_top_grid_pin_18_;
wire [0:0] cbx_1__0__3_top_grid_pin_19_;
wire [0:0] cbx_1__0__3_top_grid_pin_20_;
wire [0:0] cbx_1__0__3_top_grid_pin_21_;
wire [0:0] cbx_1__0__3_top_grid_pin_22_;
wire [0:0] cbx_1__0__3_top_grid_pin_23_;
wire [0:0] cbx_1__0__3_top_grid_pin_24_;
wire [0:0] cbx_1__0__3_top_grid_pin_25_;
wire [0:0] cbx_1__0__3_top_grid_pin_26_;
wire [0:0] cbx_1__0__3_top_grid_pin_27_;
wire [0:0] cbx_1__0__3_top_grid_pin_28_;
wire [0:0] cbx_1__0__3_top_grid_pin_29_;
wire [0:0] cbx_1__0__3_top_grid_pin_30_;
wire [0:0] cbx_1__0__3_top_grid_pin_31_;
wire [0:0] cbx_1__0__4_bottom_grid_pin_0_;
wire [0:0] cbx_1__0__4_ccff_tail;
wire [0:19] cbx_1__0__4_chanx_left_out;
wire [0:19] cbx_1__0__4_chanx_right_out;
wire [0:0] cbx_1__0__4_top_grid_pin_16_;
wire [0:0] cbx_1__0__4_top_grid_pin_17_;
wire [0:0] cbx_1__0__4_top_grid_pin_18_;
wire [0:0] cbx_1__0__4_top_grid_pin_19_;
wire [0:0] cbx_1__0__4_top_grid_pin_20_;
wire [0:0] cbx_1__0__4_top_grid_pin_21_;
wire [0:0] cbx_1__0__4_top_grid_pin_22_;
wire [0:0] cbx_1__0__4_top_grid_pin_23_;
wire [0:0] cbx_1__0__4_top_grid_pin_24_;
wire [0:0] cbx_1__0__4_top_grid_pin_25_;
wire [0:0] cbx_1__0__4_top_grid_pin_26_;
wire [0:0] cbx_1__0__4_top_grid_pin_27_;
wire [0:0] cbx_1__0__4_top_grid_pin_28_;
wire [0:0] cbx_1__0__4_top_grid_pin_29_;
wire [0:0] cbx_1__0__4_top_grid_pin_30_;
wire [0:0] cbx_1__0__4_top_grid_pin_31_;
wire [0:0] cbx_1__0__5_bottom_grid_pin_0_;
wire [0:0] cbx_1__0__5_ccff_tail;
wire [0:19] cbx_1__0__5_chanx_left_out;
wire [0:19] cbx_1__0__5_chanx_right_out;
wire [0:0] cbx_1__0__5_top_grid_pin_16_;
wire [0:0] cbx_1__0__5_top_grid_pin_17_;
wire [0:0] cbx_1__0__5_top_grid_pin_18_;
wire [0:0] cbx_1__0__5_top_grid_pin_19_;
wire [0:0] cbx_1__0__5_top_grid_pin_20_;
wire [0:0] cbx_1__0__5_top_grid_pin_21_;
wire [0:0] cbx_1__0__5_top_grid_pin_22_;
wire [0:0] cbx_1__0__5_top_grid_pin_23_;
wire [0:0] cbx_1__0__5_top_grid_pin_24_;
wire [0:0] cbx_1__0__5_top_grid_pin_25_;
wire [0:0] cbx_1__0__5_top_grid_pin_26_;
wire [0:0] cbx_1__0__5_top_grid_pin_27_;
wire [0:0] cbx_1__0__5_top_grid_pin_28_;
wire [0:0] cbx_1__0__5_top_grid_pin_29_;
wire [0:0] cbx_1__0__5_top_grid_pin_30_;
wire [0:0] cbx_1__0__5_top_grid_pin_31_;
wire [0:0] cbx_1__0__6_bottom_grid_pin_0_;
wire [0:0] cbx_1__0__6_ccff_tail;
wire [0:19] cbx_1__0__6_chanx_left_out;
wire [0:19] cbx_1__0__6_chanx_right_out;
wire [0:0] cbx_1__0__6_top_grid_pin_16_;
wire [0:0] cbx_1__0__6_top_grid_pin_17_;
wire [0:0] cbx_1__0__6_top_grid_pin_18_;
wire [0:0] cbx_1__0__6_top_grid_pin_19_;
wire [0:0] cbx_1__0__6_top_grid_pin_20_;
wire [0:0] cbx_1__0__6_top_grid_pin_21_;
wire [0:0] cbx_1__0__6_top_grid_pin_22_;
wire [0:0] cbx_1__0__6_top_grid_pin_23_;
wire [0:0] cbx_1__0__6_top_grid_pin_24_;
wire [0:0] cbx_1__0__6_top_grid_pin_25_;
wire [0:0] cbx_1__0__6_top_grid_pin_26_;
wire [0:0] cbx_1__0__6_top_grid_pin_27_;
wire [0:0] cbx_1__0__6_top_grid_pin_28_;
wire [0:0] cbx_1__0__6_top_grid_pin_29_;
wire [0:0] cbx_1__0__6_top_grid_pin_30_;
wire [0:0] cbx_1__0__6_top_grid_pin_31_;
wire [0:0] cbx_1__0__7_bottom_grid_pin_0_;
wire [0:0] cbx_1__0__7_ccff_tail;
wire [0:19] cbx_1__0__7_chanx_left_out;
wire [0:19] cbx_1__0__7_chanx_right_out;
wire [0:0] cbx_1__0__7_top_grid_pin_16_;
wire [0:0] cbx_1__0__7_top_grid_pin_17_;
wire [0:0] cbx_1__0__7_top_grid_pin_18_;
wire [0:0] cbx_1__0__7_top_grid_pin_19_;
wire [0:0] cbx_1__0__7_top_grid_pin_20_;
wire [0:0] cbx_1__0__7_top_grid_pin_21_;
wire [0:0] cbx_1__0__7_top_grid_pin_22_;
wire [0:0] cbx_1__0__7_top_grid_pin_23_;
wire [0:0] cbx_1__0__7_top_grid_pin_24_;
wire [0:0] cbx_1__0__7_top_grid_pin_25_;
wire [0:0] cbx_1__0__7_top_grid_pin_26_;
wire [0:0] cbx_1__0__7_top_grid_pin_27_;
wire [0:0] cbx_1__0__7_top_grid_pin_28_;
wire [0:0] cbx_1__0__7_top_grid_pin_29_;
wire [0:0] cbx_1__0__7_top_grid_pin_30_;
wire [0:0] cbx_1__0__7_top_grid_pin_31_;
wire [0:0] cbx_1__0__8_bottom_grid_pin_0_;
wire [0:0] cbx_1__0__8_ccff_tail;
wire [0:19] cbx_1__0__8_chanx_left_out;
wire [0:19] cbx_1__0__8_chanx_right_out;
wire [0:0] cbx_1__0__8_top_grid_pin_16_;
wire [0:0] cbx_1__0__8_top_grid_pin_17_;
wire [0:0] cbx_1__0__8_top_grid_pin_18_;
wire [0:0] cbx_1__0__8_top_grid_pin_19_;
wire [0:0] cbx_1__0__8_top_grid_pin_20_;
wire [0:0] cbx_1__0__8_top_grid_pin_21_;
wire [0:0] cbx_1__0__8_top_grid_pin_22_;
wire [0:0] cbx_1__0__8_top_grid_pin_23_;
wire [0:0] cbx_1__0__8_top_grid_pin_24_;
wire [0:0] cbx_1__0__8_top_grid_pin_25_;
wire [0:0] cbx_1__0__8_top_grid_pin_26_;
wire [0:0] cbx_1__0__8_top_grid_pin_27_;
wire [0:0] cbx_1__0__8_top_grid_pin_28_;
wire [0:0] cbx_1__0__8_top_grid_pin_29_;
wire [0:0] cbx_1__0__8_top_grid_pin_30_;
wire [0:0] cbx_1__0__8_top_grid_pin_31_;
wire [0:0] cbx_1__0__9_bottom_grid_pin_0_;
wire [0:0] cbx_1__0__9_ccff_tail;
wire [0:19] cbx_1__0__9_chanx_left_out;
wire [0:19] cbx_1__0__9_chanx_right_out;
wire [0:0] cbx_1__0__9_top_grid_pin_16_;
wire [0:0] cbx_1__0__9_top_grid_pin_17_;
wire [0:0] cbx_1__0__9_top_grid_pin_18_;
wire [0:0] cbx_1__0__9_top_grid_pin_19_;
wire [0:0] cbx_1__0__9_top_grid_pin_20_;
wire [0:0] cbx_1__0__9_top_grid_pin_21_;
wire [0:0] cbx_1__0__9_top_grid_pin_22_;
wire [0:0] cbx_1__0__9_top_grid_pin_23_;
wire [0:0] cbx_1__0__9_top_grid_pin_24_;
wire [0:0] cbx_1__0__9_top_grid_pin_25_;
wire [0:0] cbx_1__0__9_top_grid_pin_26_;
wire [0:0] cbx_1__0__9_top_grid_pin_27_;
wire [0:0] cbx_1__0__9_top_grid_pin_28_;
wire [0:0] cbx_1__0__9_top_grid_pin_29_;
wire [0:0] cbx_1__0__9_top_grid_pin_30_;
wire [0:0] cbx_1__0__9_top_grid_pin_31_;
wire [0:0] cbx_1__12__0_ccff_tail;
wire [0:19] cbx_1__12__0_chanx_left_out;
wire [0:19] cbx_1__12__0_chanx_right_out;
wire [0:0] cbx_1__12__0_top_grid_pin_0_;
wire [0:0] cbx_1__12__10_ccff_tail;
wire [0:19] cbx_1__12__10_chanx_left_out;
wire [0:19] cbx_1__12__10_chanx_right_out;
wire [0:0] cbx_1__12__10_top_grid_pin_0_;
wire [0:0] cbx_1__12__11_ccff_tail;
wire [0:19] cbx_1__12__11_chanx_left_out;
wire [0:19] cbx_1__12__11_chanx_right_out;
wire [0:0] cbx_1__12__11_top_grid_pin_0_;
wire [0:0] cbx_1__12__1_ccff_tail;
wire [0:19] cbx_1__12__1_chanx_left_out;
wire [0:19] cbx_1__12__1_chanx_right_out;
wire [0:0] cbx_1__12__1_top_grid_pin_0_;
wire [0:0] cbx_1__12__2_ccff_tail;
wire [0:19] cbx_1__12__2_chanx_left_out;
wire [0:19] cbx_1__12__2_chanx_right_out;
wire [0:0] cbx_1__12__2_top_grid_pin_0_;
wire [0:0] cbx_1__12__3_ccff_tail;
wire [0:19] cbx_1__12__3_chanx_left_out;
wire [0:19] cbx_1__12__3_chanx_right_out;
wire [0:0] cbx_1__12__3_top_grid_pin_0_;
wire [0:0] cbx_1__12__4_ccff_tail;
wire [0:19] cbx_1__12__4_chanx_left_out;
wire [0:19] cbx_1__12__4_chanx_right_out;
wire [0:0] cbx_1__12__4_top_grid_pin_0_;
wire [0:0] cbx_1__12__5_ccff_tail;
wire [0:19] cbx_1__12__5_chanx_left_out;
wire [0:19] cbx_1__12__5_chanx_right_out;
wire [0:0] cbx_1__12__5_top_grid_pin_0_;
wire [0:0] cbx_1__12__6_ccff_tail;
wire [0:19] cbx_1__12__6_chanx_left_out;
wire [0:19] cbx_1__12__6_chanx_right_out;
wire [0:0] cbx_1__12__6_top_grid_pin_0_;
wire [0:0] cbx_1__12__7_ccff_tail;
wire [0:19] cbx_1__12__7_chanx_left_out;
wire [0:19] cbx_1__12__7_chanx_right_out;
wire [0:0] cbx_1__12__7_top_grid_pin_0_;
wire [0:0] cbx_1__12__8_ccff_tail;
wire [0:19] cbx_1__12__8_chanx_left_out;
wire [0:19] cbx_1__12__8_chanx_right_out;
wire [0:0] cbx_1__12__8_top_grid_pin_0_;
wire [0:0] cbx_1__12__9_ccff_tail;
wire [0:19] cbx_1__12__9_chanx_left_out;
wire [0:19] cbx_1__12__9_chanx_right_out;
wire [0:0] cbx_1__12__9_top_grid_pin_0_;
wire [0:0] cbx_1__1__0_ccff_tail;
wire [0:19] cbx_1__1__0_chanx_left_out;
wire [0:19] cbx_1__1__0_chanx_right_out;
wire [0:0] cbx_1__1__0_top_grid_pin_16_;
wire [0:0] cbx_1__1__0_top_grid_pin_17_;
wire [0:0] cbx_1__1__0_top_grid_pin_18_;
wire [0:0] cbx_1__1__0_top_grid_pin_19_;
wire [0:0] cbx_1__1__0_top_grid_pin_20_;
wire [0:0] cbx_1__1__0_top_grid_pin_21_;
wire [0:0] cbx_1__1__0_top_grid_pin_22_;
wire [0:0] cbx_1__1__0_top_grid_pin_23_;
wire [0:0] cbx_1__1__0_top_grid_pin_24_;
wire [0:0] cbx_1__1__0_top_grid_pin_25_;
wire [0:0] cbx_1__1__0_top_grid_pin_26_;
wire [0:0] cbx_1__1__0_top_grid_pin_27_;
wire [0:0] cbx_1__1__0_top_grid_pin_28_;
wire [0:0] cbx_1__1__0_top_grid_pin_29_;
wire [0:0] cbx_1__1__0_top_grid_pin_30_;
wire [0:0] cbx_1__1__0_top_grid_pin_31_;
wire [0:0] cbx_1__1__100_ccff_tail;
wire [0:19] cbx_1__1__100_chanx_left_out;
wire [0:19] cbx_1__1__100_chanx_right_out;
wire [0:0] cbx_1__1__100_top_grid_pin_16_;
wire [0:0] cbx_1__1__100_top_grid_pin_17_;
wire [0:0] cbx_1__1__100_top_grid_pin_18_;
wire [0:0] cbx_1__1__100_top_grid_pin_19_;
wire [0:0] cbx_1__1__100_top_grid_pin_20_;
wire [0:0] cbx_1__1__100_top_grid_pin_21_;
wire [0:0] cbx_1__1__100_top_grid_pin_22_;
wire [0:0] cbx_1__1__100_top_grid_pin_23_;
wire [0:0] cbx_1__1__100_top_grid_pin_24_;
wire [0:0] cbx_1__1__100_top_grid_pin_25_;
wire [0:0] cbx_1__1__100_top_grid_pin_26_;
wire [0:0] cbx_1__1__100_top_grid_pin_27_;
wire [0:0] cbx_1__1__100_top_grid_pin_28_;
wire [0:0] cbx_1__1__100_top_grid_pin_29_;
wire [0:0] cbx_1__1__100_top_grid_pin_30_;
wire [0:0] cbx_1__1__100_top_grid_pin_31_;
wire [0:0] cbx_1__1__101_ccff_tail;
wire [0:19] cbx_1__1__101_chanx_left_out;
wire [0:19] cbx_1__1__101_chanx_right_out;
wire [0:0] cbx_1__1__101_top_grid_pin_16_;
wire [0:0] cbx_1__1__101_top_grid_pin_17_;
wire [0:0] cbx_1__1__101_top_grid_pin_18_;
wire [0:0] cbx_1__1__101_top_grid_pin_19_;
wire [0:0] cbx_1__1__101_top_grid_pin_20_;
wire [0:0] cbx_1__1__101_top_grid_pin_21_;
wire [0:0] cbx_1__1__101_top_grid_pin_22_;
wire [0:0] cbx_1__1__101_top_grid_pin_23_;
wire [0:0] cbx_1__1__101_top_grid_pin_24_;
wire [0:0] cbx_1__1__101_top_grid_pin_25_;
wire [0:0] cbx_1__1__101_top_grid_pin_26_;
wire [0:0] cbx_1__1__101_top_grid_pin_27_;
wire [0:0] cbx_1__1__101_top_grid_pin_28_;
wire [0:0] cbx_1__1__101_top_grid_pin_29_;
wire [0:0] cbx_1__1__101_top_grid_pin_30_;
wire [0:0] cbx_1__1__101_top_grid_pin_31_;
wire [0:0] cbx_1__1__102_ccff_tail;
wire [0:19] cbx_1__1__102_chanx_left_out;
wire [0:19] cbx_1__1__102_chanx_right_out;
wire [0:0] cbx_1__1__102_top_grid_pin_16_;
wire [0:0] cbx_1__1__102_top_grid_pin_17_;
wire [0:0] cbx_1__1__102_top_grid_pin_18_;
wire [0:0] cbx_1__1__102_top_grid_pin_19_;
wire [0:0] cbx_1__1__102_top_grid_pin_20_;
wire [0:0] cbx_1__1__102_top_grid_pin_21_;
wire [0:0] cbx_1__1__102_top_grid_pin_22_;
wire [0:0] cbx_1__1__102_top_grid_pin_23_;
wire [0:0] cbx_1__1__102_top_grid_pin_24_;
wire [0:0] cbx_1__1__102_top_grid_pin_25_;
wire [0:0] cbx_1__1__102_top_grid_pin_26_;
wire [0:0] cbx_1__1__102_top_grid_pin_27_;
wire [0:0] cbx_1__1__102_top_grid_pin_28_;
wire [0:0] cbx_1__1__102_top_grid_pin_29_;
wire [0:0] cbx_1__1__102_top_grid_pin_30_;
wire [0:0] cbx_1__1__102_top_grid_pin_31_;
wire [0:0] cbx_1__1__103_ccff_tail;
wire [0:19] cbx_1__1__103_chanx_left_out;
wire [0:19] cbx_1__1__103_chanx_right_out;
wire [0:0] cbx_1__1__103_top_grid_pin_16_;
wire [0:0] cbx_1__1__103_top_grid_pin_17_;
wire [0:0] cbx_1__1__103_top_grid_pin_18_;
wire [0:0] cbx_1__1__103_top_grid_pin_19_;
wire [0:0] cbx_1__1__103_top_grid_pin_20_;
wire [0:0] cbx_1__1__103_top_grid_pin_21_;
wire [0:0] cbx_1__1__103_top_grid_pin_22_;
wire [0:0] cbx_1__1__103_top_grid_pin_23_;
wire [0:0] cbx_1__1__103_top_grid_pin_24_;
wire [0:0] cbx_1__1__103_top_grid_pin_25_;
wire [0:0] cbx_1__1__103_top_grid_pin_26_;
wire [0:0] cbx_1__1__103_top_grid_pin_27_;
wire [0:0] cbx_1__1__103_top_grid_pin_28_;
wire [0:0] cbx_1__1__103_top_grid_pin_29_;
wire [0:0] cbx_1__1__103_top_grid_pin_30_;
wire [0:0] cbx_1__1__103_top_grid_pin_31_;
wire [0:0] cbx_1__1__104_ccff_tail;
wire [0:19] cbx_1__1__104_chanx_left_out;
wire [0:19] cbx_1__1__104_chanx_right_out;
wire [0:0] cbx_1__1__104_top_grid_pin_16_;
wire [0:0] cbx_1__1__104_top_grid_pin_17_;
wire [0:0] cbx_1__1__104_top_grid_pin_18_;
wire [0:0] cbx_1__1__104_top_grid_pin_19_;
wire [0:0] cbx_1__1__104_top_grid_pin_20_;
wire [0:0] cbx_1__1__104_top_grid_pin_21_;
wire [0:0] cbx_1__1__104_top_grid_pin_22_;
wire [0:0] cbx_1__1__104_top_grid_pin_23_;
wire [0:0] cbx_1__1__104_top_grid_pin_24_;
wire [0:0] cbx_1__1__104_top_grid_pin_25_;
wire [0:0] cbx_1__1__104_top_grid_pin_26_;
wire [0:0] cbx_1__1__104_top_grid_pin_27_;
wire [0:0] cbx_1__1__104_top_grid_pin_28_;
wire [0:0] cbx_1__1__104_top_grid_pin_29_;
wire [0:0] cbx_1__1__104_top_grid_pin_30_;
wire [0:0] cbx_1__1__104_top_grid_pin_31_;
wire [0:0] cbx_1__1__105_ccff_tail;
wire [0:19] cbx_1__1__105_chanx_left_out;
wire [0:19] cbx_1__1__105_chanx_right_out;
wire [0:0] cbx_1__1__105_top_grid_pin_16_;
wire [0:0] cbx_1__1__105_top_grid_pin_17_;
wire [0:0] cbx_1__1__105_top_grid_pin_18_;
wire [0:0] cbx_1__1__105_top_grid_pin_19_;
wire [0:0] cbx_1__1__105_top_grid_pin_20_;
wire [0:0] cbx_1__1__105_top_grid_pin_21_;
wire [0:0] cbx_1__1__105_top_grid_pin_22_;
wire [0:0] cbx_1__1__105_top_grid_pin_23_;
wire [0:0] cbx_1__1__105_top_grid_pin_24_;
wire [0:0] cbx_1__1__105_top_grid_pin_25_;
wire [0:0] cbx_1__1__105_top_grid_pin_26_;
wire [0:0] cbx_1__1__105_top_grid_pin_27_;
wire [0:0] cbx_1__1__105_top_grid_pin_28_;
wire [0:0] cbx_1__1__105_top_grid_pin_29_;
wire [0:0] cbx_1__1__105_top_grid_pin_30_;
wire [0:0] cbx_1__1__105_top_grid_pin_31_;
wire [0:0] cbx_1__1__106_ccff_tail;
wire [0:19] cbx_1__1__106_chanx_left_out;
wire [0:19] cbx_1__1__106_chanx_right_out;
wire [0:0] cbx_1__1__106_top_grid_pin_16_;
wire [0:0] cbx_1__1__106_top_grid_pin_17_;
wire [0:0] cbx_1__1__106_top_grid_pin_18_;
wire [0:0] cbx_1__1__106_top_grid_pin_19_;
wire [0:0] cbx_1__1__106_top_grid_pin_20_;
wire [0:0] cbx_1__1__106_top_grid_pin_21_;
wire [0:0] cbx_1__1__106_top_grid_pin_22_;
wire [0:0] cbx_1__1__106_top_grid_pin_23_;
wire [0:0] cbx_1__1__106_top_grid_pin_24_;
wire [0:0] cbx_1__1__106_top_grid_pin_25_;
wire [0:0] cbx_1__1__106_top_grid_pin_26_;
wire [0:0] cbx_1__1__106_top_grid_pin_27_;
wire [0:0] cbx_1__1__106_top_grid_pin_28_;
wire [0:0] cbx_1__1__106_top_grid_pin_29_;
wire [0:0] cbx_1__1__106_top_grid_pin_30_;
wire [0:0] cbx_1__1__106_top_grid_pin_31_;
wire [0:0] cbx_1__1__107_ccff_tail;
wire [0:19] cbx_1__1__107_chanx_left_out;
wire [0:19] cbx_1__1__107_chanx_right_out;
wire [0:0] cbx_1__1__107_top_grid_pin_16_;
wire [0:0] cbx_1__1__107_top_grid_pin_17_;
wire [0:0] cbx_1__1__107_top_grid_pin_18_;
wire [0:0] cbx_1__1__107_top_grid_pin_19_;
wire [0:0] cbx_1__1__107_top_grid_pin_20_;
wire [0:0] cbx_1__1__107_top_grid_pin_21_;
wire [0:0] cbx_1__1__107_top_grid_pin_22_;
wire [0:0] cbx_1__1__107_top_grid_pin_23_;
wire [0:0] cbx_1__1__107_top_grid_pin_24_;
wire [0:0] cbx_1__1__107_top_grid_pin_25_;
wire [0:0] cbx_1__1__107_top_grid_pin_26_;
wire [0:0] cbx_1__1__107_top_grid_pin_27_;
wire [0:0] cbx_1__1__107_top_grid_pin_28_;
wire [0:0] cbx_1__1__107_top_grid_pin_29_;
wire [0:0] cbx_1__1__107_top_grid_pin_30_;
wire [0:0] cbx_1__1__107_top_grid_pin_31_;
wire [0:0] cbx_1__1__108_ccff_tail;
wire [0:19] cbx_1__1__108_chanx_left_out;
wire [0:19] cbx_1__1__108_chanx_right_out;
wire [0:0] cbx_1__1__108_top_grid_pin_16_;
wire [0:0] cbx_1__1__108_top_grid_pin_17_;
wire [0:0] cbx_1__1__108_top_grid_pin_18_;
wire [0:0] cbx_1__1__108_top_grid_pin_19_;
wire [0:0] cbx_1__1__108_top_grid_pin_20_;
wire [0:0] cbx_1__1__108_top_grid_pin_21_;
wire [0:0] cbx_1__1__108_top_grid_pin_22_;
wire [0:0] cbx_1__1__108_top_grid_pin_23_;
wire [0:0] cbx_1__1__108_top_grid_pin_24_;
wire [0:0] cbx_1__1__108_top_grid_pin_25_;
wire [0:0] cbx_1__1__108_top_grid_pin_26_;
wire [0:0] cbx_1__1__108_top_grid_pin_27_;
wire [0:0] cbx_1__1__108_top_grid_pin_28_;
wire [0:0] cbx_1__1__108_top_grid_pin_29_;
wire [0:0] cbx_1__1__108_top_grid_pin_30_;
wire [0:0] cbx_1__1__108_top_grid_pin_31_;
wire [0:0] cbx_1__1__109_ccff_tail;
wire [0:19] cbx_1__1__109_chanx_left_out;
wire [0:19] cbx_1__1__109_chanx_right_out;
wire [0:0] cbx_1__1__109_top_grid_pin_16_;
wire [0:0] cbx_1__1__109_top_grid_pin_17_;
wire [0:0] cbx_1__1__109_top_grid_pin_18_;
wire [0:0] cbx_1__1__109_top_grid_pin_19_;
wire [0:0] cbx_1__1__109_top_grid_pin_20_;
wire [0:0] cbx_1__1__109_top_grid_pin_21_;
wire [0:0] cbx_1__1__109_top_grid_pin_22_;
wire [0:0] cbx_1__1__109_top_grid_pin_23_;
wire [0:0] cbx_1__1__109_top_grid_pin_24_;
wire [0:0] cbx_1__1__109_top_grid_pin_25_;
wire [0:0] cbx_1__1__109_top_grid_pin_26_;
wire [0:0] cbx_1__1__109_top_grid_pin_27_;
wire [0:0] cbx_1__1__109_top_grid_pin_28_;
wire [0:0] cbx_1__1__109_top_grid_pin_29_;
wire [0:0] cbx_1__1__109_top_grid_pin_30_;
wire [0:0] cbx_1__1__109_top_grid_pin_31_;
wire [0:0] cbx_1__1__10_ccff_tail;
wire [0:19] cbx_1__1__10_chanx_left_out;
wire [0:19] cbx_1__1__10_chanx_right_out;
wire [0:0] cbx_1__1__10_top_grid_pin_16_;
wire [0:0] cbx_1__1__10_top_grid_pin_17_;
wire [0:0] cbx_1__1__10_top_grid_pin_18_;
wire [0:0] cbx_1__1__10_top_grid_pin_19_;
wire [0:0] cbx_1__1__10_top_grid_pin_20_;
wire [0:0] cbx_1__1__10_top_grid_pin_21_;
wire [0:0] cbx_1__1__10_top_grid_pin_22_;
wire [0:0] cbx_1__1__10_top_grid_pin_23_;
wire [0:0] cbx_1__1__10_top_grid_pin_24_;
wire [0:0] cbx_1__1__10_top_grid_pin_25_;
wire [0:0] cbx_1__1__10_top_grid_pin_26_;
wire [0:0] cbx_1__1__10_top_grid_pin_27_;
wire [0:0] cbx_1__1__10_top_grid_pin_28_;
wire [0:0] cbx_1__1__10_top_grid_pin_29_;
wire [0:0] cbx_1__1__10_top_grid_pin_30_;
wire [0:0] cbx_1__1__10_top_grid_pin_31_;
wire [0:0] cbx_1__1__110_ccff_tail;
wire [0:19] cbx_1__1__110_chanx_left_out;
wire [0:19] cbx_1__1__110_chanx_right_out;
wire [0:0] cbx_1__1__110_top_grid_pin_16_;
wire [0:0] cbx_1__1__110_top_grid_pin_17_;
wire [0:0] cbx_1__1__110_top_grid_pin_18_;
wire [0:0] cbx_1__1__110_top_grid_pin_19_;
wire [0:0] cbx_1__1__110_top_grid_pin_20_;
wire [0:0] cbx_1__1__110_top_grid_pin_21_;
wire [0:0] cbx_1__1__110_top_grid_pin_22_;
wire [0:0] cbx_1__1__110_top_grid_pin_23_;
wire [0:0] cbx_1__1__110_top_grid_pin_24_;
wire [0:0] cbx_1__1__110_top_grid_pin_25_;
wire [0:0] cbx_1__1__110_top_grid_pin_26_;
wire [0:0] cbx_1__1__110_top_grid_pin_27_;
wire [0:0] cbx_1__1__110_top_grid_pin_28_;
wire [0:0] cbx_1__1__110_top_grid_pin_29_;
wire [0:0] cbx_1__1__110_top_grid_pin_30_;
wire [0:0] cbx_1__1__110_top_grid_pin_31_;
wire [0:0] cbx_1__1__111_ccff_tail;
wire [0:19] cbx_1__1__111_chanx_left_out;
wire [0:19] cbx_1__1__111_chanx_right_out;
wire [0:0] cbx_1__1__111_top_grid_pin_16_;
wire [0:0] cbx_1__1__111_top_grid_pin_17_;
wire [0:0] cbx_1__1__111_top_grid_pin_18_;
wire [0:0] cbx_1__1__111_top_grid_pin_19_;
wire [0:0] cbx_1__1__111_top_grid_pin_20_;
wire [0:0] cbx_1__1__111_top_grid_pin_21_;
wire [0:0] cbx_1__1__111_top_grid_pin_22_;
wire [0:0] cbx_1__1__111_top_grid_pin_23_;
wire [0:0] cbx_1__1__111_top_grid_pin_24_;
wire [0:0] cbx_1__1__111_top_grid_pin_25_;
wire [0:0] cbx_1__1__111_top_grid_pin_26_;
wire [0:0] cbx_1__1__111_top_grid_pin_27_;
wire [0:0] cbx_1__1__111_top_grid_pin_28_;
wire [0:0] cbx_1__1__111_top_grid_pin_29_;
wire [0:0] cbx_1__1__111_top_grid_pin_30_;
wire [0:0] cbx_1__1__111_top_grid_pin_31_;
wire [0:0] cbx_1__1__112_ccff_tail;
wire [0:19] cbx_1__1__112_chanx_left_out;
wire [0:19] cbx_1__1__112_chanx_right_out;
wire [0:0] cbx_1__1__112_top_grid_pin_16_;
wire [0:0] cbx_1__1__112_top_grid_pin_17_;
wire [0:0] cbx_1__1__112_top_grid_pin_18_;
wire [0:0] cbx_1__1__112_top_grid_pin_19_;
wire [0:0] cbx_1__1__112_top_grid_pin_20_;
wire [0:0] cbx_1__1__112_top_grid_pin_21_;
wire [0:0] cbx_1__1__112_top_grid_pin_22_;
wire [0:0] cbx_1__1__112_top_grid_pin_23_;
wire [0:0] cbx_1__1__112_top_grid_pin_24_;
wire [0:0] cbx_1__1__112_top_grid_pin_25_;
wire [0:0] cbx_1__1__112_top_grid_pin_26_;
wire [0:0] cbx_1__1__112_top_grid_pin_27_;
wire [0:0] cbx_1__1__112_top_grid_pin_28_;
wire [0:0] cbx_1__1__112_top_grid_pin_29_;
wire [0:0] cbx_1__1__112_top_grid_pin_30_;
wire [0:0] cbx_1__1__112_top_grid_pin_31_;
wire [0:0] cbx_1__1__113_ccff_tail;
wire [0:19] cbx_1__1__113_chanx_left_out;
wire [0:19] cbx_1__1__113_chanx_right_out;
wire [0:0] cbx_1__1__113_top_grid_pin_16_;
wire [0:0] cbx_1__1__113_top_grid_pin_17_;
wire [0:0] cbx_1__1__113_top_grid_pin_18_;
wire [0:0] cbx_1__1__113_top_grid_pin_19_;
wire [0:0] cbx_1__1__113_top_grid_pin_20_;
wire [0:0] cbx_1__1__113_top_grid_pin_21_;
wire [0:0] cbx_1__1__113_top_grid_pin_22_;
wire [0:0] cbx_1__1__113_top_grid_pin_23_;
wire [0:0] cbx_1__1__113_top_grid_pin_24_;
wire [0:0] cbx_1__1__113_top_grid_pin_25_;
wire [0:0] cbx_1__1__113_top_grid_pin_26_;
wire [0:0] cbx_1__1__113_top_grid_pin_27_;
wire [0:0] cbx_1__1__113_top_grid_pin_28_;
wire [0:0] cbx_1__1__113_top_grid_pin_29_;
wire [0:0] cbx_1__1__113_top_grid_pin_30_;
wire [0:0] cbx_1__1__113_top_grid_pin_31_;
wire [0:0] cbx_1__1__114_ccff_tail;
wire [0:19] cbx_1__1__114_chanx_left_out;
wire [0:19] cbx_1__1__114_chanx_right_out;
wire [0:0] cbx_1__1__114_top_grid_pin_16_;
wire [0:0] cbx_1__1__114_top_grid_pin_17_;
wire [0:0] cbx_1__1__114_top_grid_pin_18_;
wire [0:0] cbx_1__1__114_top_grid_pin_19_;
wire [0:0] cbx_1__1__114_top_grid_pin_20_;
wire [0:0] cbx_1__1__114_top_grid_pin_21_;
wire [0:0] cbx_1__1__114_top_grid_pin_22_;
wire [0:0] cbx_1__1__114_top_grid_pin_23_;
wire [0:0] cbx_1__1__114_top_grid_pin_24_;
wire [0:0] cbx_1__1__114_top_grid_pin_25_;
wire [0:0] cbx_1__1__114_top_grid_pin_26_;
wire [0:0] cbx_1__1__114_top_grid_pin_27_;
wire [0:0] cbx_1__1__114_top_grid_pin_28_;
wire [0:0] cbx_1__1__114_top_grid_pin_29_;
wire [0:0] cbx_1__1__114_top_grid_pin_30_;
wire [0:0] cbx_1__1__114_top_grid_pin_31_;
wire [0:0] cbx_1__1__115_ccff_tail;
wire [0:19] cbx_1__1__115_chanx_left_out;
wire [0:19] cbx_1__1__115_chanx_right_out;
wire [0:0] cbx_1__1__115_top_grid_pin_16_;
wire [0:0] cbx_1__1__115_top_grid_pin_17_;
wire [0:0] cbx_1__1__115_top_grid_pin_18_;
wire [0:0] cbx_1__1__115_top_grid_pin_19_;
wire [0:0] cbx_1__1__115_top_grid_pin_20_;
wire [0:0] cbx_1__1__115_top_grid_pin_21_;
wire [0:0] cbx_1__1__115_top_grid_pin_22_;
wire [0:0] cbx_1__1__115_top_grid_pin_23_;
wire [0:0] cbx_1__1__115_top_grid_pin_24_;
wire [0:0] cbx_1__1__115_top_grid_pin_25_;
wire [0:0] cbx_1__1__115_top_grid_pin_26_;
wire [0:0] cbx_1__1__115_top_grid_pin_27_;
wire [0:0] cbx_1__1__115_top_grid_pin_28_;
wire [0:0] cbx_1__1__115_top_grid_pin_29_;
wire [0:0] cbx_1__1__115_top_grid_pin_30_;
wire [0:0] cbx_1__1__115_top_grid_pin_31_;
wire [0:0] cbx_1__1__116_ccff_tail;
wire [0:19] cbx_1__1__116_chanx_left_out;
wire [0:19] cbx_1__1__116_chanx_right_out;
wire [0:0] cbx_1__1__116_top_grid_pin_16_;
wire [0:0] cbx_1__1__116_top_grid_pin_17_;
wire [0:0] cbx_1__1__116_top_grid_pin_18_;
wire [0:0] cbx_1__1__116_top_grid_pin_19_;
wire [0:0] cbx_1__1__116_top_grid_pin_20_;
wire [0:0] cbx_1__1__116_top_grid_pin_21_;
wire [0:0] cbx_1__1__116_top_grid_pin_22_;
wire [0:0] cbx_1__1__116_top_grid_pin_23_;
wire [0:0] cbx_1__1__116_top_grid_pin_24_;
wire [0:0] cbx_1__1__116_top_grid_pin_25_;
wire [0:0] cbx_1__1__116_top_grid_pin_26_;
wire [0:0] cbx_1__1__116_top_grid_pin_27_;
wire [0:0] cbx_1__1__116_top_grid_pin_28_;
wire [0:0] cbx_1__1__116_top_grid_pin_29_;
wire [0:0] cbx_1__1__116_top_grid_pin_30_;
wire [0:0] cbx_1__1__116_top_grid_pin_31_;
wire [0:0] cbx_1__1__117_ccff_tail;
wire [0:19] cbx_1__1__117_chanx_left_out;
wire [0:19] cbx_1__1__117_chanx_right_out;
wire [0:0] cbx_1__1__117_top_grid_pin_16_;
wire [0:0] cbx_1__1__117_top_grid_pin_17_;
wire [0:0] cbx_1__1__117_top_grid_pin_18_;
wire [0:0] cbx_1__1__117_top_grid_pin_19_;
wire [0:0] cbx_1__1__117_top_grid_pin_20_;
wire [0:0] cbx_1__1__117_top_grid_pin_21_;
wire [0:0] cbx_1__1__117_top_grid_pin_22_;
wire [0:0] cbx_1__1__117_top_grid_pin_23_;
wire [0:0] cbx_1__1__117_top_grid_pin_24_;
wire [0:0] cbx_1__1__117_top_grid_pin_25_;
wire [0:0] cbx_1__1__117_top_grid_pin_26_;
wire [0:0] cbx_1__1__117_top_grid_pin_27_;
wire [0:0] cbx_1__1__117_top_grid_pin_28_;
wire [0:0] cbx_1__1__117_top_grid_pin_29_;
wire [0:0] cbx_1__1__117_top_grid_pin_30_;
wire [0:0] cbx_1__1__117_top_grid_pin_31_;
wire [0:0] cbx_1__1__118_ccff_tail;
wire [0:19] cbx_1__1__118_chanx_left_out;
wire [0:19] cbx_1__1__118_chanx_right_out;
wire [0:0] cbx_1__1__118_top_grid_pin_16_;
wire [0:0] cbx_1__1__118_top_grid_pin_17_;
wire [0:0] cbx_1__1__118_top_grid_pin_18_;
wire [0:0] cbx_1__1__118_top_grid_pin_19_;
wire [0:0] cbx_1__1__118_top_grid_pin_20_;
wire [0:0] cbx_1__1__118_top_grid_pin_21_;
wire [0:0] cbx_1__1__118_top_grid_pin_22_;
wire [0:0] cbx_1__1__118_top_grid_pin_23_;
wire [0:0] cbx_1__1__118_top_grid_pin_24_;
wire [0:0] cbx_1__1__118_top_grid_pin_25_;
wire [0:0] cbx_1__1__118_top_grid_pin_26_;
wire [0:0] cbx_1__1__118_top_grid_pin_27_;
wire [0:0] cbx_1__1__118_top_grid_pin_28_;
wire [0:0] cbx_1__1__118_top_grid_pin_29_;
wire [0:0] cbx_1__1__118_top_grid_pin_30_;
wire [0:0] cbx_1__1__118_top_grid_pin_31_;
wire [0:0] cbx_1__1__119_ccff_tail;
wire [0:19] cbx_1__1__119_chanx_left_out;
wire [0:19] cbx_1__1__119_chanx_right_out;
wire [0:0] cbx_1__1__119_top_grid_pin_16_;
wire [0:0] cbx_1__1__119_top_grid_pin_17_;
wire [0:0] cbx_1__1__119_top_grid_pin_18_;
wire [0:0] cbx_1__1__119_top_grid_pin_19_;
wire [0:0] cbx_1__1__119_top_grid_pin_20_;
wire [0:0] cbx_1__1__119_top_grid_pin_21_;
wire [0:0] cbx_1__1__119_top_grid_pin_22_;
wire [0:0] cbx_1__1__119_top_grid_pin_23_;
wire [0:0] cbx_1__1__119_top_grid_pin_24_;
wire [0:0] cbx_1__1__119_top_grid_pin_25_;
wire [0:0] cbx_1__1__119_top_grid_pin_26_;
wire [0:0] cbx_1__1__119_top_grid_pin_27_;
wire [0:0] cbx_1__1__119_top_grid_pin_28_;
wire [0:0] cbx_1__1__119_top_grid_pin_29_;
wire [0:0] cbx_1__1__119_top_grid_pin_30_;
wire [0:0] cbx_1__1__119_top_grid_pin_31_;
wire [0:0] cbx_1__1__11_ccff_tail;
wire [0:19] cbx_1__1__11_chanx_left_out;
wire [0:19] cbx_1__1__11_chanx_right_out;
wire [0:0] cbx_1__1__11_top_grid_pin_16_;
wire [0:0] cbx_1__1__11_top_grid_pin_17_;
wire [0:0] cbx_1__1__11_top_grid_pin_18_;
wire [0:0] cbx_1__1__11_top_grid_pin_19_;
wire [0:0] cbx_1__1__11_top_grid_pin_20_;
wire [0:0] cbx_1__1__11_top_grid_pin_21_;
wire [0:0] cbx_1__1__11_top_grid_pin_22_;
wire [0:0] cbx_1__1__11_top_grid_pin_23_;
wire [0:0] cbx_1__1__11_top_grid_pin_24_;
wire [0:0] cbx_1__1__11_top_grid_pin_25_;
wire [0:0] cbx_1__1__11_top_grid_pin_26_;
wire [0:0] cbx_1__1__11_top_grid_pin_27_;
wire [0:0] cbx_1__1__11_top_grid_pin_28_;
wire [0:0] cbx_1__1__11_top_grid_pin_29_;
wire [0:0] cbx_1__1__11_top_grid_pin_30_;
wire [0:0] cbx_1__1__11_top_grid_pin_31_;
wire [0:0] cbx_1__1__120_ccff_tail;
wire [0:19] cbx_1__1__120_chanx_left_out;
wire [0:19] cbx_1__1__120_chanx_right_out;
wire [0:0] cbx_1__1__120_top_grid_pin_16_;
wire [0:0] cbx_1__1__120_top_grid_pin_17_;
wire [0:0] cbx_1__1__120_top_grid_pin_18_;
wire [0:0] cbx_1__1__120_top_grid_pin_19_;
wire [0:0] cbx_1__1__120_top_grid_pin_20_;
wire [0:0] cbx_1__1__120_top_grid_pin_21_;
wire [0:0] cbx_1__1__120_top_grid_pin_22_;
wire [0:0] cbx_1__1__120_top_grid_pin_23_;
wire [0:0] cbx_1__1__120_top_grid_pin_24_;
wire [0:0] cbx_1__1__120_top_grid_pin_25_;
wire [0:0] cbx_1__1__120_top_grid_pin_26_;
wire [0:0] cbx_1__1__120_top_grid_pin_27_;
wire [0:0] cbx_1__1__120_top_grid_pin_28_;
wire [0:0] cbx_1__1__120_top_grid_pin_29_;
wire [0:0] cbx_1__1__120_top_grid_pin_30_;
wire [0:0] cbx_1__1__120_top_grid_pin_31_;
wire [0:0] cbx_1__1__121_ccff_tail;
wire [0:19] cbx_1__1__121_chanx_left_out;
wire [0:19] cbx_1__1__121_chanx_right_out;
wire [0:0] cbx_1__1__121_top_grid_pin_16_;
wire [0:0] cbx_1__1__121_top_grid_pin_17_;
wire [0:0] cbx_1__1__121_top_grid_pin_18_;
wire [0:0] cbx_1__1__121_top_grid_pin_19_;
wire [0:0] cbx_1__1__121_top_grid_pin_20_;
wire [0:0] cbx_1__1__121_top_grid_pin_21_;
wire [0:0] cbx_1__1__121_top_grid_pin_22_;
wire [0:0] cbx_1__1__121_top_grid_pin_23_;
wire [0:0] cbx_1__1__121_top_grid_pin_24_;
wire [0:0] cbx_1__1__121_top_grid_pin_25_;
wire [0:0] cbx_1__1__121_top_grid_pin_26_;
wire [0:0] cbx_1__1__121_top_grid_pin_27_;
wire [0:0] cbx_1__1__121_top_grid_pin_28_;
wire [0:0] cbx_1__1__121_top_grid_pin_29_;
wire [0:0] cbx_1__1__121_top_grid_pin_30_;
wire [0:0] cbx_1__1__121_top_grid_pin_31_;
wire [0:0] cbx_1__1__122_ccff_tail;
wire [0:19] cbx_1__1__122_chanx_left_out;
wire [0:19] cbx_1__1__122_chanx_right_out;
wire [0:0] cbx_1__1__122_top_grid_pin_16_;
wire [0:0] cbx_1__1__122_top_grid_pin_17_;
wire [0:0] cbx_1__1__122_top_grid_pin_18_;
wire [0:0] cbx_1__1__122_top_grid_pin_19_;
wire [0:0] cbx_1__1__122_top_grid_pin_20_;
wire [0:0] cbx_1__1__122_top_grid_pin_21_;
wire [0:0] cbx_1__1__122_top_grid_pin_22_;
wire [0:0] cbx_1__1__122_top_grid_pin_23_;
wire [0:0] cbx_1__1__122_top_grid_pin_24_;
wire [0:0] cbx_1__1__122_top_grid_pin_25_;
wire [0:0] cbx_1__1__122_top_grid_pin_26_;
wire [0:0] cbx_1__1__122_top_grid_pin_27_;
wire [0:0] cbx_1__1__122_top_grid_pin_28_;
wire [0:0] cbx_1__1__122_top_grid_pin_29_;
wire [0:0] cbx_1__1__122_top_grid_pin_30_;
wire [0:0] cbx_1__1__122_top_grid_pin_31_;
wire [0:0] cbx_1__1__123_ccff_tail;
wire [0:19] cbx_1__1__123_chanx_left_out;
wire [0:19] cbx_1__1__123_chanx_right_out;
wire [0:0] cbx_1__1__123_top_grid_pin_16_;
wire [0:0] cbx_1__1__123_top_grid_pin_17_;
wire [0:0] cbx_1__1__123_top_grid_pin_18_;
wire [0:0] cbx_1__1__123_top_grid_pin_19_;
wire [0:0] cbx_1__1__123_top_grid_pin_20_;
wire [0:0] cbx_1__1__123_top_grid_pin_21_;
wire [0:0] cbx_1__1__123_top_grid_pin_22_;
wire [0:0] cbx_1__1__123_top_grid_pin_23_;
wire [0:0] cbx_1__1__123_top_grid_pin_24_;
wire [0:0] cbx_1__1__123_top_grid_pin_25_;
wire [0:0] cbx_1__1__123_top_grid_pin_26_;
wire [0:0] cbx_1__1__123_top_grid_pin_27_;
wire [0:0] cbx_1__1__123_top_grid_pin_28_;
wire [0:0] cbx_1__1__123_top_grid_pin_29_;
wire [0:0] cbx_1__1__123_top_grid_pin_30_;
wire [0:0] cbx_1__1__123_top_grid_pin_31_;
wire [0:0] cbx_1__1__124_ccff_tail;
wire [0:19] cbx_1__1__124_chanx_left_out;
wire [0:19] cbx_1__1__124_chanx_right_out;
wire [0:0] cbx_1__1__124_top_grid_pin_16_;
wire [0:0] cbx_1__1__124_top_grid_pin_17_;
wire [0:0] cbx_1__1__124_top_grid_pin_18_;
wire [0:0] cbx_1__1__124_top_grid_pin_19_;
wire [0:0] cbx_1__1__124_top_grid_pin_20_;
wire [0:0] cbx_1__1__124_top_grid_pin_21_;
wire [0:0] cbx_1__1__124_top_grid_pin_22_;
wire [0:0] cbx_1__1__124_top_grid_pin_23_;
wire [0:0] cbx_1__1__124_top_grid_pin_24_;
wire [0:0] cbx_1__1__124_top_grid_pin_25_;
wire [0:0] cbx_1__1__124_top_grid_pin_26_;
wire [0:0] cbx_1__1__124_top_grid_pin_27_;
wire [0:0] cbx_1__1__124_top_grid_pin_28_;
wire [0:0] cbx_1__1__124_top_grid_pin_29_;
wire [0:0] cbx_1__1__124_top_grid_pin_30_;
wire [0:0] cbx_1__1__124_top_grid_pin_31_;
wire [0:0] cbx_1__1__125_ccff_tail;
wire [0:19] cbx_1__1__125_chanx_left_out;
wire [0:19] cbx_1__1__125_chanx_right_out;
wire [0:0] cbx_1__1__125_top_grid_pin_16_;
wire [0:0] cbx_1__1__125_top_grid_pin_17_;
wire [0:0] cbx_1__1__125_top_grid_pin_18_;
wire [0:0] cbx_1__1__125_top_grid_pin_19_;
wire [0:0] cbx_1__1__125_top_grid_pin_20_;
wire [0:0] cbx_1__1__125_top_grid_pin_21_;
wire [0:0] cbx_1__1__125_top_grid_pin_22_;
wire [0:0] cbx_1__1__125_top_grid_pin_23_;
wire [0:0] cbx_1__1__125_top_grid_pin_24_;
wire [0:0] cbx_1__1__125_top_grid_pin_25_;
wire [0:0] cbx_1__1__125_top_grid_pin_26_;
wire [0:0] cbx_1__1__125_top_grid_pin_27_;
wire [0:0] cbx_1__1__125_top_grid_pin_28_;
wire [0:0] cbx_1__1__125_top_grid_pin_29_;
wire [0:0] cbx_1__1__125_top_grid_pin_30_;
wire [0:0] cbx_1__1__125_top_grid_pin_31_;
wire [0:0] cbx_1__1__126_ccff_tail;
wire [0:19] cbx_1__1__126_chanx_left_out;
wire [0:19] cbx_1__1__126_chanx_right_out;
wire [0:0] cbx_1__1__126_top_grid_pin_16_;
wire [0:0] cbx_1__1__126_top_grid_pin_17_;
wire [0:0] cbx_1__1__126_top_grid_pin_18_;
wire [0:0] cbx_1__1__126_top_grid_pin_19_;
wire [0:0] cbx_1__1__126_top_grid_pin_20_;
wire [0:0] cbx_1__1__126_top_grid_pin_21_;
wire [0:0] cbx_1__1__126_top_grid_pin_22_;
wire [0:0] cbx_1__1__126_top_grid_pin_23_;
wire [0:0] cbx_1__1__126_top_grid_pin_24_;
wire [0:0] cbx_1__1__126_top_grid_pin_25_;
wire [0:0] cbx_1__1__126_top_grid_pin_26_;
wire [0:0] cbx_1__1__126_top_grid_pin_27_;
wire [0:0] cbx_1__1__126_top_grid_pin_28_;
wire [0:0] cbx_1__1__126_top_grid_pin_29_;
wire [0:0] cbx_1__1__126_top_grid_pin_30_;
wire [0:0] cbx_1__1__126_top_grid_pin_31_;
wire [0:0] cbx_1__1__127_ccff_tail;
wire [0:19] cbx_1__1__127_chanx_left_out;
wire [0:19] cbx_1__1__127_chanx_right_out;
wire [0:0] cbx_1__1__127_top_grid_pin_16_;
wire [0:0] cbx_1__1__127_top_grid_pin_17_;
wire [0:0] cbx_1__1__127_top_grid_pin_18_;
wire [0:0] cbx_1__1__127_top_grid_pin_19_;
wire [0:0] cbx_1__1__127_top_grid_pin_20_;
wire [0:0] cbx_1__1__127_top_grid_pin_21_;
wire [0:0] cbx_1__1__127_top_grid_pin_22_;
wire [0:0] cbx_1__1__127_top_grid_pin_23_;
wire [0:0] cbx_1__1__127_top_grid_pin_24_;
wire [0:0] cbx_1__1__127_top_grid_pin_25_;
wire [0:0] cbx_1__1__127_top_grid_pin_26_;
wire [0:0] cbx_1__1__127_top_grid_pin_27_;
wire [0:0] cbx_1__1__127_top_grid_pin_28_;
wire [0:0] cbx_1__1__127_top_grid_pin_29_;
wire [0:0] cbx_1__1__127_top_grid_pin_30_;
wire [0:0] cbx_1__1__127_top_grid_pin_31_;
wire [0:0] cbx_1__1__128_ccff_tail;
wire [0:19] cbx_1__1__128_chanx_left_out;
wire [0:19] cbx_1__1__128_chanx_right_out;
wire [0:0] cbx_1__1__128_top_grid_pin_16_;
wire [0:0] cbx_1__1__128_top_grid_pin_17_;
wire [0:0] cbx_1__1__128_top_grid_pin_18_;
wire [0:0] cbx_1__1__128_top_grid_pin_19_;
wire [0:0] cbx_1__1__128_top_grid_pin_20_;
wire [0:0] cbx_1__1__128_top_grid_pin_21_;
wire [0:0] cbx_1__1__128_top_grid_pin_22_;
wire [0:0] cbx_1__1__128_top_grid_pin_23_;
wire [0:0] cbx_1__1__128_top_grid_pin_24_;
wire [0:0] cbx_1__1__128_top_grid_pin_25_;
wire [0:0] cbx_1__1__128_top_grid_pin_26_;
wire [0:0] cbx_1__1__128_top_grid_pin_27_;
wire [0:0] cbx_1__1__128_top_grid_pin_28_;
wire [0:0] cbx_1__1__128_top_grid_pin_29_;
wire [0:0] cbx_1__1__128_top_grid_pin_30_;
wire [0:0] cbx_1__1__128_top_grid_pin_31_;
wire [0:0] cbx_1__1__129_ccff_tail;
wire [0:19] cbx_1__1__129_chanx_left_out;
wire [0:19] cbx_1__1__129_chanx_right_out;
wire [0:0] cbx_1__1__129_top_grid_pin_16_;
wire [0:0] cbx_1__1__129_top_grid_pin_17_;
wire [0:0] cbx_1__1__129_top_grid_pin_18_;
wire [0:0] cbx_1__1__129_top_grid_pin_19_;
wire [0:0] cbx_1__1__129_top_grid_pin_20_;
wire [0:0] cbx_1__1__129_top_grid_pin_21_;
wire [0:0] cbx_1__1__129_top_grid_pin_22_;
wire [0:0] cbx_1__1__129_top_grid_pin_23_;
wire [0:0] cbx_1__1__129_top_grid_pin_24_;
wire [0:0] cbx_1__1__129_top_grid_pin_25_;
wire [0:0] cbx_1__1__129_top_grid_pin_26_;
wire [0:0] cbx_1__1__129_top_grid_pin_27_;
wire [0:0] cbx_1__1__129_top_grid_pin_28_;
wire [0:0] cbx_1__1__129_top_grid_pin_29_;
wire [0:0] cbx_1__1__129_top_grid_pin_30_;
wire [0:0] cbx_1__1__129_top_grid_pin_31_;
wire [0:0] cbx_1__1__12_ccff_tail;
wire [0:19] cbx_1__1__12_chanx_left_out;
wire [0:19] cbx_1__1__12_chanx_right_out;
wire [0:0] cbx_1__1__12_top_grid_pin_16_;
wire [0:0] cbx_1__1__12_top_grid_pin_17_;
wire [0:0] cbx_1__1__12_top_grid_pin_18_;
wire [0:0] cbx_1__1__12_top_grid_pin_19_;
wire [0:0] cbx_1__1__12_top_grid_pin_20_;
wire [0:0] cbx_1__1__12_top_grid_pin_21_;
wire [0:0] cbx_1__1__12_top_grid_pin_22_;
wire [0:0] cbx_1__1__12_top_grid_pin_23_;
wire [0:0] cbx_1__1__12_top_grid_pin_24_;
wire [0:0] cbx_1__1__12_top_grid_pin_25_;
wire [0:0] cbx_1__1__12_top_grid_pin_26_;
wire [0:0] cbx_1__1__12_top_grid_pin_27_;
wire [0:0] cbx_1__1__12_top_grid_pin_28_;
wire [0:0] cbx_1__1__12_top_grid_pin_29_;
wire [0:0] cbx_1__1__12_top_grid_pin_30_;
wire [0:0] cbx_1__1__12_top_grid_pin_31_;
wire [0:0] cbx_1__1__130_ccff_tail;
wire [0:19] cbx_1__1__130_chanx_left_out;
wire [0:19] cbx_1__1__130_chanx_right_out;
wire [0:0] cbx_1__1__130_top_grid_pin_16_;
wire [0:0] cbx_1__1__130_top_grid_pin_17_;
wire [0:0] cbx_1__1__130_top_grid_pin_18_;
wire [0:0] cbx_1__1__130_top_grid_pin_19_;
wire [0:0] cbx_1__1__130_top_grid_pin_20_;
wire [0:0] cbx_1__1__130_top_grid_pin_21_;
wire [0:0] cbx_1__1__130_top_grid_pin_22_;
wire [0:0] cbx_1__1__130_top_grid_pin_23_;
wire [0:0] cbx_1__1__130_top_grid_pin_24_;
wire [0:0] cbx_1__1__130_top_grid_pin_25_;
wire [0:0] cbx_1__1__130_top_grid_pin_26_;
wire [0:0] cbx_1__1__130_top_grid_pin_27_;
wire [0:0] cbx_1__1__130_top_grid_pin_28_;
wire [0:0] cbx_1__1__130_top_grid_pin_29_;
wire [0:0] cbx_1__1__130_top_grid_pin_30_;
wire [0:0] cbx_1__1__130_top_grid_pin_31_;
wire [0:0] cbx_1__1__131_ccff_tail;
wire [0:19] cbx_1__1__131_chanx_left_out;
wire [0:19] cbx_1__1__131_chanx_right_out;
wire [0:0] cbx_1__1__131_top_grid_pin_16_;
wire [0:0] cbx_1__1__131_top_grid_pin_17_;
wire [0:0] cbx_1__1__131_top_grid_pin_18_;
wire [0:0] cbx_1__1__131_top_grid_pin_19_;
wire [0:0] cbx_1__1__131_top_grid_pin_20_;
wire [0:0] cbx_1__1__131_top_grid_pin_21_;
wire [0:0] cbx_1__1__131_top_grid_pin_22_;
wire [0:0] cbx_1__1__131_top_grid_pin_23_;
wire [0:0] cbx_1__1__131_top_grid_pin_24_;
wire [0:0] cbx_1__1__131_top_grid_pin_25_;
wire [0:0] cbx_1__1__131_top_grid_pin_26_;
wire [0:0] cbx_1__1__131_top_grid_pin_27_;
wire [0:0] cbx_1__1__131_top_grid_pin_28_;
wire [0:0] cbx_1__1__131_top_grid_pin_29_;
wire [0:0] cbx_1__1__131_top_grid_pin_30_;
wire [0:0] cbx_1__1__131_top_grid_pin_31_;
wire [0:0] cbx_1__1__13_ccff_tail;
wire [0:19] cbx_1__1__13_chanx_left_out;
wire [0:19] cbx_1__1__13_chanx_right_out;
wire [0:0] cbx_1__1__13_top_grid_pin_16_;
wire [0:0] cbx_1__1__13_top_grid_pin_17_;
wire [0:0] cbx_1__1__13_top_grid_pin_18_;
wire [0:0] cbx_1__1__13_top_grid_pin_19_;
wire [0:0] cbx_1__1__13_top_grid_pin_20_;
wire [0:0] cbx_1__1__13_top_grid_pin_21_;
wire [0:0] cbx_1__1__13_top_grid_pin_22_;
wire [0:0] cbx_1__1__13_top_grid_pin_23_;
wire [0:0] cbx_1__1__13_top_grid_pin_24_;
wire [0:0] cbx_1__1__13_top_grid_pin_25_;
wire [0:0] cbx_1__1__13_top_grid_pin_26_;
wire [0:0] cbx_1__1__13_top_grid_pin_27_;
wire [0:0] cbx_1__1__13_top_grid_pin_28_;
wire [0:0] cbx_1__1__13_top_grid_pin_29_;
wire [0:0] cbx_1__1__13_top_grid_pin_30_;
wire [0:0] cbx_1__1__13_top_grid_pin_31_;
wire [0:0] cbx_1__1__14_ccff_tail;
wire [0:19] cbx_1__1__14_chanx_left_out;
wire [0:19] cbx_1__1__14_chanx_right_out;
wire [0:0] cbx_1__1__14_top_grid_pin_16_;
wire [0:0] cbx_1__1__14_top_grid_pin_17_;
wire [0:0] cbx_1__1__14_top_grid_pin_18_;
wire [0:0] cbx_1__1__14_top_grid_pin_19_;
wire [0:0] cbx_1__1__14_top_grid_pin_20_;
wire [0:0] cbx_1__1__14_top_grid_pin_21_;
wire [0:0] cbx_1__1__14_top_grid_pin_22_;
wire [0:0] cbx_1__1__14_top_grid_pin_23_;
wire [0:0] cbx_1__1__14_top_grid_pin_24_;
wire [0:0] cbx_1__1__14_top_grid_pin_25_;
wire [0:0] cbx_1__1__14_top_grid_pin_26_;
wire [0:0] cbx_1__1__14_top_grid_pin_27_;
wire [0:0] cbx_1__1__14_top_grid_pin_28_;
wire [0:0] cbx_1__1__14_top_grid_pin_29_;
wire [0:0] cbx_1__1__14_top_grid_pin_30_;
wire [0:0] cbx_1__1__14_top_grid_pin_31_;
wire [0:0] cbx_1__1__15_ccff_tail;
wire [0:19] cbx_1__1__15_chanx_left_out;
wire [0:19] cbx_1__1__15_chanx_right_out;
wire [0:0] cbx_1__1__15_top_grid_pin_16_;
wire [0:0] cbx_1__1__15_top_grid_pin_17_;
wire [0:0] cbx_1__1__15_top_grid_pin_18_;
wire [0:0] cbx_1__1__15_top_grid_pin_19_;
wire [0:0] cbx_1__1__15_top_grid_pin_20_;
wire [0:0] cbx_1__1__15_top_grid_pin_21_;
wire [0:0] cbx_1__1__15_top_grid_pin_22_;
wire [0:0] cbx_1__1__15_top_grid_pin_23_;
wire [0:0] cbx_1__1__15_top_grid_pin_24_;
wire [0:0] cbx_1__1__15_top_grid_pin_25_;
wire [0:0] cbx_1__1__15_top_grid_pin_26_;
wire [0:0] cbx_1__1__15_top_grid_pin_27_;
wire [0:0] cbx_1__1__15_top_grid_pin_28_;
wire [0:0] cbx_1__1__15_top_grid_pin_29_;
wire [0:0] cbx_1__1__15_top_grid_pin_30_;
wire [0:0] cbx_1__1__15_top_grid_pin_31_;
wire [0:0] cbx_1__1__16_ccff_tail;
wire [0:19] cbx_1__1__16_chanx_left_out;
wire [0:19] cbx_1__1__16_chanx_right_out;
wire [0:0] cbx_1__1__16_top_grid_pin_16_;
wire [0:0] cbx_1__1__16_top_grid_pin_17_;
wire [0:0] cbx_1__1__16_top_grid_pin_18_;
wire [0:0] cbx_1__1__16_top_grid_pin_19_;
wire [0:0] cbx_1__1__16_top_grid_pin_20_;
wire [0:0] cbx_1__1__16_top_grid_pin_21_;
wire [0:0] cbx_1__1__16_top_grid_pin_22_;
wire [0:0] cbx_1__1__16_top_grid_pin_23_;
wire [0:0] cbx_1__1__16_top_grid_pin_24_;
wire [0:0] cbx_1__1__16_top_grid_pin_25_;
wire [0:0] cbx_1__1__16_top_grid_pin_26_;
wire [0:0] cbx_1__1__16_top_grid_pin_27_;
wire [0:0] cbx_1__1__16_top_grid_pin_28_;
wire [0:0] cbx_1__1__16_top_grid_pin_29_;
wire [0:0] cbx_1__1__16_top_grid_pin_30_;
wire [0:0] cbx_1__1__16_top_grid_pin_31_;
wire [0:0] cbx_1__1__17_ccff_tail;
wire [0:19] cbx_1__1__17_chanx_left_out;
wire [0:19] cbx_1__1__17_chanx_right_out;
wire [0:0] cbx_1__1__17_top_grid_pin_16_;
wire [0:0] cbx_1__1__17_top_grid_pin_17_;
wire [0:0] cbx_1__1__17_top_grid_pin_18_;
wire [0:0] cbx_1__1__17_top_grid_pin_19_;
wire [0:0] cbx_1__1__17_top_grid_pin_20_;
wire [0:0] cbx_1__1__17_top_grid_pin_21_;
wire [0:0] cbx_1__1__17_top_grid_pin_22_;
wire [0:0] cbx_1__1__17_top_grid_pin_23_;
wire [0:0] cbx_1__1__17_top_grid_pin_24_;
wire [0:0] cbx_1__1__17_top_grid_pin_25_;
wire [0:0] cbx_1__1__17_top_grid_pin_26_;
wire [0:0] cbx_1__1__17_top_grid_pin_27_;
wire [0:0] cbx_1__1__17_top_grid_pin_28_;
wire [0:0] cbx_1__1__17_top_grid_pin_29_;
wire [0:0] cbx_1__1__17_top_grid_pin_30_;
wire [0:0] cbx_1__1__17_top_grid_pin_31_;
wire [0:0] cbx_1__1__18_ccff_tail;
wire [0:19] cbx_1__1__18_chanx_left_out;
wire [0:19] cbx_1__1__18_chanx_right_out;
wire [0:0] cbx_1__1__18_top_grid_pin_16_;
wire [0:0] cbx_1__1__18_top_grid_pin_17_;
wire [0:0] cbx_1__1__18_top_grid_pin_18_;
wire [0:0] cbx_1__1__18_top_grid_pin_19_;
wire [0:0] cbx_1__1__18_top_grid_pin_20_;
wire [0:0] cbx_1__1__18_top_grid_pin_21_;
wire [0:0] cbx_1__1__18_top_grid_pin_22_;
wire [0:0] cbx_1__1__18_top_grid_pin_23_;
wire [0:0] cbx_1__1__18_top_grid_pin_24_;
wire [0:0] cbx_1__1__18_top_grid_pin_25_;
wire [0:0] cbx_1__1__18_top_grid_pin_26_;
wire [0:0] cbx_1__1__18_top_grid_pin_27_;
wire [0:0] cbx_1__1__18_top_grid_pin_28_;
wire [0:0] cbx_1__1__18_top_grid_pin_29_;
wire [0:0] cbx_1__1__18_top_grid_pin_30_;
wire [0:0] cbx_1__1__18_top_grid_pin_31_;
wire [0:0] cbx_1__1__19_ccff_tail;
wire [0:19] cbx_1__1__19_chanx_left_out;
wire [0:19] cbx_1__1__19_chanx_right_out;
wire [0:0] cbx_1__1__19_top_grid_pin_16_;
wire [0:0] cbx_1__1__19_top_grid_pin_17_;
wire [0:0] cbx_1__1__19_top_grid_pin_18_;
wire [0:0] cbx_1__1__19_top_grid_pin_19_;
wire [0:0] cbx_1__1__19_top_grid_pin_20_;
wire [0:0] cbx_1__1__19_top_grid_pin_21_;
wire [0:0] cbx_1__1__19_top_grid_pin_22_;
wire [0:0] cbx_1__1__19_top_grid_pin_23_;
wire [0:0] cbx_1__1__19_top_grid_pin_24_;
wire [0:0] cbx_1__1__19_top_grid_pin_25_;
wire [0:0] cbx_1__1__19_top_grid_pin_26_;
wire [0:0] cbx_1__1__19_top_grid_pin_27_;
wire [0:0] cbx_1__1__19_top_grid_pin_28_;
wire [0:0] cbx_1__1__19_top_grid_pin_29_;
wire [0:0] cbx_1__1__19_top_grid_pin_30_;
wire [0:0] cbx_1__1__19_top_grid_pin_31_;
wire [0:0] cbx_1__1__1_ccff_tail;
wire [0:19] cbx_1__1__1_chanx_left_out;
wire [0:19] cbx_1__1__1_chanx_right_out;
wire [0:0] cbx_1__1__1_top_grid_pin_16_;
wire [0:0] cbx_1__1__1_top_grid_pin_17_;
wire [0:0] cbx_1__1__1_top_grid_pin_18_;
wire [0:0] cbx_1__1__1_top_grid_pin_19_;
wire [0:0] cbx_1__1__1_top_grid_pin_20_;
wire [0:0] cbx_1__1__1_top_grid_pin_21_;
wire [0:0] cbx_1__1__1_top_grid_pin_22_;
wire [0:0] cbx_1__1__1_top_grid_pin_23_;
wire [0:0] cbx_1__1__1_top_grid_pin_24_;
wire [0:0] cbx_1__1__1_top_grid_pin_25_;
wire [0:0] cbx_1__1__1_top_grid_pin_26_;
wire [0:0] cbx_1__1__1_top_grid_pin_27_;
wire [0:0] cbx_1__1__1_top_grid_pin_28_;
wire [0:0] cbx_1__1__1_top_grid_pin_29_;
wire [0:0] cbx_1__1__1_top_grid_pin_30_;
wire [0:0] cbx_1__1__1_top_grid_pin_31_;
wire [0:0] cbx_1__1__20_ccff_tail;
wire [0:19] cbx_1__1__20_chanx_left_out;
wire [0:19] cbx_1__1__20_chanx_right_out;
wire [0:0] cbx_1__1__20_top_grid_pin_16_;
wire [0:0] cbx_1__1__20_top_grid_pin_17_;
wire [0:0] cbx_1__1__20_top_grid_pin_18_;
wire [0:0] cbx_1__1__20_top_grid_pin_19_;
wire [0:0] cbx_1__1__20_top_grid_pin_20_;
wire [0:0] cbx_1__1__20_top_grid_pin_21_;
wire [0:0] cbx_1__1__20_top_grid_pin_22_;
wire [0:0] cbx_1__1__20_top_grid_pin_23_;
wire [0:0] cbx_1__1__20_top_grid_pin_24_;
wire [0:0] cbx_1__1__20_top_grid_pin_25_;
wire [0:0] cbx_1__1__20_top_grid_pin_26_;
wire [0:0] cbx_1__1__20_top_grid_pin_27_;
wire [0:0] cbx_1__1__20_top_grid_pin_28_;
wire [0:0] cbx_1__1__20_top_grid_pin_29_;
wire [0:0] cbx_1__1__20_top_grid_pin_30_;
wire [0:0] cbx_1__1__20_top_grid_pin_31_;
wire [0:0] cbx_1__1__21_ccff_tail;
wire [0:19] cbx_1__1__21_chanx_left_out;
wire [0:19] cbx_1__1__21_chanx_right_out;
wire [0:0] cbx_1__1__21_top_grid_pin_16_;
wire [0:0] cbx_1__1__21_top_grid_pin_17_;
wire [0:0] cbx_1__1__21_top_grid_pin_18_;
wire [0:0] cbx_1__1__21_top_grid_pin_19_;
wire [0:0] cbx_1__1__21_top_grid_pin_20_;
wire [0:0] cbx_1__1__21_top_grid_pin_21_;
wire [0:0] cbx_1__1__21_top_grid_pin_22_;
wire [0:0] cbx_1__1__21_top_grid_pin_23_;
wire [0:0] cbx_1__1__21_top_grid_pin_24_;
wire [0:0] cbx_1__1__21_top_grid_pin_25_;
wire [0:0] cbx_1__1__21_top_grid_pin_26_;
wire [0:0] cbx_1__1__21_top_grid_pin_27_;
wire [0:0] cbx_1__1__21_top_grid_pin_28_;
wire [0:0] cbx_1__1__21_top_grid_pin_29_;
wire [0:0] cbx_1__1__21_top_grid_pin_30_;
wire [0:0] cbx_1__1__21_top_grid_pin_31_;
wire [0:0] cbx_1__1__22_ccff_tail;
wire [0:19] cbx_1__1__22_chanx_left_out;
wire [0:19] cbx_1__1__22_chanx_right_out;
wire [0:0] cbx_1__1__22_top_grid_pin_16_;
wire [0:0] cbx_1__1__22_top_grid_pin_17_;
wire [0:0] cbx_1__1__22_top_grid_pin_18_;
wire [0:0] cbx_1__1__22_top_grid_pin_19_;
wire [0:0] cbx_1__1__22_top_grid_pin_20_;
wire [0:0] cbx_1__1__22_top_grid_pin_21_;
wire [0:0] cbx_1__1__22_top_grid_pin_22_;
wire [0:0] cbx_1__1__22_top_grid_pin_23_;
wire [0:0] cbx_1__1__22_top_grid_pin_24_;
wire [0:0] cbx_1__1__22_top_grid_pin_25_;
wire [0:0] cbx_1__1__22_top_grid_pin_26_;
wire [0:0] cbx_1__1__22_top_grid_pin_27_;
wire [0:0] cbx_1__1__22_top_grid_pin_28_;
wire [0:0] cbx_1__1__22_top_grid_pin_29_;
wire [0:0] cbx_1__1__22_top_grid_pin_30_;
wire [0:0] cbx_1__1__22_top_grid_pin_31_;
wire [0:0] cbx_1__1__23_ccff_tail;
wire [0:19] cbx_1__1__23_chanx_left_out;
wire [0:19] cbx_1__1__23_chanx_right_out;
wire [0:0] cbx_1__1__23_top_grid_pin_16_;
wire [0:0] cbx_1__1__23_top_grid_pin_17_;
wire [0:0] cbx_1__1__23_top_grid_pin_18_;
wire [0:0] cbx_1__1__23_top_grid_pin_19_;
wire [0:0] cbx_1__1__23_top_grid_pin_20_;
wire [0:0] cbx_1__1__23_top_grid_pin_21_;
wire [0:0] cbx_1__1__23_top_grid_pin_22_;
wire [0:0] cbx_1__1__23_top_grid_pin_23_;
wire [0:0] cbx_1__1__23_top_grid_pin_24_;
wire [0:0] cbx_1__1__23_top_grid_pin_25_;
wire [0:0] cbx_1__1__23_top_grid_pin_26_;
wire [0:0] cbx_1__1__23_top_grid_pin_27_;
wire [0:0] cbx_1__1__23_top_grid_pin_28_;
wire [0:0] cbx_1__1__23_top_grid_pin_29_;
wire [0:0] cbx_1__1__23_top_grid_pin_30_;
wire [0:0] cbx_1__1__23_top_grid_pin_31_;
wire [0:0] cbx_1__1__24_ccff_tail;
wire [0:19] cbx_1__1__24_chanx_left_out;
wire [0:19] cbx_1__1__24_chanx_right_out;
wire [0:0] cbx_1__1__24_top_grid_pin_16_;
wire [0:0] cbx_1__1__24_top_grid_pin_17_;
wire [0:0] cbx_1__1__24_top_grid_pin_18_;
wire [0:0] cbx_1__1__24_top_grid_pin_19_;
wire [0:0] cbx_1__1__24_top_grid_pin_20_;
wire [0:0] cbx_1__1__24_top_grid_pin_21_;
wire [0:0] cbx_1__1__24_top_grid_pin_22_;
wire [0:0] cbx_1__1__24_top_grid_pin_23_;
wire [0:0] cbx_1__1__24_top_grid_pin_24_;
wire [0:0] cbx_1__1__24_top_grid_pin_25_;
wire [0:0] cbx_1__1__24_top_grid_pin_26_;
wire [0:0] cbx_1__1__24_top_grid_pin_27_;
wire [0:0] cbx_1__1__24_top_grid_pin_28_;
wire [0:0] cbx_1__1__24_top_grid_pin_29_;
wire [0:0] cbx_1__1__24_top_grid_pin_30_;
wire [0:0] cbx_1__1__24_top_grid_pin_31_;
wire [0:0] cbx_1__1__25_ccff_tail;
wire [0:19] cbx_1__1__25_chanx_left_out;
wire [0:19] cbx_1__1__25_chanx_right_out;
wire [0:0] cbx_1__1__25_top_grid_pin_16_;
wire [0:0] cbx_1__1__25_top_grid_pin_17_;
wire [0:0] cbx_1__1__25_top_grid_pin_18_;
wire [0:0] cbx_1__1__25_top_grid_pin_19_;
wire [0:0] cbx_1__1__25_top_grid_pin_20_;
wire [0:0] cbx_1__1__25_top_grid_pin_21_;
wire [0:0] cbx_1__1__25_top_grid_pin_22_;
wire [0:0] cbx_1__1__25_top_grid_pin_23_;
wire [0:0] cbx_1__1__25_top_grid_pin_24_;
wire [0:0] cbx_1__1__25_top_grid_pin_25_;
wire [0:0] cbx_1__1__25_top_grid_pin_26_;
wire [0:0] cbx_1__1__25_top_grid_pin_27_;
wire [0:0] cbx_1__1__25_top_grid_pin_28_;
wire [0:0] cbx_1__1__25_top_grid_pin_29_;
wire [0:0] cbx_1__1__25_top_grid_pin_30_;
wire [0:0] cbx_1__1__25_top_grid_pin_31_;
wire [0:0] cbx_1__1__26_ccff_tail;
wire [0:19] cbx_1__1__26_chanx_left_out;
wire [0:19] cbx_1__1__26_chanx_right_out;
wire [0:0] cbx_1__1__26_top_grid_pin_16_;
wire [0:0] cbx_1__1__26_top_grid_pin_17_;
wire [0:0] cbx_1__1__26_top_grid_pin_18_;
wire [0:0] cbx_1__1__26_top_grid_pin_19_;
wire [0:0] cbx_1__1__26_top_grid_pin_20_;
wire [0:0] cbx_1__1__26_top_grid_pin_21_;
wire [0:0] cbx_1__1__26_top_grid_pin_22_;
wire [0:0] cbx_1__1__26_top_grid_pin_23_;
wire [0:0] cbx_1__1__26_top_grid_pin_24_;
wire [0:0] cbx_1__1__26_top_grid_pin_25_;
wire [0:0] cbx_1__1__26_top_grid_pin_26_;
wire [0:0] cbx_1__1__26_top_grid_pin_27_;
wire [0:0] cbx_1__1__26_top_grid_pin_28_;
wire [0:0] cbx_1__1__26_top_grid_pin_29_;
wire [0:0] cbx_1__1__26_top_grid_pin_30_;
wire [0:0] cbx_1__1__26_top_grid_pin_31_;
wire [0:0] cbx_1__1__27_ccff_tail;
wire [0:19] cbx_1__1__27_chanx_left_out;
wire [0:19] cbx_1__1__27_chanx_right_out;
wire [0:0] cbx_1__1__27_top_grid_pin_16_;
wire [0:0] cbx_1__1__27_top_grid_pin_17_;
wire [0:0] cbx_1__1__27_top_grid_pin_18_;
wire [0:0] cbx_1__1__27_top_grid_pin_19_;
wire [0:0] cbx_1__1__27_top_grid_pin_20_;
wire [0:0] cbx_1__1__27_top_grid_pin_21_;
wire [0:0] cbx_1__1__27_top_grid_pin_22_;
wire [0:0] cbx_1__1__27_top_grid_pin_23_;
wire [0:0] cbx_1__1__27_top_grid_pin_24_;
wire [0:0] cbx_1__1__27_top_grid_pin_25_;
wire [0:0] cbx_1__1__27_top_grid_pin_26_;
wire [0:0] cbx_1__1__27_top_grid_pin_27_;
wire [0:0] cbx_1__1__27_top_grid_pin_28_;
wire [0:0] cbx_1__1__27_top_grid_pin_29_;
wire [0:0] cbx_1__1__27_top_grid_pin_30_;
wire [0:0] cbx_1__1__27_top_grid_pin_31_;
wire [0:0] cbx_1__1__28_ccff_tail;
wire [0:19] cbx_1__1__28_chanx_left_out;
wire [0:19] cbx_1__1__28_chanx_right_out;
wire [0:0] cbx_1__1__28_top_grid_pin_16_;
wire [0:0] cbx_1__1__28_top_grid_pin_17_;
wire [0:0] cbx_1__1__28_top_grid_pin_18_;
wire [0:0] cbx_1__1__28_top_grid_pin_19_;
wire [0:0] cbx_1__1__28_top_grid_pin_20_;
wire [0:0] cbx_1__1__28_top_grid_pin_21_;
wire [0:0] cbx_1__1__28_top_grid_pin_22_;
wire [0:0] cbx_1__1__28_top_grid_pin_23_;
wire [0:0] cbx_1__1__28_top_grid_pin_24_;
wire [0:0] cbx_1__1__28_top_grid_pin_25_;
wire [0:0] cbx_1__1__28_top_grid_pin_26_;
wire [0:0] cbx_1__1__28_top_grid_pin_27_;
wire [0:0] cbx_1__1__28_top_grid_pin_28_;
wire [0:0] cbx_1__1__28_top_grid_pin_29_;
wire [0:0] cbx_1__1__28_top_grid_pin_30_;
wire [0:0] cbx_1__1__28_top_grid_pin_31_;
wire [0:0] cbx_1__1__29_ccff_tail;
wire [0:19] cbx_1__1__29_chanx_left_out;
wire [0:19] cbx_1__1__29_chanx_right_out;
wire [0:0] cbx_1__1__29_top_grid_pin_16_;
wire [0:0] cbx_1__1__29_top_grid_pin_17_;
wire [0:0] cbx_1__1__29_top_grid_pin_18_;
wire [0:0] cbx_1__1__29_top_grid_pin_19_;
wire [0:0] cbx_1__1__29_top_grid_pin_20_;
wire [0:0] cbx_1__1__29_top_grid_pin_21_;
wire [0:0] cbx_1__1__29_top_grid_pin_22_;
wire [0:0] cbx_1__1__29_top_grid_pin_23_;
wire [0:0] cbx_1__1__29_top_grid_pin_24_;
wire [0:0] cbx_1__1__29_top_grid_pin_25_;
wire [0:0] cbx_1__1__29_top_grid_pin_26_;
wire [0:0] cbx_1__1__29_top_grid_pin_27_;
wire [0:0] cbx_1__1__29_top_grid_pin_28_;
wire [0:0] cbx_1__1__29_top_grid_pin_29_;
wire [0:0] cbx_1__1__29_top_grid_pin_30_;
wire [0:0] cbx_1__1__29_top_grid_pin_31_;
wire [0:0] cbx_1__1__2_ccff_tail;
wire [0:19] cbx_1__1__2_chanx_left_out;
wire [0:19] cbx_1__1__2_chanx_right_out;
wire [0:0] cbx_1__1__2_top_grid_pin_16_;
wire [0:0] cbx_1__1__2_top_grid_pin_17_;
wire [0:0] cbx_1__1__2_top_grid_pin_18_;
wire [0:0] cbx_1__1__2_top_grid_pin_19_;
wire [0:0] cbx_1__1__2_top_grid_pin_20_;
wire [0:0] cbx_1__1__2_top_grid_pin_21_;
wire [0:0] cbx_1__1__2_top_grid_pin_22_;
wire [0:0] cbx_1__1__2_top_grid_pin_23_;
wire [0:0] cbx_1__1__2_top_grid_pin_24_;
wire [0:0] cbx_1__1__2_top_grid_pin_25_;
wire [0:0] cbx_1__1__2_top_grid_pin_26_;
wire [0:0] cbx_1__1__2_top_grid_pin_27_;
wire [0:0] cbx_1__1__2_top_grid_pin_28_;
wire [0:0] cbx_1__1__2_top_grid_pin_29_;
wire [0:0] cbx_1__1__2_top_grid_pin_30_;
wire [0:0] cbx_1__1__2_top_grid_pin_31_;
wire [0:0] cbx_1__1__30_ccff_tail;
wire [0:19] cbx_1__1__30_chanx_left_out;
wire [0:19] cbx_1__1__30_chanx_right_out;
wire [0:0] cbx_1__1__30_top_grid_pin_16_;
wire [0:0] cbx_1__1__30_top_grid_pin_17_;
wire [0:0] cbx_1__1__30_top_grid_pin_18_;
wire [0:0] cbx_1__1__30_top_grid_pin_19_;
wire [0:0] cbx_1__1__30_top_grid_pin_20_;
wire [0:0] cbx_1__1__30_top_grid_pin_21_;
wire [0:0] cbx_1__1__30_top_grid_pin_22_;
wire [0:0] cbx_1__1__30_top_grid_pin_23_;
wire [0:0] cbx_1__1__30_top_grid_pin_24_;
wire [0:0] cbx_1__1__30_top_grid_pin_25_;
wire [0:0] cbx_1__1__30_top_grid_pin_26_;
wire [0:0] cbx_1__1__30_top_grid_pin_27_;
wire [0:0] cbx_1__1__30_top_grid_pin_28_;
wire [0:0] cbx_1__1__30_top_grid_pin_29_;
wire [0:0] cbx_1__1__30_top_grid_pin_30_;
wire [0:0] cbx_1__1__30_top_grid_pin_31_;
wire [0:0] cbx_1__1__31_ccff_tail;
wire [0:19] cbx_1__1__31_chanx_left_out;
wire [0:19] cbx_1__1__31_chanx_right_out;
wire [0:0] cbx_1__1__31_top_grid_pin_16_;
wire [0:0] cbx_1__1__31_top_grid_pin_17_;
wire [0:0] cbx_1__1__31_top_grid_pin_18_;
wire [0:0] cbx_1__1__31_top_grid_pin_19_;
wire [0:0] cbx_1__1__31_top_grid_pin_20_;
wire [0:0] cbx_1__1__31_top_grid_pin_21_;
wire [0:0] cbx_1__1__31_top_grid_pin_22_;
wire [0:0] cbx_1__1__31_top_grid_pin_23_;
wire [0:0] cbx_1__1__31_top_grid_pin_24_;
wire [0:0] cbx_1__1__31_top_grid_pin_25_;
wire [0:0] cbx_1__1__31_top_grid_pin_26_;
wire [0:0] cbx_1__1__31_top_grid_pin_27_;
wire [0:0] cbx_1__1__31_top_grid_pin_28_;
wire [0:0] cbx_1__1__31_top_grid_pin_29_;
wire [0:0] cbx_1__1__31_top_grid_pin_30_;
wire [0:0] cbx_1__1__31_top_grid_pin_31_;
wire [0:0] cbx_1__1__32_ccff_tail;
wire [0:19] cbx_1__1__32_chanx_left_out;
wire [0:19] cbx_1__1__32_chanx_right_out;
wire [0:0] cbx_1__1__32_top_grid_pin_16_;
wire [0:0] cbx_1__1__32_top_grid_pin_17_;
wire [0:0] cbx_1__1__32_top_grid_pin_18_;
wire [0:0] cbx_1__1__32_top_grid_pin_19_;
wire [0:0] cbx_1__1__32_top_grid_pin_20_;
wire [0:0] cbx_1__1__32_top_grid_pin_21_;
wire [0:0] cbx_1__1__32_top_grid_pin_22_;
wire [0:0] cbx_1__1__32_top_grid_pin_23_;
wire [0:0] cbx_1__1__32_top_grid_pin_24_;
wire [0:0] cbx_1__1__32_top_grid_pin_25_;
wire [0:0] cbx_1__1__32_top_grid_pin_26_;
wire [0:0] cbx_1__1__32_top_grid_pin_27_;
wire [0:0] cbx_1__1__32_top_grid_pin_28_;
wire [0:0] cbx_1__1__32_top_grid_pin_29_;
wire [0:0] cbx_1__1__32_top_grid_pin_30_;
wire [0:0] cbx_1__1__32_top_grid_pin_31_;
wire [0:0] cbx_1__1__33_ccff_tail;
wire [0:19] cbx_1__1__33_chanx_left_out;
wire [0:19] cbx_1__1__33_chanx_right_out;
wire [0:0] cbx_1__1__33_top_grid_pin_16_;
wire [0:0] cbx_1__1__33_top_grid_pin_17_;
wire [0:0] cbx_1__1__33_top_grid_pin_18_;
wire [0:0] cbx_1__1__33_top_grid_pin_19_;
wire [0:0] cbx_1__1__33_top_grid_pin_20_;
wire [0:0] cbx_1__1__33_top_grid_pin_21_;
wire [0:0] cbx_1__1__33_top_grid_pin_22_;
wire [0:0] cbx_1__1__33_top_grid_pin_23_;
wire [0:0] cbx_1__1__33_top_grid_pin_24_;
wire [0:0] cbx_1__1__33_top_grid_pin_25_;
wire [0:0] cbx_1__1__33_top_grid_pin_26_;
wire [0:0] cbx_1__1__33_top_grid_pin_27_;
wire [0:0] cbx_1__1__33_top_grid_pin_28_;
wire [0:0] cbx_1__1__33_top_grid_pin_29_;
wire [0:0] cbx_1__1__33_top_grid_pin_30_;
wire [0:0] cbx_1__1__33_top_grid_pin_31_;
wire [0:0] cbx_1__1__34_ccff_tail;
wire [0:19] cbx_1__1__34_chanx_left_out;
wire [0:19] cbx_1__1__34_chanx_right_out;
wire [0:0] cbx_1__1__34_top_grid_pin_16_;
wire [0:0] cbx_1__1__34_top_grid_pin_17_;
wire [0:0] cbx_1__1__34_top_grid_pin_18_;
wire [0:0] cbx_1__1__34_top_grid_pin_19_;
wire [0:0] cbx_1__1__34_top_grid_pin_20_;
wire [0:0] cbx_1__1__34_top_grid_pin_21_;
wire [0:0] cbx_1__1__34_top_grid_pin_22_;
wire [0:0] cbx_1__1__34_top_grid_pin_23_;
wire [0:0] cbx_1__1__34_top_grid_pin_24_;
wire [0:0] cbx_1__1__34_top_grid_pin_25_;
wire [0:0] cbx_1__1__34_top_grid_pin_26_;
wire [0:0] cbx_1__1__34_top_grid_pin_27_;
wire [0:0] cbx_1__1__34_top_grid_pin_28_;
wire [0:0] cbx_1__1__34_top_grid_pin_29_;
wire [0:0] cbx_1__1__34_top_grid_pin_30_;
wire [0:0] cbx_1__1__34_top_grid_pin_31_;
wire [0:0] cbx_1__1__35_ccff_tail;
wire [0:19] cbx_1__1__35_chanx_left_out;
wire [0:19] cbx_1__1__35_chanx_right_out;
wire [0:0] cbx_1__1__35_top_grid_pin_16_;
wire [0:0] cbx_1__1__35_top_grid_pin_17_;
wire [0:0] cbx_1__1__35_top_grid_pin_18_;
wire [0:0] cbx_1__1__35_top_grid_pin_19_;
wire [0:0] cbx_1__1__35_top_grid_pin_20_;
wire [0:0] cbx_1__1__35_top_grid_pin_21_;
wire [0:0] cbx_1__1__35_top_grid_pin_22_;
wire [0:0] cbx_1__1__35_top_grid_pin_23_;
wire [0:0] cbx_1__1__35_top_grid_pin_24_;
wire [0:0] cbx_1__1__35_top_grid_pin_25_;
wire [0:0] cbx_1__1__35_top_grid_pin_26_;
wire [0:0] cbx_1__1__35_top_grid_pin_27_;
wire [0:0] cbx_1__1__35_top_grid_pin_28_;
wire [0:0] cbx_1__1__35_top_grid_pin_29_;
wire [0:0] cbx_1__1__35_top_grid_pin_30_;
wire [0:0] cbx_1__1__35_top_grid_pin_31_;
wire [0:0] cbx_1__1__36_ccff_tail;
wire [0:19] cbx_1__1__36_chanx_left_out;
wire [0:19] cbx_1__1__36_chanx_right_out;
wire [0:0] cbx_1__1__36_top_grid_pin_16_;
wire [0:0] cbx_1__1__36_top_grid_pin_17_;
wire [0:0] cbx_1__1__36_top_grid_pin_18_;
wire [0:0] cbx_1__1__36_top_grid_pin_19_;
wire [0:0] cbx_1__1__36_top_grid_pin_20_;
wire [0:0] cbx_1__1__36_top_grid_pin_21_;
wire [0:0] cbx_1__1__36_top_grid_pin_22_;
wire [0:0] cbx_1__1__36_top_grid_pin_23_;
wire [0:0] cbx_1__1__36_top_grid_pin_24_;
wire [0:0] cbx_1__1__36_top_grid_pin_25_;
wire [0:0] cbx_1__1__36_top_grid_pin_26_;
wire [0:0] cbx_1__1__36_top_grid_pin_27_;
wire [0:0] cbx_1__1__36_top_grid_pin_28_;
wire [0:0] cbx_1__1__36_top_grid_pin_29_;
wire [0:0] cbx_1__1__36_top_grid_pin_30_;
wire [0:0] cbx_1__1__36_top_grid_pin_31_;
wire [0:0] cbx_1__1__37_ccff_tail;
wire [0:19] cbx_1__1__37_chanx_left_out;
wire [0:19] cbx_1__1__37_chanx_right_out;
wire [0:0] cbx_1__1__37_top_grid_pin_16_;
wire [0:0] cbx_1__1__37_top_grid_pin_17_;
wire [0:0] cbx_1__1__37_top_grid_pin_18_;
wire [0:0] cbx_1__1__37_top_grid_pin_19_;
wire [0:0] cbx_1__1__37_top_grid_pin_20_;
wire [0:0] cbx_1__1__37_top_grid_pin_21_;
wire [0:0] cbx_1__1__37_top_grid_pin_22_;
wire [0:0] cbx_1__1__37_top_grid_pin_23_;
wire [0:0] cbx_1__1__37_top_grid_pin_24_;
wire [0:0] cbx_1__1__37_top_grid_pin_25_;
wire [0:0] cbx_1__1__37_top_grid_pin_26_;
wire [0:0] cbx_1__1__37_top_grid_pin_27_;
wire [0:0] cbx_1__1__37_top_grid_pin_28_;
wire [0:0] cbx_1__1__37_top_grid_pin_29_;
wire [0:0] cbx_1__1__37_top_grid_pin_30_;
wire [0:0] cbx_1__1__37_top_grid_pin_31_;
wire [0:0] cbx_1__1__38_ccff_tail;
wire [0:19] cbx_1__1__38_chanx_left_out;
wire [0:19] cbx_1__1__38_chanx_right_out;
wire [0:0] cbx_1__1__38_top_grid_pin_16_;
wire [0:0] cbx_1__1__38_top_grid_pin_17_;
wire [0:0] cbx_1__1__38_top_grid_pin_18_;
wire [0:0] cbx_1__1__38_top_grid_pin_19_;
wire [0:0] cbx_1__1__38_top_grid_pin_20_;
wire [0:0] cbx_1__1__38_top_grid_pin_21_;
wire [0:0] cbx_1__1__38_top_grid_pin_22_;
wire [0:0] cbx_1__1__38_top_grid_pin_23_;
wire [0:0] cbx_1__1__38_top_grid_pin_24_;
wire [0:0] cbx_1__1__38_top_grid_pin_25_;
wire [0:0] cbx_1__1__38_top_grid_pin_26_;
wire [0:0] cbx_1__1__38_top_grid_pin_27_;
wire [0:0] cbx_1__1__38_top_grid_pin_28_;
wire [0:0] cbx_1__1__38_top_grid_pin_29_;
wire [0:0] cbx_1__1__38_top_grid_pin_30_;
wire [0:0] cbx_1__1__38_top_grid_pin_31_;
wire [0:0] cbx_1__1__39_ccff_tail;
wire [0:19] cbx_1__1__39_chanx_left_out;
wire [0:19] cbx_1__1__39_chanx_right_out;
wire [0:0] cbx_1__1__39_top_grid_pin_16_;
wire [0:0] cbx_1__1__39_top_grid_pin_17_;
wire [0:0] cbx_1__1__39_top_grid_pin_18_;
wire [0:0] cbx_1__1__39_top_grid_pin_19_;
wire [0:0] cbx_1__1__39_top_grid_pin_20_;
wire [0:0] cbx_1__1__39_top_grid_pin_21_;
wire [0:0] cbx_1__1__39_top_grid_pin_22_;
wire [0:0] cbx_1__1__39_top_grid_pin_23_;
wire [0:0] cbx_1__1__39_top_grid_pin_24_;
wire [0:0] cbx_1__1__39_top_grid_pin_25_;
wire [0:0] cbx_1__1__39_top_grid_pin_26_;
wire [0:0] cbx_1__1__39_top_grid_pin_27_;
wire [0:0] cbx_1__1__39_top_grid_pin_28_;
wire [0:0] cbx_1__1__39_top_grid_pin_29_;
wire [0:0] cbx_1__1__39_top_grid_pin_30_;
wire [0:0] cbx_1__1__39_top_grid_pin_31_;
wire [0:0] cbx_1__1__3_ccff_tail;
wire [0:19] cbx_1__1__3_chanx_left_out;
wire [0:19] cbx_1__1__3_chanx_right_out;
wire [0:0] cbx_1__1__3_top_grid_pin_16_;
wire [0:0] cbx_1__1__3_top_grid_pin_17_;
wire [0:0] cbx_1__1__3_top_grid_pin_18_;
wire [0:0] cbx_1__1__3_top_grid_pin_19_;
wire [0:0] cbx_1__1__3_top_grid_pin_20_;
wire [0:0] cbx_1__1__3_top_grid_pin_21_;
wire [0:0] cbx_1__1__3_top_grid_pin_22_;
wire [0:0] cbx_1__1__3_top_grid_pin_23_;
wire [0:0] cbx_1__1__3_top_grid_pin_24_;
wire [0:0] cbx_1__1__3_top_grid_pin_25_;
wire [0:0] cbx_1__1__3_top_grid_pin_26_;
wire [0:0] cbx_1__1__3_top_grid_pin_27_;
wire [0:0] cbx_1__1__3_top_grid_pin_28_;
wire [0:0] cbx_1__1__3_top_grid_pin_29_;
wire [0:0] cbx_1__1__3_top_grid_pin_30_;
wire [0:0] cbx_1__1__3_top_grid_pin_31_;
wire [0:0] cbx_1__1__40_ccff_tail;
wire [0:19] cbx_1__1__40_chanx_left_out;
wire [0:19] cbx_1__1__40_chanx_right_out;
wire [0:0] cbx_1__1__40_top_grid_pin_16_;
wire [0:0] cbx_1__1__40_top_grid_pin_17_;
wire [0:0] cbx_1__1__40_top_grid_pin_18_;
wire [0:0] cbx_1__1__40_top_grid_pin_19_;
wire [0:0] cbx_1__1__40_top_grid_pin_20_;
wire [0:0] cbx_1__1__40_top_grid_pin_21_;
wire [0:0] cbx_1__1__40_top_grid_pin_22_;
wire [0:0] cbx_1__1__40_top_grid_pin_23_;
wire [0:0] cbx_1__1__40_top_grid_pin_24_;
wire [0:0] cbx_1__1__40_top_grid_pin_25_;
wire [0:0] cbx_1__1__40_top_grid_pin_26_;
wire [0:0] cbx_1__1__40_top_grid_pin_27_;
wire [0:0] cbx_1__1__40_top_grid_pin_28_;
wire [0:0] cbx_1__1__40_top_grid_pin_29_;
wire [0:0] cbx_1__1__40_top_grid_pin_30_;
wire [0:0] cbx_1__1__40_top_grid_pin_31_;
wire [0:0] cbx_1__1__41_ccff_tail;
wire [0:19] cbx_1__1__41_chanx_left_out;
wire [0:19] cbx_1__1__41_chanx_right_out;
wire [0:0] cbx_1__1__41_top_grid_pin_16_;
wire [0:0] cbx_1__1__41_top_grid_pin_17_;
wire [0:0] cbx_1__1__41_top_grid_pin_18_;
wire [0:0] cbx_1__1__41_top_grid_pin_19_;
wire [0:0] cbx_1__1__41_top_grid_pin_20_;
wire [0:0] cbx_1__1__41_top_grid_pin_21_;
wire [0:0] cbx_1__1__41_top_grid_pin_22_;
wire [0:0] cbx_1__1__41_top_grid_pin_23_;
wire [0:0] cbx_1__1__41_top_grid_pin_24_;
wire [0:0] cbx_1__1__41_top_grid_pin_25_;
wire [0:0] cbx_1__1__41_top_grid_pin_26_;
wire [0:0] cbx_1__1__41_top_grid_pin_27_;
wire [0:0] cbx_1__1__41_top_grid_pin_28_;
wire [0:0] cbx_1__1__41_top_grid_pin_29_;
wire [0:0] cbx_1__1__41_top_grid_pin_30_;
wire [0:0] cbx_1__1__41_top_grid_pin_31_;
wire [0:0] cbx_1__1__42_ccff_tail;
wire [0:19] cbx_1__1__42_chanx_left_out;
wire [0:19] cbx_1__1__42_chanx_right_out;
wire [0:0] cbx_1__1__42_top_grid_pin_16_;
wire [0:0] cbx_1__1__42_top_grid_pin_17_;
wire [0:0] cbx_1__1__42_top_grid_pin_18_;
wire [0:0] cbx_1__1__42_top_grid_pin_19_;
wire [0:0] cbx_1__1__42_top_grid_pin_20_;
wire [0:0] cbx_1__1__42_top_grid_pin_21_;
wire [0:0] cbx_1__1__42_top_grid_pin_22_;
wire [0:0] cbx_1__1__42_top_grid_pin_23_;
wire [0:0] cbx_1__1__42_top_grid_pin_24_;
wire [0:0] cbx_1__1__42_top_grid_pin_25_;
wire [0:0] cbx_1__1__42_top_grid_pin_26_;
wire [0:0] cbx_1__1__42_top_grid_pin_27_;
wire [0:0] cbx_1__1__42_top_grid_pin_28_;
wire [0:0] cbx_1__1__42_top_grid_pin_29_;
wire [0:0] cbx_1__1__42_top_grid_pin_30_;
wire [0:0] cbx_1__1__42_top_grid_pin_31_;
wire [0:0] cbx_1__1__43_ccff_tail;
wire [0:19] cbx_1__1__43_chanx_left_out;
wire [0:19] cbx_1__1__43_chanx_right_out;
wire [0:0] cbx_1__1__43_top_grid_pin_16_;
wire [0:0] cbx_1__1__43_top_grid_pin_17_;
wire [0:0] cbx_1__1__43_top_grid_pin_18_;
wire [0:0] cbx_1__1__43_top_grid_pin_19_;
wire [0:0] cbx_1__1__43_top_grid_pin_20_;
wire [0:0] cbx_1__1__43_top_grid_pin_21_;
wire [0:0] cbx_1__1__43_top_grid_pin_22_;
wire [0:0] cbx_1__1__43_top_grid_pin_23_;
wire [0:0] cbx_1__1__43_top_grid_pin_24_;
wire [0:0] cbx_1__1__43_top_grid_pin_25_;
wire [0:0] cbx_1__1__43_top_grid_pin_26_;
wire [0:0] cbx_1__1__43_top_grid_pin_27_;
wire [0:0] cbx_1__1__43_top_grid_pin_28_;
wire [0:0] cbx_1__1__43_top_grid_pin_29_;
wire [0:0] cbx_1__1__43_top_grid_pin_30_;
wire [0:0] cbx_1__1__43_top_grid_pin_31_;
wire [0:0] cbx_1__1__44_ccff_tail;
wire [0:19] cbx_1__1__44_chanx_left_out;
wire [0:19] cbx_1__1__44_chanx_right_out;
wire [0:0] cbx_1__1__44_top_grid_pin_16_;
wire [0:0] cbx_1__1__44_top_grid_pin_17_;
wire [0:0] cbx_1__1__44_top_grid_pin_18_;
wire [0:0] cbx_1__1__44_top_grid_pin_19_;
wire [0:0] cbx_1__1__44_top_grid_pin_20_;
wire [0:0] cbx_1__1__44_top_grid_pin_21_;
wire [0:0] cbx_1__1__44_top_grid_pin_22_;
wire [0:0] cbx_1__1__44_top_grid_pin_23_;
wire [0:0] cbx_1__1__44_top_grid_pin_24_;
wire [0:0] cbx_1__1__44_top_grid_pin_25_;
wire [0:0] cbx_1__1__44_top_grid_pin_26_;
wire [0:0] cbx_1__1__44_top_grid_pin_27_;
wire [0:0] cbx_1__1__44_top_grid_pin_28_;
wire [0:0] cbx_1__1__44_top_grid_pin_29_;
wire [0:0] cbx_1__1__44_top_grid_pin_30_;
wire [0:0] cbx_1__1__44_top_grid_pin_31_;
wire [0:0] cbx_1__1__45_ccff_tail;
wire [0:19] cbx_1__1__45_chanx_left_out;
wire [0:19] cbx_1__1__45_chanx_right_out;
wire [0:0] cbx_1__1__45_top_grid_pin_16_;
wire [0:0] cbx_1__1__45_top_grid_pin_17_;
wire [0:0] cbx_1__1__45_top_grid_pin_18_;
wire [0:0] cbx_1__1__45_top_grid_pin_19_;
wire [0:0] cbx_1__1__45_top_grid_pin_20_;
wire [0:0] cbx_1__1__45_top_grid_pin_21_;
wire [0:0] cbx_1__1__45_top_grid_pin_22_;
wire [0:0] cbx_1__1__45_top_grid_pin_23_;
wire [0:0] cbx_1__1__45_top_grid_pin_24_;
wire [0:0] cbx_1__1__45_top_grid_pin_25_;
wire [0:0] cbx_1__1__45_top_grid_pin_26_;
wire [0:0] cbx_1__1__45_top_grid_pin_27_;
wire [0:0] cbx_1__1__45_top_grid_pin_28_;
wire [0:0] cbx_1__1__45_top_grid_pin_29_;
wire [0:0] cbx_1__1__45_top_grid_pin_30_;
wire [0:0] cbx_1__1__45_top_grid_pin_31_;
wire [0:0] cbx_1__1__46_ccff_tail;
wire [0:19] cbx_1__1__46_chanx_left_out;
wire [0:19] cbx_1__1__46_chanx_right_out;
wire [0:0] cbx_1__1__46_top_grid_pin_16_;
wire [0:0] cbx_1__1__46_top_grid_pin_17_;
wire [0:0] cbx_1__1__46_top_grid_pin_18_;
wire [0:0] cbx_1__1__46_top_grid_pin_19_;
wire [0:0] cbx_1__1__46_top_grid_pin_20_;
wire [0:0] cbx_1__1__46_top_grid_pin_21_;
wire [0:0] cbx_1__1__46_top_grid_pin_22_;
wire [0:0] cbx_1__1__46_top_grid_pin_23_;
wire [0:0] cbx_1__1__46_top_grid_pin_24_;
wire [0:0] cbx_1__1__46_top_grid_pin_25_;
wire [0:0] cbx_1__1__46_top_grid_pin_26_;
wire [0:0] cbx_1__1__46_top_grid_pin_27_;
wire [0:0] cbx_1__1__46_top_grid_pin_28_;
wire [0:0] cbx_1__1__46_top_grid_pin_29_;
wire [0:0] cbx_1__1__46_top_grid_pin_30_;
wire [0:0] cbx_1__1__46_top_grid_pin_31_;
wire [0:0] cbx_1__1__47_ccff_tail;
wire [0:19] cbx_1__1__47_chanx_left_out;
wire [0:19] cbx_1__1__47_chanx_right_out;
wire [0:0] cbx_1__1__47_top_grid_pin_16_;
wire [0:0] cbx_1__1__47_top_grid_pin_17_;
wire [0:0] cbx_1__1__47_top_grid_pin_18_;
wire [0:0] cbx_1__1__47_top_grid_pin_19_;
wire [0:0] cbx_1__1__47_top_grid_pin_20_;
wire [0:0] cbx_1__1__47_top_grid_pin_21_;
wire [0:0] cbx_1__1__47_top_grid_pin_22_;
wire [0:0] cbx_1__1__47_top_grid_pin_23_;
wire [0:0] cbx_1__1__47_top_grid_pin_24_;
wire [0:0] cbx_1__1__47_top_grid_pin_25_;
wire [0:0] cbx_1__1__47_top_grid_pin_26_;
wire [0:0] cbx_1__1__47_top_grid_pin_27_;
wire [0:0] cbx_1__1__47_top_grid_pin_28_;
wire [0:0] cbx_1__1__47_top_grid_pin_29_;
wire [0:0] cbx_1__1__47_top_grid_pin_30_;
wire [0:0] cbx_1__1__47_top_grid_pin_31_;
wire [0:0] cbx_1__1__48_ccff_tail;
wire [0:19] cbx_1__1__48_chanx_left_out;
wire [0:19] cbx_1__1__48_chanx_right_out;
wire [0:0] cbx_1__1__48_top_grid_pin_16_;
wire [0:0] cbx_1__1__48_top_grid_pin_17_;
wire [0:0] cbx_1__1__48_top_grid_pin_18_;
wire [0:0] cbx_1__1__48_top_grid_pin_19_;
wire [0:0] cbx_1__1__48_top_grid_pin_20_;
wire [0:0] cbx_1__1__48_top_grid_pin_21_;
wire [0:0] cbx_1__1__48_top_grid_pin_22_;
wire [0:0] cbx_1__1__48_top_grid_pin_23_;
wire [0:0] cbx_1__1__48_top_grid_pin_24_;
wire [0:0] cbx_1__1__48_top_grid_pin_25_;
wire [0:0] cbx_1__1__48_top_grid_pin_26_;
wire [0:0] cbx_1__1__48_top_grid_pin_27_;
wire [0:0] cbx_1__1__48_top_grid_pin_28_;
wire [0:0] cbx_1__1__48_top_grid_pin_29_;
wire [0:0] cbx_1__1__48_top_grid_pin_30_;
wire [0:0] cbx_1__1__48_top_grid_pin_31_;
wire [0:0] cbx_1__1__49_ccff_tail;
wire [0:19] cbx_1__1__49_chanx_left_out;
wire [0:19] cbx_1__1__49_chanx_right_out;
wire [0:0] cbx_1__1__49_top_grid_pin_16_;
wire [0:0] cbx_1__1__49_top_grid_pin_17_;
wire [0:0] cbx_1__1__49_top_grid_pin_18_;
wire [0:0] cbx_1__1__49_top_grid_pin_19_;
wire [0:0] cbx_1__1__49_top_grid_pin_20_;
wire [0:0] cbx_1__1__49_top_grid_pin_21_;
wire [0:0] cbx_1__1__49_top_grid_pin_22_;
wire [0:0] cbx_1__1__49_top_grid_pin_23_;
wire [0:0] cbx_1__1__49_top_grid_pin_24_;
wire [0:0] cbx_1__1__49_top_grid_pin_25_;
wire [0:0] cbx_1__1__49_top_grid_pin_26_;
wire [0:0] cbx_1__1__49_top_grid_pin_27_;
wire [0:0] cbx_1__1__49_top_grid_pin_28_;
wire [0:0] cbx_1__1__49_top_grid_pin_29_;
wire [0:0] cbx_1__1__49_top_grid_pin_30_;
wire [0:0] cbx_1__1__49_top_grid_pin_31_;
wire [0:0] cbx_1__1__4_ccff_tail;
wire [0:19] cbx_1__1__4_chanx_left_out;
wire [0:19] cbx_1__1__4_chanx_right_out;
wire [0:0] cbx_1__1__4_top_grid_pin_16_;
wire [0:0] cbx_1__1__4_top_grid_pin_17_;
wire [0:0] cbx_1__1__4_top_grid_pin_18_;
wire [0:0] cbx_1__1__4_top_grid_pin_19_;
wire [0:0] cbx_1__1__4_top_grid_pin_20_;
wire [0:0] cbx_1__1__4_top_grid_pin_21_;
wire [0:0] cbx_1__1__4_top_grid_pin_22_;
wire [0:0] cbx_1__1__4_top_grid_pin_23_;
wire [0:0] cbx_1__1__4_top_grid_pin_24_;
wire [0:0] cbx_1__1__4_top_grid_pin_25_;
wire [0:0] cbx_1__1__4_top_grid_pin_26_;
wire [0:0] cbx_1__1__4_top_grid_pin_27_;
wire [0:0] cbx_1__1__4_top_grid_pin_28_;
wire [0:0] cbx_1__1__4_top_grid_pin_29_;
wire [0:0] cbx_1__1__4_top_grid_pin_30_;
wire [0:0] cbx_1__1__4_top_grid_pin_31_;
wire [0:0] cbx_1__1__50_ccff_tail;
wire [0:19] cbx_1__1__50_chanx_left_out;
wire [0:19] cbx_1__1__50_chanx_right_out;
wire [0:0] cbx_1__1__50_top_grid_pin_16_;
wire [0:0] cbx_1__1__50_top_grid_pin_17_;
wire [0:0] cbx_1__1__50_top_grid_pin_18_;
wire [0:0] cbx_1__1__50_top_grid_pin_19_;
wire [0:0] cbx_1__1__50_top_grid_pin_20_;
wire [0:0] cbx_1__1__50_top_grid_pin_21_;
wire [0:0] cbx_1__1__50_top_grid_pin_22_;
wire [0:0] cbx_1__1__50_top_grid_pin_23_;
wire [0:0] cbx_1__1__50_top_grid_pin_24_;
wire [0:0] cbx_1__1__50_top_grid_pin_25_;
wire [0:0] cbx_1__1__50_top_grid_pin_26_;
wire [0:0] cbx_1__1__50_top_grid_pin_27_;
wire [0:0] cbx_1__1__50_top_grid_pin_28_;
wire [0:0] cbx_1__1__50_top_grid_pin_29_;
wire [0:0] cbx_1__1__50_top_grid_pin_30_;
wire [0:0] cbx_1__1__50_top_grid_pin_31_;
wire [0:0] cbx_1__1__51_ccff_tail;
wire [0:19] cbx_1__1__51_chanx_left_out;
wire [0:19] cbx_1__1__51_chanx_right_out;
wire [0:0] cbx_1__1__51_top_grid_pin_16_;
wire [0:0] cbx_1__1__51_top_grid_pin_17_;
wire [0:0] cbx_1__1__51_top_grid_pin_18_;
wire [0:0] cbx_1__1__51_top_grid_pin_19_;
wire [0:0] cbx_1__1__51_top_grid_pin_20_;
wire [0:0] cbx_1__1__51_top_grid_pin_21_;
wire [0:0] cbx_1__1__51_top_grid_pin_22_;
wire [0:0] cbx_1__1__51_top_grid_pin_23_;
wire [0:0] cbx_1__1__51_top_grid_pin_24_;
wire [0:0] cbx_1__1__51_top_grid_pin_25_;
wire [0:0] cbx_1__1__51_top_grid_pin_26_;
wire [0:0] cbx_1__1__51_top_grid_pin_27_;
wire [0:0] cbx_1__1__51_top_grid_pin_28_;
wire [0:0] cbx_1__1__51_top_grid_pin_29_;
wire [0:0] cbx_1__1__51_top_grid_pin_30_;
wire [0:0] cbx_1__1__51_top_grid_pin_31_;
wire [0:0] cbx_1__1__52_ccff_tail;
wire [0:19] cbx_1__1__52_chanx_left_out;
wire [0:19] cbx_1__1__52_chanx_right_out;
wire [0:0] cbx_1__1__52_top_grid_pin_16_;
wire [0:0] cbx_1__1__52_top_grid_pin_17_;
wire [0:0] cbx_1__1__52_top_grid_pin_18_;
wire [0:0] cbx_1__1__52_top_grid_pin_19_;
wire [0:0] cbx_1__1__52_top_grid_pin_20_;
wire [0:0] cbx_1__1__52_top_grid_pin_21_;
wire [0:0] cbx_1__1__52_top_grid_pin_22_;
wire [0:0] cbx_1__1__52_top_grid_pin_23_;
wire [0:0] cbx_1__1__52_top_grid_pin_24_;
wire [0:0] cbx_1__1__52_top_grid_pin_25_;
wire [0:0] cbx_1__1__52_top_grid_pin_26_;
wire [0:0] cbx_1__1__52_top_grid_pin_27_;
wire [0:0] cbx_1__1__52_top_grid_pin_28_;
wire [0:0] cbx_1__1__52_top_grid_pin_29_;
wire [0:0] cbx_1__1__52_top_grid_pin_30_;
wire [0:0] cbx_1__1__52_top_grid_pin_31_;
wire [0:0] cbx_1__1__53_ccff_tail;
wire [0:19] cbx_1__1__53_chanx_left_out;
wire [0:19] cbx_1__1__53_chanx_right_out;
wire [0:0] cbx_1__1__53_top_grid_pin_16_;
wire [0:0] cbx_1__1__53_top_grid_pin_17_;
wire [0:0] cbx_1__1__53_top_grid_pin_18_;
wire [0:0] cbx_1__1__53_top_grid_pin_19_;
wire [0:0] cbx_1__1__53_top_grid_pin_20_;
wire [0:0] cbx_1__1__53_top_grid_pin_21_;
wire [0:0] cbx_1__1__53_top_grid_pin_22_;
wire [0:0] cbx_1__1__53_top_grid_pin_23_;
wire [0:0] cbx_1__1__53_top_grid_pin_24_;
wire [0:0] cbx_1__1__53_top_grid_pin_25_;
wire [0:0] cbx_1__1__53_top_grid_pin_26_;
wire [0:0] cbx_1__1__53_top_grid_pin_27_;
wire [0:0] cbx_1__1__53_top_grid_pin_28_;
wire [0:0] cbx_1__1__53_top_grid_pin_29_;
wire [0:0] cbx_1__1__53_top_grid_pin_30_;
wire [0:0] cbx_1__1__53_top_grid_pin_31_;
wire [0:0] cbx_1__1__54_ccff_tail;
wire [0:19] cbx_1__1__54_chanx_left_out;
wire [0:19] cbx_1__1__54_chanx_right_out;
wire [0:0] cbx_1__1__54_top_grid_pin_16_;
wire [0:0] cbx_1__1__54_top_grid_pin_17_;
wire [0:0] cbx_1__1__54_top_grid_pin_18_;
wire [0:0] cbx_1__1__54_top_grid_pin_19_;
wire [0:0] cbx_1__1__54_top_grid_pin_20_;
wire [0:0] cbx_1__1__54_top_grid_pin_21_;
wire [0:0] cbx_1__1__54_top_grid_pin_22_;
wire [0:0] cbx_1__1__54_top_grid_pin_23_;
wire [0:0] cbx_1__1__54_top_grid_pin_24_;
wire [0:0] cbx_1__1__54_top_grid_pin_25_;
wire [0:0] cbx_1__1__54_top_grid_pin_26_;
wire [0:0] cbx_1__1__54_top_grid_pin_27_;
wire [0:0] cbx_1__1__54_top_grid_pin_28_;
wire [0:0] cbx_1__1__54_top_grid_pin_29_;
wire [0:0] cbx_1__1__54_top_grid_pin_30_;
wire [0:0] cbx_1__1__54_top_grid_pin_31_;
wire [0:0] cbx_1__1__55_ccff_tail;
wire [0:19] cbx_1__1__55_chanx_left_out;
wire [0:19] cbx_1__1__55_chanx_right_out;
wire [0:0] cbx_1__1__55_top_grid_pin_16_;
wire [0:0] cbx_1__1__55_top_grid_pin_17_;
wire [0:0] cbx_1__1__55_top_grid_pin_18_;
wire [0:0] cbx_1__1__55_top_grid_pin_19_;
wire [0:0] cbx_1__1__55_top_grid_pin_20_;
wire [0:0] cbx_1__1__55_top_grid_pin_21_;
wire [0:0] cbx_1__1__55_top_grid_pin_22_;
wire [0:0] cbx_1__1__55_top_grid_pin_23_;
wire [0:0] cbx_1__1__55_top_grid_pin_24_;
wire [0:0] cbx_1__1__55_top_grid_pin_25_;
wire [0:0] cbx_1__1__55_top_grid_pin_26_;
wire [0:0] cbx_1__1__55_top_grid_pin_27_;
wire [0:0] cbx_1__1__55_top_grid_pin_28_;
wire [0:0] cbx_1__1__55_top_grid_pin_29_;
wire [0:0] cbx_1__1__55_top_grid_pin_30_;
wire [0:0] cbx_1__1__55_top_grid_pin_31_;
wire [0:0] cbx_1__1__56_ccff_tail;
wire [0:19] cbx_1__1__56_chanx_left_out;
wire [0:19] cbx_1__1__56_chanx_right_out;
wire [0:0] cbx_1__1__56_top_grid_pin_16_;
wire [0:0] cbx_1__1__56_top_grid_pin_17_;
wire [0:0] cbx_1__1__56_top_grid_pin_18_;
wire [0:0] cbx_1__1__56_top_grid_pin_19_;
wire [0:0] cbx_1__1__56_top_grid_pin_20_;
wire [0:0] cbx_1__1__56_top_grid_pin_21_;
wire [0:0] cbx_1__1__56_top_grid_pin_22_;
wire [0:0] cbx_1__1__56_top_grid_pin_23_;
wire [0:0] cbx_1__1__56_top_grid_pin_24_;
wire [0:0] cbx_1__1__56_top_grid_pin_25_;
wire [0:0] cbx_1__1__56_top_grid_pin_26_;
wire [0:0] cbx_1__1__56_top_grid_pin_27_;
wire [0:0] cbx_1__1__56_top_grid_pin_28_;
wire [0:0] cbx_1__1__56_top_grid_pin_29_;
wire [0:0] cbx_1__1__56_top_grid_pin_30_;
wire [0:0] cbx_1__1__56_top_grid_pin_31_;
wire [0:0] cbx_1__1__57_ccff_tail;
wire [0:19] cbx_1__1__57_chanx_left_out;
wire [0:19] cbx_1__1__57_chanx_right_out;
wire [0:0] cbx_1__1__57_top_grid_pin_16_;
wire [0:0] cbx_1__1__57_top_grid_pin_17_;
wire [0:0] cbx_1__1__57_top_grid_pin_18_;
wire [0:0] cbx_1__1__57_top_grid_pin_19_;
wire [0:0] cbx_1__1__57_top_grid_pin_20_;
wire [0:0] cbx_1__1__57_top_grid_pin_21_;
wire [0:0] cbx_1__1__57_top_grid_pin_22_;
wire [0:0] cbx_1__1__57_top_grid_pin_23_;
wire [0:0] cbx_1__1__57_top_grid_pin_24_;
wire [0:0] cbx_1__1__57_top_grid_pin_25_;
wire [0:0] cbx_1__1__57_top_grid_pin_26_;
wire [0:0] cbx_1__1__57_top_grid_pin_27_;
wire [0:0] cbx_1__1__57_top_grid_pin_28_;
wire [0:0] cbx_1__1__57_top_grid_pin_29_;
wire [0:0] cbx_1__1__57_top_grid_pin_30_;
wire [0:0] cbx_1__1__57_top_grid_pin_31_;
wire [0:0] cbx_1__1__58_ccff_tail;
wire [0:19] cbx_1__1__58_chanx_left_out;
wire [0:19] cbx_1__1__58_chanx_right_out;
wire [0:0] cbx_1__1__58_top_grid_pin_16_;
wire [0:0] cbx_1__1__58_top_grid_pin_17_;
wire [0:0] cbx_1__1__58_top_grid_pin_18_;
wire [0:0] cbx_1__1__58_top_grid_pin_19_;
wire [0:0] cbx_1__1__58_top_grid_pin_20_;
wire [0:0] cbx_1__1__58_top_grid_pin_21_;
wire [0:0] cbx_1__1__58_top_grid_pin_22_;
wire [0:0] cbx_1__1__58_top_grid_pin_23_;
wire [0:0] cbx_1__1__58_top_grid_pin_24_;
wire [0:0] cbx_1__1__58_top_grid_pin_25_;
wire [0:0] cbx_1__1__58_top_grid_pin_26_;
wire [0:0] cbx_1__1__58_top_grid_pin_27_;
wire [0:0] cbx_1__1__58_top_grid_pin_28_;
wire [0:0] cbx_1__1__58_top_grid_pin_29_;
wire [0:0] cbx_1__1__58_top_grid_pin_30_;
wire [0:0] cbx_1__1__58_top_grid_pin_31_;
wire [0:0] cbx_1__1__59_ccff_tail;
wire [0:19] cbx_1__1__59_chanx_left_out;
wire [0:19] cbx_1__1__59_chanx_right_out;
wire [0:0] cbx_1__1__59_top_grid_pin_16_;
wire [0:0] cbx_1__1__59_top_grid_pin_17_;
wire [0:0] cbx_1__1__59_top_grid_pin_18_;
wire [0:0] cbx_1__1__59_top_grid_pin_19_;
wire [0:0] cbx_1__1__59_top_grid_pin_20_;
wire [0:0] cbx_1__1__59_top_grid_pin_21_;
wire [0:0] cbx_1__1__59_top_grid_pin_22_;
wire [0:0] cbx_1__1__59_top_grid_pin_23_;
wire [0:0] cbx_1__1__59_top_grid_pin_24_;
wire [0:0] cbx_1__1__59_top_grid_pin_25_;
wire [0:0] cbx_1__1__59_top_grid_pin_26_;
wire [0:0] cbx_1__1__59_top_grid_pin_27_;
wire [0:0] cbx_1__1__59_top_grid_pin_28_;
wire [0:0] cbx_1__1__59_top_grid_pin_29_;
wire [0:0] cbx_1__1__59_top_grid_pin_30_;
wire [0:0] cbx_1__1__59_top_grid_pin_31_;
wire [0:0] cbx_1__1__5_ccff_tail;
wire [0:19] cbx_1__1__5_chanx_left_out;
wire [0:19] cbx_1__1__5_chanx_right_out;
wire [0:0] cbx_1__1__5_top_grid_pin_16_;
wire [0:0] cbx_1__1__5_top_grid_pin_17_;
wire [0:0] cbx_1__1__5_top_grid_pin_18_;
wire [0:0] cbx_1__1__5_top_grid_pin_19_;
wire [0:0] cbx_1__1__5_top_grid_pin_20_;
wire [0:0] cbx_1__1__5_top_grid_pin_21_;
wire [0:0] cbx_1__1__5_top_grid_pin_22_;
wire [0:0] cbx_1__1__5_top_grid_pin_23_;
wire [0:0] cbx_1__1__5_top_grid_pin_24_;
wire [0:0] cbx_1__1__5_top_grid_pin_25_;
wire [0:0] cbx_1__1__5_top_grid_pin_26_;
wire [0:0] cbx_1__1__5_top_grid_pin_27_;
wire [0:0] cbx_1__1__5_top_grid_pin_28_;
wire [0:0] cbx_1__1__5_top_grid_pin_29_;
wire [0:0] cbx_1__1__5_top_grid_pin_30_;
wire [0:0] cbx_1__1__5_top_grid_pin_31_;
wire [0:0] cbx_1__1__60_ccff_tail;
wire [0:19] cbx_1__1__60_chanx_left_out;
wire [0:19] cbx_1__1__60_chanx_right_out;
wire [0:0] cbx_1__1__60_top_grid_pin_16_;
wire [0:0] cbx_1__1__60_top_grid_pin_17_;
wire [0:0] cbx_1__1__60_top_grid_pin_18_;
wire [0:0] cbx_1__1__60_top_grid_pin_19_;
wire [0:0] cbx_1__1__60_top_grid_pin_20_;
wire [0:0] cbx_1__1__60_top_grid_pin_21_;
wire [0:0] cbx_1__1__60_top_grid_pin_22_;
wire [0:0] cbx_1__1__60_top_grid_pin_23_;
wire [0:0] cbx_1__1__60_top_grid_pin_24_;
wire [0:0] cbx_1__1__60_top_grid_pin_25_;
wire [0:0] cbx_1__1__60_top_grid_pin_26_;
wire [0:0] cbx_1__1__60_top_grid_pin_27_;
wire [0:0] cbx_1__1__60_top_grid_pin_28_;
wire [0:0] cbx_1__1__60_top_grid_pin_29_;
wire [0:0] cbx_1__1__60_top_grid_pin_30_;
wire [0:0] cbx_1__1__60_top_grid_pin_31_;
wire [0:0] cbx_1__1__61_ccff_tail;
wire [0:19] cbx_1__1__61_chanx_left_out;
wire [0:19] cbx_1__1__61_chanx_right_out;
wire [0:0] cbx_1__1__61_top_grid_pin_16_;
wire [0:0] cbx_1__1__61_top_grid_pin_17_;
wire [0:0] cbx_1__1__61_top_grid_pin_18_;
wire [0:0] cbx_1__1__61_top_grid_pin_19_;
wire [0:0] cbx_1__1__61_top_grid_pin_20_;
wire [0:0] cbx_1__1__61_top_grid_pin_21_;
wire [0:0] cbx_1__1__61_top_grid_pin_22_;
wire [0:0] cbx_1__1__61_top_grid_pin_23_;
wire [0:0] cbx_1__1__61_top_grid_pin_24_;
wire [0:0] cbx_1__1__61_top_grid_pin_25_;
wire [0:0] cbx_1__1__61_top_grid_pin_26_;
wire [0:0] cbx_1__1__61_top_grid_pin_27_;
wire [0:0] cbx_1__1__61_top_grid_pin_28_;
wire [0:0] cbx_1__1__61_top_grid_pin_29_;
wire [0:0] cbx_1__1__61_top_grid_pin_30_;
wire [0:0] cbx_1__1__61_top_grid_pin_31_;
wire [0:0] cbx_1__1__62_ccff_tail;
wire [0:19] cbx_1__1__62_chanx_left_out;
wire [0:19] cbx_1__1__62_chanx_right_out;
wire [0:0] cbx_1__1__62_top_grid_pin_16_;
wire [0:0] cbx_1__1__62_top_grid_pin_17_;
wire [0:0] cbx_1__1__62_top_grid_pin_18_;
wire [0:0] cbx_1__1__62_top_grid_pin_19_;
wire [0:0] cbx_1__1__62_top_grid_pin_20_;
wire [0:0] cbx_1__1__62_top_grid_pin_21_;
wire [0:0] cbx_1__1__62_top_grid_pin_22_;
wire [0:0] cbx_1__1__62_top_grid_pin_23_;
wire [0:0] cbx_1__1__62_top_grid_pin_24_;
wire [0:0] cbx_1__1__62_top_grid_pin_25_;
wire [0:0] cbx_1__1__62_top_grid_pin_26_;
wire [0:0] cbx_1__1__62_top_grid_pin_27_;
wire [0:0] cbx_1__1__62_top_grid_pin_28_;
wire [0:0] cbx_1__1__62_top_grid_pin_29_;
wire [0:0] cbx_1__1__62_top_grid_pin_30_;
wire [0:0] cbx_1__1__62_top_grid_pin_31_;
wire [0:0] cbx_1__1__63_ccff_tail;
wire [0:19] cbx_1__1__63_chanx_left_out;
wire [0:19] cbx_1__1__63_chanx_right_out;
wire [0:0] cbx_1__1__63_top_grid_pin_16_;
wire [0:0] cbx_1__1__63_top_grid_pin_17_;
wire [0:0] cbx_1__1__63_top_grid_pin_18_;
wire [0:0] cbx_1__1__63_top_grid_pin_19_;
wire [0:0] cbx_1__1__63_top_grid_pin_20_;
wire [0:0] cbx_1__1__63_top_grid_pin_21_;
wire [0:0] cbx_1__1__63_top_grid_pin_22_;
wire [0:0] cbx_1__1__63_top_grid_pin_23_;
wire [0:0] cbx_1__1__63_top_grid_pin_24_;
wire [0:0] cbx_1__1__63_top_grid_pin_25_;
wire [0:0] cbx_1__1__63_top_grid_pin_26_;
wire [0:0] cbx_1__1__63_top_grid_pin_27_;
wire [0:0] cbx_1__1__63_top_grid_pin_28_;
wire [0:0] cbx_1__1__63_top_grid_pin_29_;
wire [0:0] cbx_1__1__63_top_grid_pin_30_;
wire [0:0] cbx_1__1__63_top_grid_pin_31_;
wire [0:0] cbx_1__1__64_ccff_tail;
wire [0:19] cbx_1__1__64_chanx_left_out;
wire [0:19] cbx_1__1__64_chanx_right_out;
wire [0:0] cbx_1__1__64_top_grid_pin_16_;
wire [0:0] cbx_1__1__64_top_grid_pin_17_;
wire [0:0] cbx_1__1__64_top_grid_pin_18_;
wire [0:0] cbx_1__1__64_top_grid_pin_19_;
wire [0:0] cbx_1__1__64_top_grid_pin_20_;
wire [0:0] cbx_1__1__64_top_grid_pin_21_;
wire [0:0] cbx_1__1__64_top_grid_pin_22_;
wire [0:0] cbx_1__1__64_top_grid_pin_23_;
wire [0:0] cbx_1__1__64_top_grid_pin_24_;
wire [0:0] cbx_1__1__64_top_grid_pin_25_;
wire [0:0] cbx_1__1__64_top_grid_pin_26_;
wire [0:0] cbx_1__1__64_top_grid_pin_27_;
wire [0:0] cbx_1__1__64_top_grid_pin_28_;
wire [0:0] cbx_1__1__64_top_grid_pin_29_;
wire [0:0] cbx_1__1__64_top_grid_pin_30_;
wire [0:0] cbx_1__1__64_top_grid_pin_31_;
wire [0:0] cbx_1__1__65_ccff_tail;
wire [0:19] cbx_1__1__65_chanx_left_out;
wire [0:19] cbx_1__1__65_chanx_right_out;
wire [0:0] cbx_1__1__65_top_grid_pin_16_;
wire [0:0] cbx_1__1__65_top_grid_pin_17_;
wire [0:0] cbx_1__1__65_top_grid_pin_18_;
wire [0:0] cbx_1__1__65_top_grid_pin_19_;
wire [0:0] cbx_1__1__65_top_grid_pin_20_;
wire [0:0] cbx_1__1__65_top_grid_pin_21_;
wire [0:0] cbx_1__1__65_top_grid_pin_22_;
wire [0:0] cbx_1__1__65_top_grid_pin_23_;
wire [0:0] cbx_1__1__65_top_grid_pin_24_;
wire [0:0] cbx_1__1__65_top_grid_pin_25_;
wire [0:0] cbx_1__1__65_top_grid_pin_26_;
wire [0:0] cbx_1__1__65_top_grid_pin_27_;
wire [0:0] cbx_1__1__65_top_grid_pin_28_;
wire [0:0] cbx_1__1__65_top_grid_pin_29_;
wire [0:0] cbx_1__1__65_top_grid_pin_30_;
wire [0:0] cbx_1__1__65_top_grid_pin_31_;
wire [0:0] cbx_1__1__66_ccff_tail;
wire [0:19] cbx_1__1__66_chanx_left_out;
wire [0:19] cbx_1__1__66_chanx_right_out;
wire [0:0] cbx_1__1__66_top_grid_pin_16_;
wire [0:0] cbx_1__1__66_top_grid_pin_17_;
wire [0:0] cbx_1__1__66_top_grid_pin_18_;
wire [0:0] cbx_1__1__66_top_grid_pin_19_;
wire [0:0] cbx_1__1__66_top_grid_pin_20_;
wire [0:0] cbx_1__1__66_top_grid_pin_21_;
wire [0:0] cbx_1__1__66_top_grid_pin_22_;
wire [0:0] cbx_1__1__66_top_grid_pin_23_;
wire [0:0] cbx_1__1__66_top_grid_pin_24_;
wire [0:0] cbx_1__1__66_top_grid_pin_25_;
wire [0:0] cbx_1__1__66_top_grid_pin_26_;
wire [0:0] cbx_1__1__66_top_grid_pin_27_;
wire [0:0] cbx_1__1__66_top_grid_pin_28_;
wire [0:0] cbx_1__1__66_top_grid_pin_29_;
wire [0:0] cbx_1__1__66_top_grid_pin_30_;
wire [0:0] cbx_1__1__66_top_grid_pin_31_;
wire [0:0] cbx_1__1__67_ccff_tail;
wire [0:19] cbx_1__1__67_chanx_left_out;
wire [0:19] cbx_1__1__67_chanx_right_out;
wire [0:0] cbx_1__1__67_top_grid_pin_16_;
wire [0:0] cbx_1__1__67_top_grid_pin_17_;
wire [0:0] cbx_1__1__67_top_grid_pin_18_;
wire [0:0] cbx_1__1__67_top_grid_pin_19_;
wire [0:0] cbx_1__1__67_top_grid_pin_20_;
wire [0:0] cbx_1__1__67_top_grid_pin_21_;
wire [0:0] cbx_1__1__67_top_grid_pin_22_;
wire [0:0] cbx_1__1__67_top_grid_pin_23_;
wire [0:0] cbx_1__1__67_top_grid_pin_24_;
wire [0:0] cbx_1__1__67_top_grid_pin_25_;
wire [0:0] cbx_1__1__67_top_grid_pin_26_;
wire [0:0] cbx_1__1__67_top_grid_pin_27_;
wire [0:0] cbx_1__1__67_top_grid_pin_28_;
wire [0:0] cbx_1__1__67_top_grid_pin_29_;
wire [0:0] cbx_1__1__67_top_grid_pin_30_;
wire [0:0] cbx_1__1__67_top_grid_pin_31_;
wire [0:0] cbx_1__1__68_ccff_tail;
wire [0:19] cbx_1__1__68_chanx_left_out;
wire [0:19] cbx_1__1__68_chanx_right_out;
wire [0:0] cbx_1__1__68_top_grid_pin_16_;
wire [0:0] cbx_1__1__68_top_grid_pin_17_;
wire [0:0] cbx_1__1__68_top_grid_pin_18_;
wire [0:0] cbx_1__1__68_top_grid_pin_19_;
wire [0:0] cbx_1__1__68_top_grid_pin_20_;
wire [0:0] cbx_1__1__68_top_grid_pin_21_;
wire [0:0] cbx_1__1__68_top_grid_pin_22_;
wire [0:0] cbx_1__1__68_top_grid_pin_23_;
wire [0:0] cbx_1__1__68_top_grid_pin_24_;
wire [0:0] cbx_1__1__68_top_grid_pin_25_;
wire [0:0] cbx_1__1__68_top_grid_pin_26_;
wire [0:0] cbx_1__1__68_top_grid_pin_27_;
wire [0:0] cbx_1__1__68_top_grid_pin_28_;
wire [0:0] cbx_1__1__68_top_grid_pin_29_;
wire [0:0] cbx_1__1__68_top_grid_pin_30_;
wire [0:0] cbx_1__1__68_top_grid_pin_31_;
wire [0:0] cbx_1__1__69_ccff_tail;
wire [0:19] cbx_1__1__69_chanx_left_out;
wire [0:19] cbx_1__1__69_chanx_right_out;
wire [0:0] cbx_1__1__69_top_grid_pin_16_;
wire [0:0] cbx_1__1__69_top_grid_pin_17_;
wire [0:0] cbx_1__1__69_top_grid_pin_18_;
wire [0:0] cbx_1__1__69_top_grid_pin_19_;
wire [0:0] cbx_1__1__69_top_grid_pin_20_;
wire [0:0] cbx_1__1__69_top_grid_pin_21_;
wire [0:0] cbx_1__1__69_top_grid_pin_22_;
wire [0:0] cbx_1__1__69_top_grid_pin_23_;
wire [0:0] cbx_1__1__69_top_grid_pin_24_;
wire [0:0] cbx_1__1__69_top_grid_pin_25_;
wire [0:0] cbx_1__1__69_top_grid_pin_26_;
wire [0:0] cbx_1__1__69_top_grid_pin_27_;
wire [0:0] cbx_1__1__69_top_grid_pin_28_;
wire [0:0] cbx_1__1__69_top_grid_pin_29_;
wire [0:0] cbx_1__1__69_top_grid_pin_30_;
wire [0:0] cbx_1__1__69_top_grid_pin_31_;
wire [0:0] cbx_1__1__6_ccff_tail;
wire [0:19] cbx_1__1__6_chanx_left_out;
wire [0:19] cbx_1__1__6_chanx_right_out;
wire [0:0] cbx_1__1__6_top_grid_pin_16_;
wire [0:0] cbx_1__1__6_top_grid_pin_17_;
wire [0:0] cbx_1__1__6_top_grid_pin_18_;
wire [0:0] cbx_1__1__6_top_grid_pin_19_;
wire [0:0] cbx_1__1__6_top_grid_pin_20_;
wire [0:0] cbx_1__1__6_top_grid_pin_21_;
wire [0:0] cbx_1__1__6_top_grid_pin_22_;
wire [0:0] cbx_1__1__6_top_grid_pin_23_;
wire [0:0] cbx_1__1__6_top_grid_pin_24_;
wire [0:0] cbx_1__1__6_top_grid_pin_25_;
wire [0:0] cbx_1__1__6_top_grid_pin_26_;
wire [0:0] cbx_1__1__6_top_grid_pin_27_;
wire [0:0] cbx_1__1__6_top_grid_pin_28_;
wire [0:0] cbx_1__1__6_top_grid_pin_29_;
wire [0:0] cbx_1__1__6_top_grid_pin_30_;
wire [0:0] cbx_1__1__6_top_grid_pin_31_;
wire [0:0] cbx_1__1__70_ccff_tail;
wire [0:19] cbx_1__1__70_chanx_left_out;
wire [0:19] cbx_1__1__70_chanx_right_out;
wire [0:0] cbx_1__1__70_top_grid_pin_16_;
wire [0:0] cbx_1__1__70_top_grid_pin_17_;
wire [0:0] cbx_1__1__70_top_grid_pin_18_;
wire [0:0] cbx_1__1__70_top_grid_pin_19_;
wire [0:0] cbx_1__1__70_top_grid_pin_20_;
wire [0:0] cbx_1__1__70_top_grid_pin_21_;
wire [0:0] cbx_1__1__70_top_grid_pin_22_;
wire [0:0] cbx_1__1__70_top_grid_pin_23_;
wire [0:0] cbx_1__1__70_top_grid_pin_24_;
wire [0:0] cbx_1__1__70_top_grid_pin_25_;
wire [0:0] cbx_1__1__70_top_grid_pin_26_;
wire [0:0] cbx_1__1__70_top_grid_pin_27_;
wire [0:0] cbx_1__1__70_top_grid_pin_28_;
wire [0:0] cbx_1__1__70_top_grid_pin_29_;
wire [0:0] cbx_1__1__70_top_grid_pin_30_;
wire [0:0] cbx_1__1__70_top_grid_pin_31_;
wire [0:0] cbx_1__1__71_ccff_tail;
wire [0:19] cbx_1__1__71_chanx_left_out;
wire [0:19] cbx_1__1__71_chanx_right_out;
wire [0:0] cbx_1__1__71_top_grid_pin_16_;
wire [0:0] cbx_1__1__71_top_grid_pin_17_;
wire [0:0] cbx_1__1__71_top_grid_pin_18_;
wire [0:0] cbx_1__1__71_top_grid_pin_19_;
wire [0:0] cbx_1__1__71_top_grid_pin_20_;
wire [0:0] cbx_1__1__71_top_grid_pin_21_;
wire [0:0] cbx_1__1__71_top_grid_pin_22_;
wire [0:0] cbx_1__1__71_top_grid_pin_23_;
wire [0:0] cbx_1__1__71_top_grid_pin_24_;
wire [0:0] cbx_1__1__71_top_grid_pin_25_;
wire [0:0] cbx_1__1__71_top_grid_pin_26_;
wire [0:0] cbx_1__1__71_top_grid_pin_27_;
wire [0:0] cbx_1__1__71_top_grid_pin_28_;
wire [0:0] cbx_1__1__71_top_grid_pin_29_;
wire [0:0] cbx_1__1__71_top_grid_pin_30_;
wire [0:0] cbx_1__1__71_top_grid_pin_31_;
wire [0:0] cbx_1__1__72_ccff_tail;
wire [0:19] cbx_1__1__72_chanx_left_out;
wire [0:19] cbx_1__1__72_chanx_right_out;
wire [0:0] cbx_1__1__72_top_grid_pin_16_;
wire [0:0] cbx_1__1__72_top_grid_pin_17_;
wire [0:0] cbx_1__1__72_top_grid_pin_18_;
wire [0:0] cbx_1__1__72_top_grid_pin_19_;
wire [0:0] cbx_1__1__72_top_grid_pin_20_;
wire [0:0] cbx_1__1__72_top_grid_pin_21_;
wire [0:0] cbx_1__1__72_top_grid_pin_22_;
wire [0:0] cbx_1__1__72_top_grid_pin_23_;
wire [0:0] cbx_1__1__72_top_grid_pin_24_;
wire [0:0] cbx_1__1__72_top_grid_pin_25_;
wire [0:0] cbx_1__1__72_top_grid_pin_26_;
wire [0:0] cbx_1__1__72_top_grid_pin_27_;
wire [0:0] cbx_1__1__72_top_grid_pin_28_;
wire [0:0] cbx_1__1__72_top_grid_pin_29_;
wire [0:0] cbx_1__1__72_top_grid_pin_30_;
wire [0:0] cbx_1__1__72_top_grid_pin_31_;
wire [0:0] cbx_1__1__73_ccff_tail;
wire [0:19] cbx_1__1__73_chanx_left_out;
wire [0:19] cbx_1__1__73_chanx_right_out;
wire [0:0] cbx_1__1__73_top_grid_pin_16_;
wire [0:0] cbx_1__1__73_top_grid_pin_17_;
wire [0:0] cbx_1__1__73_top_grid_pin_18_;
wire [0:0] cbx_1__1__73_top_grid_pin_19_;
wire [0:0] cbx_1__1__73_top_grid_pin_20_;
wire [0:0] cbx_1__1__73_top_grid_pin_21_;
wire [0:0] cbx_1__1__73_top_grid_pin_22_;
wire [0:0] cbx_1__1__73_top_grid_pin_23_;
wire [0:0] cbx_1__1__73_top_grid_pin_24_;
wire [0:0] cbx_1__1__73_top_grid_pin_25_;
wire [0:0] cbx_1__1__73_top_grid_pin_26_;
wire [0:0] cbx_1__1__73_top_grid_pin_27_;
wire [0:0] cbx_1__1__73_top_grid_pin_28_;
wire [0:0] cbx_1__1__73_top_grid_pin_29_;
wire [0:0] cbx_1__1__73_top_grid_pin_30_;
wire [0:0] cbx_1__1__73_top_grid_pin_31_;
wire [0:0] cbx_1__1__74_ccff_tail;
wire [0:19] cbx_1__1__74_chanx_left_out;
wire [0:19] cbx_1__1__74_chanx_right_out;
wire [0:0] cbx_1__1__74_top_grid_pin_16_;
wire [0:0] cbx_1__1__74_top_grid_pin_17_;
wire [0:0] cbx_1__1__74_top_grid_pin_18_;
wire [0:0] cbx_1__1__74_top_grid_pin_19_;
wire [0:0] cbx_1__1__74_top_grid_pin_20_;
wire [0:0] cbx_1__1__74_top_grid_pin_21_;
wire [0:0] cbx_1__1__74_top_grid_pin_22_;
wire [0:0] cbx_1__1__74_top_grid_pin_23_;
wire [0:0] cbx_1__1__74_top_grid_pin_24_;
wire [0:0] cbx_1__1__74_top_grid_pin_25_;
wire [0:0] cbx_1__1__74_top_grid_pin_26_;
wire [0:0] cbx_1__1__74_top_grid_pin_27_;
wire [0:0] cbx_1__1__74_top_grid_pin_28_;
wire [0:0] cbx_1__1__74_top_grid_pin_29_;
wire [0:0] cbx_1__1__74_top_grid_pin_30_;
wire [0:0] cbx_1__1__74_top_grid_pin_31_;
wire [0:0] cbx_1__1__75_ccff_tail;
wire [0:19] cbx_1__1__75_chanx_left_out;
wire [0:19] cbx_1__1__75_chanx_right_out;
wire [0:0] cbx_1__1__75_top_grid_pin_16_;
wire [0:0] cbx_1__1__75_top_grid_pin_17_;
wire [0:0] cbx_1__1__75_top_grid_pin_18_;
wire [0:0] cbx_1__1__75_top_grid_pin_19_;
wire [0:0] cbx_1__1__75_top_grid_pin_20_;
wire [0:0] cbx_1__1__75_top_grid_pin_21_;
wire [0:0] cbx_1__1__75_top_grid_pin_22_;
wire [0:0] cbx_1__1__75_top_grid_pin_23_;
wire [0:0] cbx_1__1__75_top_grid_pin_24_;
wire [0:0] cbx_1__1__75_top_grid_pin_25_;
wire [0:0] cbx_1__1__75_top_grid_pin_26_;
wire [0:0] cbx_1__1__75_top_grid_pin_27_;
wire [0:0] cbx_1__1__75_top_grid_pin_28_;
wire [0:0] cbx_1__1__75_top_grid_pin_29_;
wire [0:0] cbx_1__1__75_top_grid_pin_30_;
wire [0:0] cbx_1__1__75_top_grid_pin_31_;
wire [0:0] cbx_1__1__76_ccff_tail;
wire [0:19] cbx_1__1__76_chanx_left_out;
wire [0:19] cbx_1__1__76_chanx_right_out;
wire [0:0] cbx_1__1__76_top_grid_pin_16_;
wire [0:0] cbx_1__1__76_top_grid_pin_17_;
wire [0:0] cbx_1__1__76_top_grid_pin_18_;
wire [0:0] cbx_1__1__76_top_grid_pin_19_;
wire [0:0] cbx_1__1__76_top_grid_pin_20_;
wire [0:0] cbx_1__1__76_top_grid_pin_21_;
wire [0:0] cbx_1__1__76_top_grid_pin_22_;
wire [0:0] cbx_1__1__76_top_grid_pin_23_;
wire [0:0] cbx_1__1__76_top_grid_pin_24_;
wire [0:0] cbx_1__1__76_top_grid_pin_25_;
wire [0:0] cbx_1__1__76_top_grid_pin_26_;
wire [0:0] cbx_1__1__76_top_grid_pin_27_;
wire [0:0] cbx_1__1__76_top_grid_pin_28_;
wire [0:0] cbx_1__1__76_top_grid_pin_29_;
wire [0:0] cbx_1__1__76_top_grid_pin_30_;
wire [0:0] cbx_1__1__76_top_grid_pin_31_;
wire [0:0] cbx_1__1__77_ccff_tail;
wire [0:19] cbx_1__1__77_chanx_left_out;
wire [0:19] cbx_1__1__77_chanx_right_out;
wire [0:0] cbx_1__1__77_top_grid_pin_16_;
wire [0:0] cbx_1__1__77_top_grid_pin_17_;
wire [0:0] cbx_1__1__77_top_grid_pin_18_;
wire [0:0] cbx_1__1__77_top_grid_pin_19_;
wire [0:0] cbx_1__1__77_top_grid_pin_20_;
wire [0:0] cbx_1__1__77_top_grid_pin_21_;
wire [0:0] cbx_1__1__77_top_grid_pin_22_;
wire [0:0] cbx_1__1__77_top_grid_pin_23_;
wire [0:0] cbx_1__1__77_top_grid_pin_24_;
wire [0:0] cbx_1__1__77_top_grid_pin_25_;
wire [0:0] cbx_1__1__77_top_grid_pin_26_;
wire [0:0] cbx_1__1__77_top_grid_pin_27_;
wire [0:0] cbx_1__1__77_top_grid_pin_28_;
wire [0:0] cbx_1__1__77_top_grid_pin_29_;
wire [0:0] cbx_1__1__77_top_grid_pin_30_;
wire [0:0] cbx_1__1__77_top_grid_pin_31_;
wire [0:0] cbx_1__1__78_ccff_tail;
wire [0:19] cbx_1__1__78_chanx_left_out;
wire [0:19] cbx_1__1__78_chanx_right_out;
wire [0:0] cbx_1__1__78_top_grid_pin_16_;
wire [0:0] cbx_1__1__78_top_grid_pin_17_;
wire [0:0] cbx_1__1__78_top_grid_pin_18_;
wire [0:0] cbx_1__1__78_top_grid_pin_19_;
wire [0:0] cbx_1__1__78_top_grid_pin_20_;
wire [0:0] cbx_1__1__78_top_grid_pin_21_;
wire [0:0] cbx_1__1__78_top_grid_pin_22_;
wire [0:0] cbx_1__1__78_top_grid_pin_23_;
wire [0:0] cbx_1__1__78_top_grid_pin_24_;
wire [0:0] cbx_1__1__78_top_grid_pin_25_;
wire [0:0] cbx_1__1__78_top_grid_pin_26_;
wire [0:0] cbx_1__1__78_top_grid_pin_27_;
wire [0:0] cbx_1__1__78_top_grid_pin_28_;
wire [0:0] cbx_1__1__78_top_grid_pin_29_;
wire [0:0] cbx_1__1__78_top_grid_pin_30_;
wire [0:0] cbx_1__1__78_top_grid_pin_31_;
wire [0:0] cbx_1__1__79_ccff_tail;
wire [0:19] cbx_1__1__79_chanx_left_out;
wire [0:19] cbx_1__1__79_chanx_right_out;
wire [0:0] cbx_1__1__79_top_grid_pin_16_;
wire [0:0] cbx_1__1__79_top_grid_pin_17_;
wire [0:0] cbx_1__1__79_top_grid_pin_18_;
wire [0:0] cbx_1__1__79_top_grid_pin_19_;
wire [0:0] cbx_1__1__79_top_grid_pin_20_;
wire [0:0] cbx_1__1__79_top_grid_pin_21_;
wire [0:0] cbx_1__1__79_top_grid_pin_22_;
wire [0:0] cbx_1__1__79_top_grid_pin_23_;
wire [0:0] cbx_1__1__79_top_grid_pin_24_;
wire [0:0] cbx_1__1__79_top_grid_pin_25_;
wire [0:0] cbx_1__1__79_top_grid_pin_26_;
wire [0:0] cbx_1__1__79_top_grid_pin_27_;
wire [0:0] cbx_1__1__79_top_grid_pin_28_;
wire [0:0] cbx_1__1__79_top_grid_pin_29_;
wire [0:0] cbx_1__1__79_top_grid_pin_30_;
wire [0:0] cbx_1__1__79_top_grid_pin_31_;
wire [0:0] cbx_1__1__7_ccff_tail;
wire [0:19] cbx_1__1__7_chanx_left_out;
wire [0:19] cbx_1__1__7_chanx_right_out;
wire [0:0] cbx_1__1__7_top_grid_pin_16_;
wire [0:0] cbx_1__1__7_top_grid_pin_17_;
wire [0:0] cbx_1__1__7_top_grid_pin_18_;
wire [0:0] cbx_1__1__7_top_grid_pin_19_;
wire [0:0] cbx_1__1__7_top_grid_pin_20_;
wire [0:0] cbx_1__1__7_top_grid_pin_21_;
wire [0:0] cbx_1__1__7_top_grid_pin_22_;
wire [0:0] cbx_1__1__7_top_grid_pin_23_;
wire [0:0] cbx_1__1__7_top_grid_pin_24_;
wire [0:0] cbx_1__1__7_top_grid_pin_25_;
wire [0:0] cbx_1__1__7_top_grid_pin_26_;
wire [0:0] cbx_1__1__7_top_grid_pin_27_;
wire [0:0] cbx_1__1__7_top_grid_pin_28_;
wire [0:0] cbx_1__1__7_top_grid_pin_29_;
wire [0:0] cbx_1__1__7_top_grid_pin_30_;
wire [0:0] cbx_1__1__7_top_grid_pin_31_;
wire [0:0] cbx_1__1__80_ccff_tail;
wire [0:19] cbx_1__1__80_chanx_left_out;
wire [0:19] cbx_1__1__80_chanx_right_out;
wire [0:0] cbx_1__1__80_top_grid_pin_16_;
wire [0:0] cbx_1__1__80_top_grid_pin_17_;
wire [0:0] cbx_1__1__80_top_grid_pin_18_;
wire [0:0] cbx_1__1__80_top_grid_pin_19_;
wire [0:0] cbx_1__1__80_top_grid_pin_20_;
wire [0:0] cbx_1__1__80_top_grid_pin_21_;
wire [0:0] cbx_1__1__80_top_grid_pin_22_;
wire [0:0] cbx_1__1__80_top_grid_pin_23_;
wire [0:0] cbx_1__1__80_top_grid_pin_24_;
wire [0:0] cbx_1__1__80_top_grid_pin_25_;
wire [0:0] cbx_1__1__80_top_grid_pin_26_;
wire [0:0] cbx_1__1__80_top_grid_pin_27_;
wire [0:0] cbx_1__1__80_top_grid_pin_28_;
wire [0:0] cbx_1__1__80_top_grid_pin_29_;
wire [0:0] cbx_1__1__80_top_grid_pin_30_;
wire [0:0] cbx_1__1__80_top_grid_pin_31_;
wire [0:0] cbx_1__1__81_ccff_tail;
wire [0:19] cbx_1__1__81_chanx_left_out;
wire [0:19] cbx_1__1__81_chanx_right_out;
wire [0:0] cbx_1__1__81_top_grid_pin_16_;
wire [0:0] cbx_1__1__81_top_grid_pin_17_;
wire [0:0] cbx_1__1__81_top_grid_pin_18_;
wire [0:0] cbx_1__1__81_top_grid_pin_19_;
wire [0:0] cbx_1__1__81_top_grid_pin_20_;
wire [0:0] cbx_1__1__81_top_grid_pin_21_;
wire [0:0] cbx_1__1__81_top_grid_pin_22_;
wire [0:0] cbx_1__1__81_top_grid_pin_23_;
wire [0:0] cbx_1__1__81_top_grid_pin_24_;
wire [0:0] cbx_1__1__81_top_grid_pin_25_;
wire [0:0] cbx_1__1__81_top_grid_pin_26_;
wire [0:0] cbx_1__1__81_top_grid_pin_27_;
wire [0:0] cbx_1__1__81_top_grid_pin_28_;
wire [0:0] cbx_1__1__81_top_grid_pin_29_;
wire [0:0] cbx_1__1__81_top_grid_pin_30_;
wire [0:0] cbx_1__1__81_top_grid_pin_31_;
wire [0:0] cbx_1__1__82_ccff_tail;
wire [0:19] cbx_1__1__82_chanx_left_out;
wire [0:19] cbx_1__1__82_chanx_right_out;
wire [0:0] cbx_1__1__82_top_grid_pin_16_;
wire [0:0] cbx_1__1__82_top_grid_pin_17_;
wire [0:0] cbx_1__1__82_top_grid_pin_18_;
wire [0:0] cbx_1__1__82_top_grid_pin_19_;
wire [0:0] cbx_1__1__82_top_grid_pin_20_;
wire [0:0] cbx_1__1__82_top_grid_pin_21_;
wire [0:0] cbx_1__1__82_top_grid_pin_22_;
wire [0:0] cbx_1__1__82_top_grid_pin_23_;
wire [0:0] cbx_1__1__82_top_grid_pin_24_;
wire [0:0] cbx_1__1__82_top_grid_pin_25_;
wire [0:0] cbx_1__1__82_top_grid_pin_26_;
wire [0:0] cbx_1__1__82_top_grid_pin_27_;
wire [0:0] cbx_1__1__82_top_grid_pin_28_;
wire [0:0] cbx_1__1__82_top_grid_pin_29_;
wire [0:0] cbx_1__1__82_top_grid_pin_30_;
wire [0:0] cbx_1__1__82_top_grid_pin_31_;
wire [0:0] cbx_1__1__83_ccff_tail;
wire [0:19] cbx_1__1__83_chanx_left_out;
wire [0:19] cbx_1__1__83_chanx_right_out;
wire [0:0] cbx_1__1__83_top_grid_pin_16_;
wire [0:0] cbx_1__1__83_top_grid_pin_17_;
wire [0:0] cbx_1__1__83_top_grid_pin_18_;
wire [0:0] cbx_1__1__83_top_grid_pin_19_;
wire [0:0] cbx_1__1__83_top_grid_pin_20_;
wire [0:0] cbx_1__1__83_top_grid_pin_21_;
wire [0:0] cbx_1__1__83_top_grid_pin_22_;
wire [0:0] cbx_1__1__83_top_grid_pin_23_;
wire [0:0] cbx_1__1__83_top_grid_pin_24_;
wire [0:0] cbx_1__1__83_top_grid_pin_25_;
wire [0:0] cbx_1__1__83_top_grid_pin_26_;
wire [0:0] cbx_1__1__83_top_grid_pin_27_;
wire [0:0] cbx_1__1__83_top_grid_pin_28_;
wire [0:0] cbx_1__1__83_top_grid_pin_29_;
wire [0:0] cbx_1__1__83_top_grid_pin_30_;
wire [0:0] cbx_1__1__83_top_grid_pin_31_;
wire [0:0] cbx_1__1__84_ccff_tail;
wire [0:19] cbx_1__1__84_chanx_left_out;
wire [0:19] cbx_1__1__84_chanx_right_out;
wire [0:0] cbx_1__1__84_top_grid_pin_16_;
wire [0:0] cbx_1__1__84_top_grid_pin_17_;
wire [0:0] cbx_1__1__84_top_grid_pin_18_;
wire [0:0] cbx_1__1__84_top_grid_pin_19_;
wire [0:0] cbx_1__1__84_top_grid_pin_20_;
wire [0:0] cbx_1__1__84_top_grid_pin_21_;
wire [0:0] cbx_1__1__84_top_grid_pin_22_;
wire [0:0] cbx_1__1__84_top_grid_pin_23_;
wire [0:0] cbx_1__1__84_top_grid_pin_24_;
wire [0:0] cbx_1__1__84_top_grid_pin_25_;
wire [0:0] cbx_1__1__84_top_grid_pin_26_;
wire [0:0] cbx_1__1__84_top_grid_pin_27_;
wire [0:0] cbx_1__1__84_top_grid_pin_28_;
wire [0:0] cbx_1__1__84_top_grid_pin_29_;
wire [0:0] cbx_1__1__84_top_grid_pin_30_;
wire [0:0] cbx_1__1__84_top_grid_pin_31_;
wire [0:0] cbx_1__1__85_ccff_tail;
wire [0:19] cbx_1__1__85_chanx_left_out;
wire [0:19] cbx_1__1__85_chanx_right_out;
wire [0:0] cbx_1__1__85_top_grid_pin_16_;
wire [0:0] cbx_1__1__85_top_grid_pin_17_;
wire [0:0] cbx_1__1__85_top_grid_pin_18_;
wire [0:0] cbx_1__1__85_top_grid_pin_19_;
wire [0:0] cbx_1__1__85_top_grid_pin_20_;
wire [0:0] cbx_1__1__85_top_grid_pin_21_;
wire [0:0] cbx_1__1__85_top_grid_pin_22_;
wire [0:0] cbx_1__1__85_top_grid_pin_23_;
wire [0:0] cbx_1__1__85_top_grid_pin_24_;
wire [0:0] cbx_1__1__85_top_grid_pin_25_;
wire [0:0] cbx_1__1__85_top_grid_pin_26_;
wire [0:0] cbx_1__1__85_top_grid_pin_27_;
wire [0:0] cbx_1__1__85_top_grid_pin_28_;
wire [0:0] cbx_1__1__85_top_grid_pin_29_;
wire [0:0] cbx_1__1__85_top_grid_pin_30_;
wire [0:0] cbx_1__1__85_top_grid_pin_31_;
wire [0:0] cbx_1__1__86_ccff_tail;
wire [0:19] cbx_1__1__86_chanx_left_out;
wire [0:19] cbx_1__1__86_chanx_right_out;
wire [0:0] cbx_1__1__86_top_grid_pin_16_;
wire [0:0] cbx_1__1__86_top_grid_pin_17_;
wire [0:0] cbx_1__1__86_top_grid_pin_18_;
wire [0:0] cbx_1__1__86_top_grid_pin_19_;
wire [0:0] cbx_1__1__86_top_grid_pin_20_;
wire [0:0] cbx_1__1__86_top_grid_pin_21_;
wire [0:0] cbx_1__1__86_top_grid_pin_22_;
wire [0:0] cbx_1__1__86_top_grid_pin_23_;
wire [0:0] cbx_1__1__86_top_grid_pin_24_;
wire [0:0] cbx_1__1__86_top_grid_pin_25_;
wire [0:0] cbx_1__1__86_top_grid_pin_26_;
wire [0:0] cbx_1__1__86_top_grid_pin_27_;
wire [0:0] cbx_1__1__86_top_grid_pin_28_;
wire [0:0] cbx_1__1__86_top_grid_pin_29_;
wire [0:0] cbx_1__1__86_top_grid_pin_30_;
wire [0:0] cbx_1__1__86_top_grid_pin_31_;
wire [0:0] cbx_1__1__87_ccff_tail;
wire [0:19] cbx_1__1__87_chanx_left_out;
wire [0:19] cbx_1__1__87_chanx_right_out;
wire [0:0] cbx_1__1__87_top_grid_pin_16_;
wire [0:0] cbx_1__1__87_top_grid_pin_17_;
wire [0:0] cbx_1__1__87_top_grid_pin_18_;
wire [0:0] cbx_1__1__87_top_grid_pin_19_;
wire [0:0] cbx_1__1__87_top_grid_pin_20_;
wire [0:0] cbx_1__1__87_top_grid_pin_21_;
wire [0:0] cbx_1__1__87_top_grid_pin_22_;
wire [0:0] cbx_1__1__87_top_grid_pin_23_;
wire [0:0] cbx_1__1__87_top_grid_pin_24_;
wire [0:0] cbx_1__1__87_top_grid_pin_25_;
wire [0:0] cbx_1__1__87_top_grid_pin_26_;
wire [0:0] cbx_1__1__87_top_grid_pin_27_;
wire [0:0] cbx_1__1__87_top_grid_pin_28_;
wire [0:0] cbx_1__1__87_top_grid_pin_29_;
wire [0:0] cbx_1__1__87_top_grid_pin_30_;
wire [0:0] cbx_1__1__87_top_grid_pin_31_;
wire [0:0] cbx_1__1__88_ccff_tail;
wire [0:19] cbx_1__1__88_chanx_left_out;
wire [0:19] cbx_1__1__88_chanx_right_out;
wire [0:0] cbx_1__1__88_top_grid_pin_16_;
wire [0:0] cbx_1__1__88_top_grid_pin_17_;
wire [0:0] cbx_1__1__88_top_grid_pin_18_;
wire [0:0] cbx_1__1__88_top_grid_pin_19_;
wire [0:0] cbx_1__1__88_top_grid_pin_20_;
wire [0:0] cbx_1__1__88_top_grid_pin_21_;
wire [0:0] cbx_1__1__88_top_grid_pin_22_;
wire [0:0] cbx_1__1__88_top_grid_pin_23_;
wire [0:0] cbx_1__1__88_top_grid_pin_24_;
wire [0:0] cbx_1__1__88_top_grid_pin_25_;
wire [0:0] cbx_1__1__88_top_grid_pin_26_;
wire [0:0] cbx_1__1__88_top_grid_pin_27_;
wire [0:0] cbx_1__1__88_top_grid_pin_28_;
wire [0:0] cbx_1__1__88_top_grid_pin_29_;
wire [0:0] cbx_1__1__88_top_grid_pin_30_;
wire [0:0] cbx_1__1__88_top_grid_pin_31_;
wire [0:0] cbx_1__1__89_ccff_tail;
wire [0:19] cbx_1__1__89_chanx_left_out;
wire [0:19] cbx_1__1__89_chanx_right_out;
wire [0:0] cbx_1__1__89_top_grid_pin_16_;
wire [0:0] cbx_1__1__89_top_grid_pin_17_;
wire [0:0] cbx_1__1__89_top_grid_pin_18_;
wire [0:0] cbx_1__1__89_top_grid_pin_19_;
wire [0:0] cbx_1__1__89_top_grid_pin_20_;
wire [0:0] cbx_1__1__89_top_grid_pin_21_;
wire [0:0] cbx_1__1__89_top_grid_pin_22_;
wire [0:0] cbx_1__1__89_top_grid_pin_23_;
wire [0:0] cbx_1__1__89_top_grid_pin_24_;
wire [0:0] cbx_1__1__89_top_grid_pin_25_;
wire [0:0] cbx_1__1__89_top_grid_pin_26_;
wire [0:0] cbx_1__1__89_top_grid_pin_27_;
wire [0:0] cbx_1__1__89_top_grid_pin_28_;
wire [0:0] cbx_1__1__89_top_grid_pin_29_;
wire [0:0] cbx_1__1__89_top_grid_pin_30_;
wire [0:0] cbx_1__1__89_top_grid_pin_31_;
wire [0:0] cbx_1__1__8_ccff_tail;
wire [0:19] cbx_1__1__8_chanx_left_out;
wire [0:19] cbx_1__1__8_chanx_right_out;
wire [0:0] cbx_1__1__8_top_grid_pin_16_;
wire [0:0] cbx_1__1__8_top_grid_pin_17_;
wire [0:0] cbx_1__1__8_top_grid_pin_18_;
wire [0:0] cbx_1__1__8_top_grid_pin_19_;
wire [0:0] cbx_1__1__8_top_grid_pin_20_;
wire [0:0] cbx_1__1__8_top_grid_pin_21_;
wire [0:0] cbx_1__1__8_top_grid_pin_22_;
wire [0:0] cbx_1__1__8_top_grid_pin_23_;
wire [0:0] cbx_1__1__8_top_grid_pin_24_;
wire [0:0] cbx_1__1__8_top_grid_pin_25_;
wire [0:0] cbx_1__1__8_top_grid_pin_26_;
wire [0:0] cbx_1__1__8_top_grid_pin_27_;
wire [0:0] cbx_1__1__8_top_grid_pin_28_;
wire [0:0] cbx_1__1__8_top_grid_pin_29_;
wire [0:0] cbx_1__1__8_top_grid_pin_30_;
wire [0:0] cbx_1__1__8_top_grid_pin_31_;
wire [0:0] cbx_1__1__90_ccff_tail;
wire [0:19] cbx_1__1__90_chanx_left_out;
wire [0:19] cbx_1__1__90_chanx_right_out;
wire [0:0] cbx_1__1__90_top_grid_pin_16_;
wire [0:0] cbx_1__1__90_top_grid_pin_17_;
wire [0:0] cbx_1__1__90_top_grid_pin_18_;
wire [0:0] cbx_1__1__90_top_grid_pin_19_;
wire [0:0] cbx_1__1__90_top_grid_pin_20_;
wire [0:0] cbx_1__1__90_top_grid_pin_21_;
wire [0:0] cbx_1__1__90_top_grid_pin_22_;
wire [0:0] cbx_1__1__90_top_grid_pin_23_;
wire [0:0] cbx_1__1__90_top_grid_pin_24_;
wire [0:0] cbx_1__1__90_top_grid_pin_25_;
wire [0:0] cbx_1__1__90_top_grid_pin_26_;
wire [0:0] cbx_1__1__90_top_grid_pin_27_;
wire [0:0] cbx_1__1__90_top_grid_pin_28_;
wire [0:0] cbx_1__1__90_top_grid_pin_29_;
wire [0:0] cbx_1__1__90_top_grid_pin_30_;
wire [0:0] cbx_1__1__90_top_grid_pin_31_;
wire [0:0] cbx_1__1__91_ccff_tail;
wire [0:19] cbx_1__1__91_chanx_left_out;
wire [0:19] cbx_1__1__91_chanx_right_out;
wire [0:0] cbx_1__1__91_top_grid_pin_16_;
wire [0:0] cbx_1__1__91_top_grid_pin_17_;
wire [0:0] cbx_1__1__91_top_grid_pin_18_;
wire [0:0] cbx_1__1__91_top_grid_pin_19_;
wire [0:0] cbx_1__1__91_top_grid_pin_20_;
wire [0:0] cbx_1__1__91_top_grid_pin_21_;
wire [0:0] cbx_1__1__91_top_grid_pin_22_;
wire [0:0] cbx_1__1__91_top_grid_pin_23_;
wire [0:0] cbx_1__1__91_top_grid_pin_24_;
wire [0:0] cbx_1__1__91_top_grid_pin_25_;
wire [0:0] cbx_1__1__91_top_grid_pin_26_;
wire [0:0] cbx_1__1__91_top_grid_pin_27_;
wire [0:0] cbx_1__1__91_top_grid_pin_28_;
wire [0:0] cbx_1__1__91_top_grid_pin_29_;
wire [0:0] cbx_1__1__91_top_grid_pin_30_;
wire [0:0] cbx_1__1__91_top_grid_pin_31_;
wire [0:0] cbx_1__1__92_ccff_tail;
wire [0:19] cbx_1__1__92_chanx_left_out;
wire [0:19] cbx_1__1__92_chanx_right_out;
wire [0:0] cbx_1__1__92_top_grid_pin_16_;
wire [0:0] cbx_1__1__92_top_grid_pin_17_;
wire [0:0] cbx_1__1__92_top_grid_pin_18_;
wire [0:0] cbx_1__1__92_top_grid_pin_19_;
wire [0:0] cbx_1__1__92_top_grid_pin_20_;
wire [0:0] cbx_1__1__92_top_grid_pin_21_;
wire [0:0] cbx_1__1__92_top_grid_pin_22_;
wire [0:0] cbx_1__1__92_top_grid_pin_23_;
wire [0:0] cbx_1__1__92_top_grid_pin_24_;
wire [0:0] cbx_1__1__92_top_grid_pin_25_;
wire [0:0] cbx_1__1__92_top_grid_pin_26_;
wire [0:0] cbx_1__1__92_top_grid_pin_27_;
wire [0:0] cbx_1__1__92_top_grid_pin_28_;
wire [0:0] cbx_1__1__92_top_grid_pin_29_;
wire [0:0] cbx_1__1__92_top_grid_pin_30_;
wire [0:0] cbx_1__1__92_top_grid_pin_31_;
wire [0:0] cbx_1__1__93_ccff_tail;
wire [0:19] cbx_1__1__93_chanx_left_out;
wire [0:19] cbx_1__1__93_chanx_right_out;
wire [0:0] cbx_1__1__93_top_grid_pin_16_;
wire [0:0] cbx_1__1__93_top_grid_pin_17_;
wire [0:0] cbx_1__1__93_top_grid_pin_18_;
wire [0:0] cbx_1__1__93_top_grid_pin_19_;
wire [0:0] cbx_1__1__93_top_grid_pin_20_;
wire [0:0] cbx_1__1__93_top_grid_pin_21_;
wire [0:0] cbx_1__1__93_top_grid_pin_22_;
wire [0:0] cbx_1__1__93_top_grid_pin_23_;
wire [0:0] cbx_1__1__93_top_grid_pin_24_;
wire [0:0] cbx_1__1__93_top_grid_pin_25_;
wire [0:0] cbx_1__1__93_top_grid_pin_26_;
wire [0:0] cbx_1__1__93_top_grid_pin_27_;
wire [0:0] cbx_1__1__93_top_grid_pin_28_;
wire [0:0] cbx_1__1__93_top_grid_pin_29_;
wire [0:0] cbx_1__1__93_top_grid_pin_30_;
wire [0:0] cbx_1__1__93_top_grid_pin_31_;
wire [0:0] cbx_1__1__94_ccff_tail;
wire [0:19] cbx_1__1__94_chanx_left_out;
wire [0:19] cbx_1__1__94_chanx_right_out;
wire [0:0] cbx_1__1__94_top_grid_pin_16_;
wire [0:0] cbx_1__1__94_top_grid_pin_17_;
wire [0:0] cbx_1__1__94_top_grid_pin_18_;
wire [0:0] cbx_1__1__94_top_grid_pin_19_;
wire [0:0] cbx_1__1__94_top_grid_pin_20_;
wire [0:0] cbx_1__1__94_top_grid_pin_21_;
wire [0:0] cbx_1__1__94_top_grid_pin_22_;
wire [0:0] cbx_1__1__94_top_grid_pin_23_;
wire [0:0] cbx_1__1__94_top_grid_pin_24_;
wire [0:0] cbx_1__1__94_top_grid_pin_25_;
wire [0:0] cbx_1__1__94_top_grid_pin_26_;
wire [0:0] cbx_1__1__94_top_grid_pin_27_;
wire [0:0] cbx_1__1__94_top_grid_pin_28_;
wire [0:0] cbx_1__1__94_top_grid_pin_29_;
wire [0:0] cbx_1__1__94_top_grid_pin_30_;
wire [0:0] cbx_1__1__94_top_grid_pin_31_;
wire [0:0] cbx_1__1__95_ccff_tail;
wire [0:19] cbx_1__1__95_chanx_left_out;
wire [0:19] cbx_1__1__95_chanx_right_out;
wire [0:0] cbx_1__1__95_top_grid_pin_16_;
wire [0:0] cbx_1__1__95_top_grid_pin_17_;
wire [0:0] cbx_1__1__95_top_grid_pin_18_;
wire [0:0] cbx_1__1__95_top_grid_pin_19_;
wire [0:0] cbx_1__1__95_top_grid_pin_20_;
wire [0:0] cbx_1__1__95_top_grid_pin_21_;
wire [0:0] cbx_1__1__95_top_grid_pin_22_;
wire [0:0] cbx_1__1__95_top_grid_pin_23_;
wire [0:0] cbx_1__1__95_top_grid_pin_24_;
wire [0:0] cbx_1__1__95_top_grid_pin_25_;
wire [0:0] cbx_1__1__95_top_grid_pin_26_;
wire [0:0] cbx_1__1__95_top_grid_pin_27_;
wire [0:0] cbx_1__1__95_top_grid_pin_28_;
wire [0:0] cbx_1__1__95_top_grid_pin_29_;
wire [0:0] cbx_1__1__95_top_grid_pin_30_;
wire [0:0] cbx_1__1__95_top_grid_pin_31_;
wire [0:0] cbx_1__1__96_ccff_tail;
wire [0:19] cbx_1__1__96_chanx_left_out;
wire [0:19] cbx_1__1__96_chanx_right_out;
wire [0:0] cbx_1__1__96_top_grid_pin_16_;
wire [0:0] cbx_1__1__96_top_grid_pin_17_;
wire [0:0] cbx_1__1__96_top_grid_pin_18_;
wire [0:0] cbx_1__1__96_top_grid_pin_19_;
wire [0:0] cbx_1__1__96_top_grid_pin_20_;
wire [0:0] cbx_1__1__96_top_grid_pin_21_;
wire [0:0] cbx_1__1__96_top_grid_pin_22_;
wire [0:0] cbx_1__1__96_top_grid_pin_23_;
wire [0:0] cbx_1__1__96_top_grid_pin_24_;
wire [0:0] cbx_1__1__96_top_grid_pin_25_;
wire [0:0] cbx_1__1__96_top_grid_pin_26_;
wire [0:0] cbx_1__1__96_top_grid_pin_27_;
wire [0:0] cbx_1__1__96_top_grid_pin_28_;
wire [0:0] cbx_1__1__96_top_grid_pin_29_;
wire [0:0] cbx_1__1__96_top_grid_pin_30_;
wire [0:0] cbx_1__1__96_top_grid_pin_31_;
wire [0:0] cbx_1__1__97_ccff_tail;
wire [0:19] cbx_1__1__97_chanx_left_out;
wire [0:19] cbx_1__1__97_chanx_right_out;
wire [0:0] cbx_1__1__97_top_grid_pin_16_;
wire [0:0] cbx_1__1__97_top_grid_pin_17_;
wire [0:0] cbx_1__1__97_top_grid_pin_18_;
wire [0:0] cbx_1__1__97_top_grid_pin_19_;
wire [0:0] cbx_1__1__97_top_grid_pin_20_;
wire [0:0] cbx_1__1__97_top_grid_pin_21_;
wire [0:0] cbx_1__1__97_top_grid_pin_22_;
wire [0:0] cbx_1__1__97_top_grid_pin_23_;
wire [0:0] cbx_1__1__97_top_grid_pin_24_;
wire [0:0] cbx_1__1__97_top_grid_pin_25_;
wire [0:0] cbx_1__1__97_top_grid_pin_26_;
wire [0:0] cbx_1__1__97_top_grid_pin_27_;
wire [0:0] cbx_1__1__97_top_grid_pin_28_;
wire [0:0] cbx_1__1__97_top_grid_pin_29_;
wire [0:0] cbx_1__1__97_top_grid_pin_30_;
wire [0:0] cbx_1__1__97_top_grid_pin_31_;
wire [0:0] cbx_1__1__98_ccff_tail;
wire [0:19] cbx_1__1__98_chanx_left_out;
wire [0:19] cbx_1__1__98_chanx_right_out;
wire [0:0] cbx_1__1__98_top_grid_pin_16_;
wire [0:0] cbx_1__1__98_top_grid_pin_17_;
wire [0:0] cbx_1__1__98_top_grid_pin_18_;
wire [0:0] cbx_1__1__98_top_grid_pin_19_;
wire [0:0] cbx_1__1__98_top_grid_pin_20_;
wire [0:0] cbx_1__1__98_top_grid_pin_21_;
wire [0:0] cbx_1__1__98_top_grid_pin_22_;
wire [0:0] cbx_1__1__98_top_grid_pin_23_;
wire [0:0] cbx_1__1__98_top_grid_pin_24_;
wire [0:0] cbx_1__1__98_top_grid_pin_25_;
wire [0:0] cbx_1__1__98_top_grid_pin_26_;
wire [0:0] cbx_1__1__98_top_grid_pin_27_;
wire [0:0] cbx_1__1__98_top_grid_pin_28_;
wire [0:0] cbx_1__1__98_top_grid_pin_29_;
wire [0:0] cbx_1__1__98_top_grid_pin_30_;
wire [0:0] cbx_1__1__98_top_grid_pin_31_;
wire [0:0] cbx_1__1__99_ccff_tail;
wire [0:19] cbx_1__1__99_chanx_left_out;
wire [0:19] cbx_1__1__99_chanx_right_out;
wire [0:0] cbx_1__1__99_top_grid_pin_16_;
wire [0:0] cbx_1__1__99_top_grid_pin_17_;
wire [0:0] cbx_1__1__99_top_grid_pin_18_;
wire [0:0] cbx_1__1__99_top_grid_pin_19_;
wire [0:0] cbx_1__1__99_top_grid_pin_20_;
wire [0:0] cbx_1__1__99_top_grid_pin_21_;
wire [0:0] cbx_1__1__99_top_grid_pin_22_;
wire [0:0] cbx_1__1__99_top_grid_pin_23_;
wire [0:0] cbx_1__1__99_top_grid_pin_24_;
wire [0:0] cbx_1__1__99_top_grid_pin_25_;
wire [0:0] cbx_1__1__99_top_grid_pin_26_;
wire [0:0] cbx_1__1__99_top_grid_pin_27_;
wire [0:0] cbx_1__1__99_top_grid_pin_28_;
wire [0:0] cbx_1__1__99_top_grid_pin_29_;
wire [0:0] cbx_1__1__99_top_grid_pin_30_;
wire [0:0] cbx_1__1__99_top_grid_pin_31_;
wire [0:0] cbx_1__1__9_ccff_tail;
wire [0:19] cbx_1__1__9_chanx_left_out;
wire [0:19] cbx_1__1__9_chanx_right_out;
wire [0:0] cbx_1__1__9_top_grid_pin_16_;
wire [0:0] cbx_1__1__9_top_grid_pin_17_;
wire [0:0] cbx_1__1__9_top_grid_pin_18_;
wire [0:0] cbx_1__1__9_top_grid_pin_19_;
wire [0:0] cbx_1__1__9_top_grid_pin_20_;
wire [0:0] cbx_1__1__9_top_grid_pin_21_;
wire [0:0] cbx_1__1__9_top_grid_pin_22_;
wire [0:0] cbx_1__1__9_top_grid_pin_23_;
wire [0:0] cbx_1__1__9_top_grid_pin_24_;
wire [0:0] cbx_1__1__9_top_grid_pin_25_;
wire [0:0] cbx_1__1__9_top_grid_pin_26_;
wire [0:0] cbx_1__1__9_top_grid_pin_27_;
wire [0:0] cbx_1__1__9_top_grid_pin_28_;
wire [0:0] cbx_1__1__9_top_grid_pin_29_;
wire [0:0] cbx_1__1__9_top_grid_pin_30_;
wire [0:0] cbx_1__1__9_top_grid_pin_31_;
wire [0:0] cby_0__1__0_ccff_tail;
wire [0:19] cby_0__1__0_chany_bottom_out;
wire [0:19] cby_0__1__0_chany_top_out;
wire [0:0] cby_0__1__0_left_grid_pin_0_;
wire [0:0] cby_0__1__0_right_grid_pin_52_;
wire [0:0] cby_0__1__10_ccff_tail;
wire [0:19] cby_0__1__10_chany_bottom_out;
wire [0:19] cby_0__1__10_chany_top_out;
wire [0:0] cby_0__1__10_left_grid_pin_0_;
wire [0:0] cby_0__1__10_right_grid_pin_52_;
wire [0:0] cby_0__1__11_ccff_tail;
wire [0:19] cby_0__1__11_chany_bottom_out;
wire [0:19] cby_0__1__11_chany_top_out;
wire [0:0] cby_0__1__11_left_grid_pin_0_;
wire [0:0] cby_0__1__11_right_grid_pin_52_;
wire [0:0] cby_0__1__1_ccff_tail;
wire [0:19] cby_0__1__1_chany_bottom_out;
wire [0:19] cby_0__1__1_chany_top_out;
wire [0:0] cby_0__1__1_left_grid_pin_0_;
wire [0:0] cby_0__1__1_right_grid_pin_52_;
wire [0:0] cby_0__1__2_ccff_tail;
wire [0:19] cby_0__1__2_chany_bottom_out;
wire [0:19] cby_0__1__2_chany_top_out;
wire [0:0] cby_0__1__2_left_grid_pin_0_;
wire [0:0] cby_0__1__2_right_grid_pin_52_;
wire [0:0] cby_0__1__3_ccff_tail;
wire [0:19] cby_0__1__3_chany_bottom_out;
wire [0:19] cby_0__1__3_chany_top_out;
wire [0:0] cby_0__1__3_left_grid_pin_0_;
wire [0:0] cby_0__1__3_right_grid_pin_52_;
wire [0:0] cby_0__1__4_ccff_tail;
wire [0:19] cby_0__1__4_chany_bottom_out;
wire [0:19] cby_0__1__4_chany_top_out;
wire [0:0] cby_0__1__4_left_grid_pin_0_;
wire [0:0] cby_0__1__4_right_grid_pin_52_;
wire [0:0] cby_0__1__5_ccff_tail;
wire [0:19] cby_0__1__5_chany_bottom_out;
wire [0:19] cby_0__1__5_chany_top_out;
wire [0:0] cby_0__1__5_left_grid_pin_0_;
wire [0:0] cby_0__1__5_right_grid_pin_52_;
wire [0:0] cby_0__1__6_ccff_tail;
wire [0:19] cby_0__1__6_chany_bottom_out;
wire [0:19] cby_0__1__6_chany_top_out;
wire [0:0] cby_0__1__6_left_grid_pin_0_;
wire [0:0] cby_0__1__6_right_grid_pin_52_;
wire [0:0] cby_0__1__7_ccff_tail;
wire [0:19] cby_0__1__7_chany_bottom_out;
wire [0:19] cby_0__1__7_chany_top_out;
wire [0:0] cby_0__1__7_left_grid_pin_0_;
wire [0:0] cby_0__1__7_right_grid_pin_52_;
wire [0:0] cby_0__1__8_ccff_tail;
wire [0:19] cby_0__1__8_chany_bottom_out;
wire [0:19] cby_0__1__8_chany_top_out;
wire [0:0] cby_0__1__8_left_grid_pin_0_;
wire [0:0] cby_0__1__8_right_grid_pin_52_;
wire [0:0] cby_0__1__9_ccff_tail;
wire [0:19] cby_0__1__9_chany_bottom_out;
wire [0:19] cby_0__1__9_chany_top_out;
wire [0:0] cby_0__1__9_left_grid_pin_0_;
wire [0:0] cby_0__1__9_right_grid_pin_52_;
wire [0:0] cby_1__1__0_ccff_tail;
wire [0:19] cby_1__1__0_chany_bottom_out;
wire [0:19] cby_1__1__0_chany_top_out;
wire [0:0] cby_1__1__0_left_grid_pin_0_;
wire [0:0] cby_1__1__0_left_grid_pin_10_;
wire [0:0] cby_1__1__0_left_grid_pin_11_;
wire [0:0] cby_1__1__0_left_grid_pin_12_;
wire [0:0] cby_1__1__0_left_grid_pin_13_;
wire [0:0] cby_1__1__0_left_grid_pin_14_;
wire [0:0] cby_1__1__0_left_grid_pin_15_;
wire [0:0] cby_1__1__0_left_grid_pin_1_;
wire [0:0] cby_1__1__0_left_grid_pin_2_;
wire [0:0] cby_1__1__0_left_grid_pin_3_;
wire [0:0] cby_1__1__0_left_grid_pin_4_;
wire [0:0] cby_1__1__0_left_grid_pin_5_;
wire [0:0] cby_1__1__0_left_grid_pin_6_;
wire [0:0] cby_1__1__0_left_grid_pin_7_;
wire [0:0] cby_1__1__0_left_grid_pin_8_;
wire [0:0] cby_1__1__0_left_grid_pin_9_;
wire [0:0] cby_1__1__0_right_grid_pin_52_;
wire [0:0] cby_1__1__100_ccff_tail;
wire [0:19] cby_1__1__100_chany_bottom_out;
wire [0:19] cby_1__1__100_chany_top_out;
wire [0:0] cby_1__1__100_left_grid_pin_0_;
wire [0:0] cby_1__1__100_left_grid_pin_10_;
wire [0:0] cby_1__1__100_left_grid_pin_11_;
wire [0:0] cby_1__1__100_left_grid_pin_12_;
wire [0:0] cby_1__1__100_left_grid_pin_13_;
wire [0:0] cby_1__1__100_left_grid_pin_14_;
wire [0:0] cby_1__1__100_left_grid_pin_15_;
wire [0:0] cby_1__1__100_left_grid_pin_1_;
wire [0:0] cby_1__1__100_left_grid_pin_2_;
wire [0:0] cby_1__1__100_left_grid_pin_3_;
wire [0:0] cby_1__1__100_left_grid_pin_4_;
wire [0:0] cby_1__1__100_left_grid_pin_5_;
wire [0:0] cby_1__1__100_left_grid_pin_6_;
wire [0:0] cby_1__1__100_left_grid_pin_7_;
wire [0:0] cby_1__1__100_left_grid_pin_8_;
wire [0:0] cby_1__1__100_left_grid_pin_9_;
wire [0:0] cby_1__1__100_right_grid_pin_52_;
wire [0:0] cby_1__1__101_ccff_tail;
wire [0:19] cby_1__1__101_chany_bottom_out;
wire [0:19] cby_1__1__101_chany_top_out;
wire [0:0] cby_1__1__101_left_grid_pin_0_;
wire [0:0] cby_1__1__101_left_grid_pin_10_;
wire [0:0] cby_1__1__101_left_grid_pin_11_;
wire [0:0] cby_1__1__101_left_grid_pin_12_;
wire [0:0] cby_1__1__101_left_grid_pin_13_;
wire [0:0] cby_1__1__101_left_grid_pin_14_;
wire [0:0] cby_1__1__101_left_grid_pin_15_;
wire [0:0] cby_1__1__101_left_grid_pin_1_;
wire [0:0] cby_1__1__101_left_grid_pin_2_;
wire [0:0] cby_1__1__101_left_grid_pin_3_;
wire [0:0] cby_1__1__101_left_grid_pin_4_;
wire [0:0] cby_1__1__101_left_grid_pin_5_;
wire [0:0] cby_1__1__101_left_grid_pin_6_;
wire [0:0] cby_1__1__101_left_grid_pin_7_;
wire [0:0] cby_1__1__101_left_grid_pin_8_;
wire [0:0] cby_1__1__101_left_grid_pin_9_;
wire [0:0] cby_1__1__101_right_grid_pin_52_;
wire [0:0] cby_1__1__102_ccff_tail;
wire [0:19] cby_1__1__102_chany_bottom_out;
wire [0:19] cby_1__1__102_chany_top_out;
wire [0:0] cby_1__1__102_left_grid_pin_0_;
wire [0:0] cby_1__1__102_left_grid_pin_10_;
wire [0:0] cby_1__1__102_left_grid_pin_11_;
wire [0:0] cby_1__1__102_left_grid_pin_12_;
wire [0:0] cby_1__1__102_left_grid_pin_13_;
wire [0:0] cby_1__1__102_left_grid_pin_14_;
wire [0:0] cby_1__1__102_left_grid_pin_15_;
wire [0:0] cby_1__1__102_left_grid_pin_1_;
wire [0:0] cby_1__1__102_left_grid_pin_2_;
wire [0:0] cby_1__1__102_left_grid_pin_3_;
wire [0:0] cby_1__1__102_left_grid_pin_4_;
wire [0:0] cby_1__1__102_left_grid_pin_5_;
wire [0:0] cby_1__1__102_left_grid_pin_6_;
wire [0:0] cby_1__1__102_left_grid_pin_7_;
wire [0:0] cby_1__1__102_left_grid_pin_8_;
wire [0:0] cby_1__1__102_left_grid_pin_9_;
wire [0:0] cby_1__1__102_right_grid_pin_52_;
wire [0:0] cby_1__1__103_ccff_tail;
wire [0:19] cby_1__1__103_chany_bottom_out;
wire [0:19] cby_1__1__103_chany_top_out;
wire [0:0] cby_1__1__103_left_grid_pin_0_;
wire [0:0] cby_1__1__103_left_grid_pin_10_;
wire [0:0] cby_1__1__103_left_grid_pin_11_;
wire [0:0] cby_1__1__103_left_grid_pin_12_;
wire [0:0] cby_1__1__103_left_grid_pin_13_;
wire [0:0] cby_1__1__103_left_grid_pin_14_;
wire [0:0] cby_1__1__103_left_grid_pin_15_;
wire [0:0] cby_1__1__103_left_grid_pin_1_;
wire [0:0] cby_1__1__103_left_grid_pin_2_;
wire [0:0] cby_1__1__103_left_grid_pin_3_;
wire [0:0] cby_1__1__103_left_grid_pin_4_;
wire [0:0] cby_1__1__103_left_grid_pin_5_;
wire [0:0] cby_1__1__103_left_grid_pin_6_;
wire [0:0] cby_1__1__103_left_grid_pin_7_;
wire [0:0] cby_1__1__103_left_grid_pin_8_;
wire [0:0] cby_1__1__103_left_grid_pin_9_;
wire [0:0] cby_1__1__103_right_grid_pin_52_;
wire [0:0] cby_1__1__104_ccff_tail;
wire [0:19] cby_1__1__104_chany_bottom_out;
wire [0:19] cby_1__1__104_chany_top_out;
wire [0:0] cby_1__1__104_left_grid_pin_0_;
wire [0:0] cby_1__1__104_left_grid_pin_10_;
wire [0:0] cby_1__1__104_left_grid_pin_11_;
wire [0:0] cby_1__1__104_left_grid_pin_12_;
wire [0:0] cby_1__1__104_left_grid_pin_13_;
wire [0:0] cby_1__1__104_left_grid_pin_14_;
wire [0:0] cby_1__1__104_left_grid_pin_15_;
wire [0:0] cby_1__1__104_left_grid_pin_1_;
wire [0:0] cby_1__1__104_left_grid_pin_2_;
wire [0:0] cby_1__1__104_left_grid_pin_3_;
wire [0:0] cby_1__1__104_left_grid_pin_4_;
wire [0:0] cby_1__1__104_left_grid_pin_5_;
wire [0:0] cby_1__1__104_left_grid_pin_6_;
wire [0:0] cby_1__1__104_left_grid_pin_7_;
wire [0:0] cby_1__1__104_left_grid_pin_8_;
wire [0:0] cby_1__1__104_left_grid_pin_9_;
wire [0:0] cby_1__1__104_right_grid_pin_52_;
wire [0:0] cby_1__1__105_ccff_tail;
wire [0:19] cby_1__1__105_chany_bottom_out;
wire [0:19] cby_1__1__105_chany_top_out;
wire [0:0] cby_1__1__105_left_grid_pin_0_;
wire [0:0] cby_1__1__105_left_grid_pin_10_;
wire [0:0] cby_1__1__105_left_grid_pin_11_;
wire [0:0] cby_1__1__105_left_grid_pin_12_;
wire [0:0] cby_1__1__105_left_grid_pin_13_;
wire [0:0] cby_1__1__105_left_grid_pin_14_;
wire [0:0] cby_1__1__105_left_grid_pin_15_;
wire [0:0] cby_1__1__105_left_grid_pin_1_;
wire [0:0] cby_1__1__105_left_grid_pin_2_;
wire [0:0] cby_1__1__105_left_grid_pin_3_;
wire [0:0] cby_1__1__105_left_grid_pin_4_;
wire [0:0] cby_1__1__105_left_grid_pin_5_;
wire [0:0] cby_1__1__105_left_grid_pin_6_;
wire [0:0] cby_1__1__105_left_grid_pin_7_;
wire [0:0] cby_1__1__105_left_grid_pin_8_;
wire [0:0] cby_1__1__105_left_grid_pin_9_;
wire [0:0] cby_1__1__105_right_grid_pin_52_;
wire [0:0] cby_1__1__106_ccff_tail;
wire [0:19] cby_1__1__106_chany_bottom_out;
wire [0:19] cby_1__1__106_chany_top_out;
wire [0:0] cby_1__1__106_left_grid_pin_0_;
wire [0:0] cby_1__1__106_left_grid_pin_10_;
wire [0:0] cby_1__1__106_left_grid_pin_11_;
wire [0:0] cby_1__1__106_left_grid_pin_12_;
wire [0:0] cby_1__1__106_left_grid_pin_13_;
wire [0:0] cby_1__1__106_left_grid_pin_14_;
wire [0:0] cby_1__1__106_left_grid_pin_15_;
wire [0:0] cby_1__1__106_left_grid_pin_1_;
wire [0:0] cby_1__1__106_left_grid_pin_2_;
wire [0:0] cby_1__1__106_left_grid_pin_3_;
wire [0:0] cby_1__1__106_left_grid_pin_4_;
wire [0:0] cby_1__1__106_left_grid_pin_5_;
wire [0:0] cby_1__1__106_left_grid_pin_6_;
wire [0:0] cby_1__1__106_left_grid_pin_7_;
wire [0:0] cby_1__1__106_left_grid_pin_8_;
wire [0:0] cby_1__1__106_left_grid_pin_9_;
wire [0:0] cby_1__1__106_right_grid_pin_52_;
wire [0:0] cby_1__1__107_ccff_tail;
wire [0:19] cby_1__1__107_chany_bottom_out;
wire [0:19] cby_1__1__107_chany_top_out;
wire [0:0] cby_1__1__107_left_grid_pin_0_;
wire [0:0] cby_1__1__107_left_grid_pin_10_;
wire [0:0] cby_1__1__107_left_grid_pin_11_;
wire [0:0] cby_1__1__107_left_grid_pin_12_;
wire [0:0] cby_1__1__107_left_grid_pin_13_;
wire [0:0] cby_1__1__107_left_grid_pin_14_;
wire [0:0] cby_1__1__107_left_grid_pin_15_;
wire [0:0] cby_1__1__107_left_grid_pin_1_;
wire [0:0] cby_1__1__107_left_grid_pin_2_;
wire [0:0] cby_1__1__107_left_grid_pin_3_;
wire [0:0] cby_1__1__107_left_grid_pin_4_;
wire [0:0] cby_1__1__107_left_grid_pin_5_;
wire [0:0] cby_1__1__107_left_grid_pin_6_;
wire [0:0] cby_1__1__107_left_grid_pin_7_;
wire [0:0] cby_1__1__107_left_grid_pin_8_;
wire [0:0] cby_1__1__107_left_grid_pin_9_;
wire [0:0] cby_1__1__107_right_grid_pin_52_;
wire [0:0] cby_1__1__108_ccff_tail;
wire [0:19] cby_1__1__108_chany_bottom_out;
wire [0:19] cby_1__1__108_chany_top_out;
wire [0:0] cby_1__1__108_left_grid_pin_0_;
wire [0:0] cby_1__1__108_left_grid_pin_10_;
wire [0:0] cby_1__1__108_left_grid_pin_11_;
wire [0:0] cby_1__1__108_left_grid_pin_12_;
wire [0:0] cby_1__1__108_left_grid_pin_13_;
wire [0:0] cby_1__1__108_left_grid_pin_14_;
wire [0:0] cby_1__1__108_left_grid_pin_15_;
wire [0:0] cby_1__1__108_left_grid_pin_1_;
wire [0:0] cby_1__1__108_left_grid_pin_2_;
wire [0:0] cby_1__1__108_left_grid_pin_3_;
wire [0:0] cby_1__1__108_left_grid_pin_4_;
wire [0:0] cby_1__1__108_left_grid_pin_5_;
wire [0:0] cby_1__1__108_left_grid_pin_6_;
wire [0:0] cby_1__1__108_left_grid_pin_7_;
wire [0:0] cby_1__1__108_left_grid_pin_8_;
wire [0:0] cby_1__1__108_left_grid_pin_9_;
wire [0:0] cby_1__1__108_right_grid_pin_52_;
wire [0:0] cby_1__1__109_ccff_tail;
wire [0:19] cby_1__1__109_chany_bottom_out;
wire [0:19] cby_1__1__109_chany_top_out;
wire [0:0] cby_1__1__109_left_grid_pin_0_;
wire [0:0] cby_1__1__109_left_grid_pin_10_;
wire [0:0] cby_1__1__109_left_grid_pin_11_;
wire [0:0] cby_1__1__109_left_grid_pin_12_;
wire [0:0] cby_1__1__109_left_grid_pin_13_;
wire [0:0] cby_1__1__109_left_grid_pin_14_;
wire [0:0] cby_1__1__109_left_grid_pin_15_;
wire [0:0] cby_1__1__109_left_grid_pin_1_;
wire [0:0] cby_1__1__109_left_grid_pin_2_;
wire [0:0] cby_1__1__109_left_grid_pin_3_;
wire [0:0] cby_1__1__109_left_grid_pin_4_;
wire [0:0] cby_1__1__109_left_grid_pin_5_;
wire [0:0] cby_1__1__109_left_grid_pin_6_;
wire [0:0] cby_1__1__109_left_grid_pin_7_;
wire [0:0] cby_1__1__109_left_grid_pin_8_;
wire [0:0] cby_1__1__109_left_grid_pin_9_;
wire [0:0] cby_1__1__109_right_grid_pin_52_;
wire [0:0] cby_1__1__10_ccff_tail;
wire [0:19] cby_1__1__10_chany_bottom_out;
wire [0:19] cby_1__1__10_chany_top_out;
wire [0:0] cby_1__1__10_left_grid_pin_0_;
wire [0:0] cby_1__1__10_left_grid_pin_10_;
wire [0:0] cby_1__1__10_left_grid_pin_11_;
wire [0:0] cby_1__1__10_left_grid_pin_12_;
wire [0:0] cby_1__1__10_left_grid_pin_13_;
wire [0:0] cby_1__1__10_left_grid_pin_14_;
wire [0:0] cby_1__1__10_left_grid_pin_15_;
wire [0:0] cby_1__1__10_left_grid_pin_1_;
wire [0:0] cby_1__1__10_left_grid_pin_2_;
wire [0:0] cby_1__1__10_left_grid_pin_3_;
wire [0:0] cby_1__1__10_left_grid_pin_4_;
wire [0:0] cby_1__1__10_left_grid_pin_5_;
wire [0:0] cby_1__1__10_left_grid_pin_6_;
wire [0:0] cby_1__1__10_left_grid_pin_7_;
wire [0:0] cby_1__1__10_left_grid_pin_8_;
wire [0:0] cby_1__1__10_left_grid_pin_9_;
wire [0:0] cby_1__1__10_right_grid_pin_52_;
wire [0:0] cby_1__1__110_ccff_tail;
wire [0:19] cby_1__1__110_chany_bottom_out;
wire [0:19] cby_1__1__110_chany_top_out;
wire [0:0] cby_1__1__110_left_grid_pin_0_;
wire [0:0] cby_1__1__110_left_grid_pin_10_;
wire [0:0] cby_1__1__110_left_grid_pin_11_;
wire [0:0] cby_1__1__110_left_grid_pin_12_;
wire [0:0] cby_1__1__110_left_grid_pin_13_;
wire [0:0] cby_1__1__110_left_grid_pin_14_;
wire [0:0] cby_1__1__110_left_grid_pin_15_;
wire [0:0] cby_1__1__110_left_grid_pin_1_;
wire [0:0] cby_1__1__110_left_grid_pin_2_;
wire [0:0] cby_1__1__110_left_grid_pin_3_;
wire [0:0] cby_1__1__110_left_grid_pin_4_;
wire [0:0] cby_1__1__110_left_grid_pin_5_;
wire [0:0] cby_1__1__110_left_grid_pin_6_;
wire [0:0] cby_1__1__110_left_grid_pin_7_;
wire [0:0] cby_1__1__110_left_grid_pin_8_;
wire [0:0] cby_1__1__110_left_grid_pin_9_;
wire [0:0] cby_1__1__110_right_grid_pin_52_;
wire [0:0] cby_1__1__111_ccff_tail;
wire [0:19] cby_1__1__111_chany_bottom_out;
wire [0:19] cby_1__1__111_chany_top_out;
wire [0:0] cby_1__1__111_left_grid_pin_0_;
wire [0:0] cby_1__1__111_left_grid_pin_10_;
wire [0:0] cby_1__1__111_left_grid_pin_11_;
wire [0:0] cby_1__1__111_left_grid_pin_12_;
wire [0:0] cby_1__1__111_left_grid_pin_13_;
wire [0:0] cby_1__1__111_left_grid_pin_14_;
wire [0:0] cby_1__1__111_left_grid_pin_15_;
wire [0:0] cby_1__1__111_left_grid_pin_1_;
wire [0:0] cby_1__1__111_left_grid_pin_2_;
wire [0:0] cby_1__1__111_left_grid_pin_3_;
wire [0:0] cby_1__1__111_left_grid_pin_4_;
wire [0:0] cby_1__1__111_left_grid_pin_5_;
wire [0:0] cby_1__1__111_left_grid_pin_6_;
wire [0:0] cby_1__1__111_left_grid_pin_7_;
wire [0:0] cby_1__1__111_left_grid_pin_8_;
wire [0:0] cby_1__1__111_left_grid_pin_9_;
wire [0:0] cby_1__1__111_right_grid_pin_52_;
wire [0:0] cby_1__1__112_ccff_tail;
wire [0:19] cby_1__1__112_chany_bottom_out;
wire [0:19] cby_1__1__112_chany_top_out;
wire [0:0] cby_1__1__112_left_grid_pin_0_;
wire [0:0] cby_1__1__112_left_grid_pin_10_;
wire [0:0] cby_1__1__112_left_grid_pin_11_;
wire [0:0] cby_1__1__112_left_grid_pin_12_;
wire [0:0] cby_1__1__112_left_grid_pin_13_;
wire [0:0] cby_1__1__112_left_grid_pin_14_;
wire [0:0] cby_1__1__112_left_grid_pin_15_;
wire [0:0] cby_1__1__112_left_grid_pin_1_;
wire [0:0] cby_1__1__112_left_grid_pin_2_;
wire [0:0] cby_1__1__112_left_grid_pin_3_;
wire [0:0] cby_1__1__112_left_grid_pin_4_;
wire [0:0] cby_1__1__112_left_grid_pin_5_;
wire [0:0] cby_1__1__112_left_grid_pin_6_;
wire [0:0] cby_1__1__112_left_grid_pin_7_;
wire [0:0] cby_1__1__112_left_grid_pin_8_;
wire [0:0] cby_1__1__112_left_grid_pin_9_;
wire [0:0] cby_1__1__112_right_grid_pin_52_;
wire [0:0] cby_1__1__113_ccff_tail;
wire [0:19] cby_1__1__113_chany_bottom_out;
wire [0:19] cby_1__1__113_chany_top_out;
wire [0:0] cby_1__1__113_left_grid_pin_0_;
wire [0:0] cby_1__1__113_left_grid_pin_10_;
wire [0:0] cby_1__1__113_left_grid_pin_11_;
wire [0:0] cby_1__1__113_left_grid_pin_12_;
wire [0:0] cby_1__1__113_left_grid_pin_13_;
wire [0:0] cby_1__1__113_left_grid_pin_14_;
wire [0:0] cby_1__1__113_left_grid_pin_15_;
wire [0:0] cby_1__1__113_left_grid_pin_1_;
wire [0:0] cby_1__1__113_left_grid_pin_2_;
wire [0:0] cby_1__1__113_left_grid_pin_3_;
wire [0:0] cby_1__1__113_left_grid_pin_4_;
wire [0:0] cby_1__1__113_left_grid_pin_5_;
wire [0:0] cby_1__1__113_left_grid_pin_6_;
wire [0:0] cby_1__1__113_left_grid_pin_7_;
wire [0:0] cby_1__1__113_left_grid_pin_8_;
wire [0:0] cby_1__1__113_left_grid_pin_9_;
wire [0:0] cby_1__1__113_right_grid_pin_52_;
wire [0:0] cby_1__1__114_ccff_tail;
wire [0:19] cby_1__1__114_chany_bottom_out;
wire [0:19] cby_1__1__114_chany_top_out;
wire [0:0] cby_1__1__114_left_grid_pin_0_;
wire [0:0] cby_1__1__114_left_grid_pin_10_;
wire [0:0] cby_1__1__114_left_grid_pin_11_;
wire [0:0] cby_1__1__114_left_grid_pin_12_;
wire [0:0] cby_1__1__114_left_grid_pin_13_;
wire [0:0] cby_1__1__114_left_grid_pin_14_;
wire [0:0] cby_1__1__114_left_grid_pin_15_;
wire [0:0] cby_1__1__114_left_grid_pin_1_;
wire [0:0] cby_1__1__114_left_grid_pin_2_;
wire [0:0] cby_1__1__114_left_grid_pin_3_;
wire [0:0] cby_1__1__114_left_grid_pin_4_;
wire [0:0] cby_1__1__114_left_grid_pin_5_;
wire [0:0] cby_1__1__114_left_grid_pin_6_;
wire [0:0] cby_1__1__114_left_grid_pin_7_;
wire [0:0] cby_1__1__114_left_grid_pin_8_;
wire [0:0] cby_1__1__114_left_grid_pin_9_;
wire [0:0] cby_1__1__114_right_grid_pin_52_;
wire [0:0] cby_1__1__115_ccff_tail;
wire [0:19] cby_1__1__115_chany_bottom_out;
wire [0:19] cby_1__1__115_chany_top_out;
wire [0:0] cby_1__1__115_left_grid_pin_0_;
wire [0:0] cby_1__1__115_left_grid_pin_10_;
wire [0:0] cby_1__1__115_left_grid_pin_11_;
wire [0:0] cby_1__1__115_left_grid_pin_12_;
wire [0:0] cby_1__1__115_left_grid_pin_13_;
wire [0:0] cby_1__1__115_left_grid_pin_14_;
wire [0:0] cby_1__1__115_left_grid_pin_15_;
wire [0:0] cby_1__1__115_left_grid_pin_1_;
wire [0:0] cby_1__1__115_left_grid_pin_2_;
wire [0:0] cby_1__1__115_left_grid_pin_3_;
wire [0:0] cby_1__1__115_left_grid_pin_4_;
wire [0:0] cby_1__1__115_left_grid_pin_5_;
wire [0:0] cby_1__1__115_left_grid_pin_6_;
wire [0:0] cby_1__1__115_left_grid_pin_7_;
wire [0:0] cby_1__1__115_left_grid_pin_8_;
wire [0:0] cby_1__1__115_left_grid_pin_9_;
wire [0:0] cby_1__1__115_right_grid_pin_52_;
wire [0:0] cby_1__1__116_ccff_tail;
wire [0:19] cby_1__1__116_chany_bottom_out;
wire [0:19] cby_1__1__116_chany_top_out;
wire [0:0] cby_1__1__116_left_grid_pin_0_;
wire [0:0] cby_1__1__116_left_grid_pin_10_;
wire [0:0] cby_1__1__116_left_grid_pin_11_;
wire [0:0] cby_1__1__116_left_grid_pin_12_;
wire [0:0] cby_1__1__116_left_grid_pin_13_;
wire [0:0] cby_1__1__116_left_grid_pin_14_;
wire [0:0] cby_1__1__116_left_grid_pin_15_;
wire [0:0] cby_1__1__116_left_grid_pin_1_;
wire [0:0] cby_1__1__116_left_grid_pin_2_;
wire [0:0] cby_1__1__116_left_grid_pin_3_;
wire [0:0] cby_1__1__116_left_grid_pin_4_;
wire [0:0] cby_1__1__116_left_grid_pin_5_;
wire [0:0] cby_1__1__116_left_grid_pin_6_;
wire [0:0] cby_1__1__116_left_grid_pin_7_;
wire [0:0] cby_1__1__116_left_grid_pin_8_;
wire [0:0] cby_1__1__116_left_grid_pin_9_;
wire [0:0] cby_1__1__116_right_grid_pin_52_;
wire [0:0] cby_1__1__117_ccff_tail;
wire [0:19] cby_1__1__117_chany_bottom_out;
wire [0:19] cby_1__1__117_chany_top_out;
wire [0:0] cby_1__1__117_left_grid_pin_0_;
wire [0:0] cby_1__1__117_left_grid_pin_10_;
wire [0:0] cby_1__1__117_left_grid_pin_11_;
wire [0:0] cby_1__1__117_left_grid_pin_12_;
wire [0:0] cby_1__1__117_left_grid_pin_13_;
wire [0:0] cby_1__1__117_left_grid_pin_14_;
wire [0:0] cby_1__1__117_left_grid_pin_15_;
wire [0:0] cby_1__1__117_left_grid_pin_1_;
wire [0:0] cby_1__1__117_left_grid_pin_2_;
wire [0:0] cby_1__1__117_left_grid_pin_3_;
wire [0:0] cby_1__1__117_left_grid_pin_4_;
wire [0:0] cby_1__1__117_left_grid_pin_5_;
wire [0:0] cby_1__1__117_left_grid_pin_6_;
wire [0:0] cby_1__1__117_left_grid_pin_7_;
wire [0:0] cby_1__1__117_left_grid_pin_8_;
wire [0:0] cby_1__1__117_left_grid_pin_9_;
wire [0:0] cby_1__1__117_right_grid_pin_52_;
wire [0:0] cby_1__1__118_ccff_tail;
wire [0:19] cby_1__1__118_chany_bottom_out;
wire [0:19] cby_1__1__118_chany_top_out;
wire [0:0] cby_1__1__118_left_grid_pin_0_;
wire [0:0] cby_1__1__118_left_grid_pin_10_;
wire [0:0] cby_1__1__118_left_grid_pin_11_;
wire [0:0] cby_1__1__118_left_grid_pin_12_;
wire [0:0] cby_1__1__118_left_grid_pin_13_;
wire [0:0] cby_1__1__118_left_grid_pin_14_;
wire [0:0] cby_1__1__118_left_grid_pin_15_;
wire [0:0] cby_1__1__118_left_grid_pin_1_;
wire [0:0] cby_1__1__118_left_grid_pin_2_;
wire [0:0] cby_1__1__118_left_grid_pin_3_;
wire [0:0] cby_1__1__118_left_grid_pin_4_;
wire [0:0] cby_1__1__118_left_grid_pin_5_;
wire [0:0] cby_1__1__118_left_grid_pin_6_;
wire [0:0] cby_1__1__118_left_grid_pin_7_;
wire [0:0] cby_1__1__118_left_grid_pin_8_;
wire [0:0] cby_1__1__118_left_grid_pin_9_;
wire [0:0] cby_1__1__118_right_grid_pin_52_;
wire [0:0] cby_1__1__119_ccff_tail;
wire [0:19] cby_1__1__119_chany_bottom_out;
wire [0:19] cby_1__1__119_chany_top_out;
wire [0:0] cby_1__1__119_left_grid_pin_0_;
wire [0:0] cby_1__1__119_left_grid_pin_10_;
wire [0:0] cby_1__1__119_left_grid_pin_11_;
wire [0:0] cby_1__1__119_left_grid_pin_12_;
wire [0:0] cby_1__1__119_left_grid_pin_13_;
wire [0:0] cby_1__1__119_left_grid_pin_14_;
wire [0:0] cby_1__1__119_left_grid_pin_15_;
wire [0:0] cby_1__1__119_left_grid_pin_1_;
wire [0:0] cby_1__1__119_left_grid_pin_2_;
wire [0:0] cby_1__1__119_left_grid_pin_3_;
wire [0:0] cby_1__1__119_left_grid_pin_4_;
wire [0:0] cby_1__1__119_left_grid_pin_5_;
wire [0:0] cby_1__1__119_left_grid_pin_6_;
wire [0:0] cby_1__1__119_left_grid_pin_7_;
wire [0:0] cby_1__1__119_left_grid_pin_8_;
wire [0:0] cby_1__1__119_left_grid_pin_9_;
wire [0:0] cby_1__1__119_right_grid_pin_52_;
wire [0:0] cby_1__1__11_ccff_tail;
wire [0:19] cby_1__1__11_chany_bottom_out;
wire [0:19] cby_1__1__11_chany_top_out;
wire [0:0] cby_1__1__11_left_grid_pin_0_;
wire [0:0] cby_1__1__11_left_grid_pin_10_;
wire [0:0] cby_1__1__11_left_grid_pin_11_;
wire [0:0] cby_1__1__11_left_grid_pin_12_;
wire [0:0] cby_1__1__11_left_grid_pin_13_;
wire [0:0] cby_1__1__11_left_grid_pin_14_;
wire [0:0] cby_1__1__11_left_grid_pin_15_;
wire [0:0] cby_1__1__11_left_grid_pin_1_;
wire [0:0] cby_1__1__11_left_grid_pin_2_;
wire [0:0] cby_1__1__11_left_grid_pin_3_;
wire [0:0] cby_1__1__11_left_grid_pin_4_;
wire [0:0] cby_1__1__11_left_grid_pin_5_;
wire [0:0] cby_1__1__11_left_grid_pin_6_;
wire [0:0] cby_1__1__11_left_grid_pin_7_;
wire [0:0] cby_1__1__11_left_grid_pin_8_;
wire [0:0] cby_1__1__11_left_grid_pin_9_;
wire [0:0] cby_1__1__11_right_grid_pin_52_;
wire [0:0] cby_1__1__120_ccff_tail;
wire [0:19] cby_1__1__120_chany_bottom_out;
wire [0:19] cby_1__1__120_chany_top_out;
wire [0:0] cby_1__1__120_left_grid_pin_0_;
wire [0:0] cby_1__1__120_left_grid_pin_10_;
wire [0:0] cby_1__1__120_left_grid_pin_11_;
wire [0:0] cby_1__1__120_left_grid_pin_12_;
wire [0:0] cby_1__1__120_left_grid_pin_13_;
wire [0:0] cby_1__1__120_left_grid_pin_14_;
wire [0:0] cby_1__1__120_left_grid_pin_15_;
wire [0:0] cby_1__1__120_left_grid_pin_1_;
wire [0:0] cby_1__1__120_left_grid_pin_2_;
wire [0:0] cby_1__1__120_left_grid_pin_3_;
wire [0:0] cby_1__1__120_left_grid_pin_4_;
wire [0:0] cby_1__1__120_left_grid_pin_5_;
wire [0:0] cby_1__1__120_left_grid_pin_6_;
wire [0:0] cby_1__1__120_left_grid_pin_7_;
wire [0:0] cby_1__1__120_left_grid_pin_8_;
wire [0:0] cby_1__1__120_left_grid_pin_9_;
wire [0:0] cby_1__1__120_right_grid_pin_52_;
wire [0:0] cby_1__1__121_ccff_tail;
wire [0:19] cby_1__1__121_chany_bottom_out;
wire [0:19] cby_1__1__121_chany_top_out;
wire [0:0] cby_1__1__121_left_grid_pin_0_;
wire [0:0] cby_1__1__121_left_grid_pin_10_;
wire [0:0] cby_1__1__121_left_grid_pin_11_;
wire [0:0] cby_1__1__121_left_grid_pin_12_;
wire [0:0] cby_1__1__121_left_grid_pin_13_;
wire [0:0] cby_1__1__121_left_grid_pin_14_;
wire [0:0] cby_1__1__121_left_grid_pin_15_;
wire [0:0] cby_1__1__121_left_grid_pin_1_;
wire [0:0] cby_1__1__121_left_grid_pin_2_;
wire [0:0] cby_1__1__121_left_grid_pin_3_;
wire [0:0] cby_1__1__121_left_grid_pin_4_;
wire [0:0] cby_1__1__121_left_grid_pin_5_;
wire [0:0] cby_1__1__121_left_grid_pin_6_;
wire [0:0] cby_1__1__121_left_grid_pin_7_;
wire [0:0] cby_1__1__121_left_grid_pin_8_;
wire [0:0] cby_1__1__121_left_grid_pin_9_;
wire [0:0] cby_1__1__121_right_grid_pin_52_;
wire [0:0] cby_1__1__122_ccff_tail;
wire [0:19] cby_1__1__122_chany_bottom_out;
wire [0:19] cby_1__1__122_chany_top_out;
wire [0:0] cby_1__1__122_left_grid_pin_0_;
wire [0:0] cby_1__1__122_left_grid_pin_10_;
wire [0:0] cby_1__1__122_left_grid_pin_11_;
wire [0:0] cby_1__1__122_left_grid_pin_12_;
wire [0:0] cby_1__1__122_left_grid_pin_13_;
wire [0:0] cby_1__1__122_left_grid_pin_14_;
wire [0:0] cby_1__1__122_left_grid_pin_15_;
wire [0:0] cby_1__1__122_left_grid_pin_1_;
wire [0:0] cby_1__1__122_left_grid_pin_2_;
wire [0:0] cby_1__1__122_left_grid_pin_3_;
wire [0:0] cby_1__1__122_left_grid_pin_4_;
wire [0:0] cby_1__1__122_left_grid_pin_5_;
wire [0:0] cby_1__1__122_left_grid_pin_6_;
wire [0:0] cby_1__1__122_left_grid_pin_7_;
wire [0:0] cby_1__1__122_left_grid_pin_8_;
wire [0:0] cby_1__1__122_left_grid_pin_9_;
wire [0:0] cby_1__1__122_right_grid_pin_52_;
wire [0:0] cby_1__1__123_ccff_tail;
wire [0:19] cby_1__1__123_chany_bottom_out;
wire [0:19] cby_1__1__123_chany_top_out;
wire [0:0] cby_1__1__123_left_grid_pin_0_;
wire [0:0] cby_1__1__123_left_grid_pin_10_;
wire [0:0] cby_1__1__123_left_grid_pin_11_;
wire [0:0] cby_1__1__123_left_grid_pin_12_;
wire [0:0] cby_1__1__123_left_grid_pin_13_;
wire [0:0] cby_1__1__123_left_grid_pin_14_;
wire [0:0] cby_1__1__123_left_grid_pin_15_;
wire [0:0] cby_1__1__123_left_grid_pin_1_;
wire [0:0] cby_1__1__123_left_grid_pin_2_;
wire [0:0] cby_1__1__123_left_grid_pin_3_;
wire [0:0] cby_1__1__123_left_grid_pin_4_;
wire [0:0] cby_1__1__123_left_grid_pin_5_;
wire [0:0] cby_1__1__123_left_grid_pin_6_;
wire [0:0] cby_1__1__123_left_grid_pin_7_;
wire [0:0] cby_1__1__123_left_grid_pin_8_;
wire [0:0] cby_1__1__123_left_grid_pin_9_;
wire [0:0] cby_1__1__123_right_grid_pin_52_;
wire [0:0] cby_1__1__124_ccff_tail;
wire [0:19] cby_1__1__124_chany_bottom_out;
wire [0:19] cby_1__1__124_chany_top_out;
wire [0:0] cby_1__1__124_left_grid_pin_0_;
wire [0:0] cby_1__1__124_left_grid_pin_10_;
wire [0:0] cby_1__1__124_left_grid_pin_11_;
wire [0:0] cby_1__1__124_left_grid_pin_12_;
wire [0:0] cby_1__1__124_left_grid_pin_13_;
wire [0:0] cby_1__1__124_left_grid_pin_14_;
wire [0:0] cby_1__1__124_left_grid_pin_15_;
wire [0:0] cby_1__1__124_left_grid_pin_1_;
wire [0:0] cby_1__1__124_left_grid_pin_2_;
wire [0:0] cby_1__1__124_left_grid_pin_3_;
wire [0:0] cby_1__1__124_left_grid_pin_4_;
wire [0:0] cby_1__1__124_left_grid_pin_5_;
wire [0:0] cby_1__1__124_left_grid_pin_6_;
wire [0:0] cby_1__1__124_left_grid_pin_7_;
wire [0:0] cby_1__1__124_left_grid_pin_8_;
wire [0:0] cby_1__1__124_left_grid_pin_9_;
wire [0:0] cby_1__1__124_right_grid_pin_52_;
wire [0:0] cby_1__1__125_ccff_tail;
wire [0:19] cby_1__1__125_chany_bottom_out;
wire [0:19] cby_1__1__125_chany_top_out;
wire [0:0] cby_1__1__125_left_grid_pin_0_;
wire [0:0] cby_1__1__125_left_grid_pin_10_;
wire [0:0] cby_1__1__125_left_grid_pin_11_;
wire [0:0] cby_1__1__125_left_grid_pin_12_;
wire [0:0] cby_1__1__125_left_grid_pin_13_;
wire [0:0] cby_1__1__125_left_grid_pin_14_;
wire [0:0] cby_1__1__125_left_grid_pin_15_;
wire [0:0] cby_1__1__125_left_grid_pin_1_;
wire [0:0] cby_1__1__125_left_grid_pin_2_;
wire [0:0] cby_1__1__125_left_grid_pin_3_;
wire [0:0] cby_1__1__125_left_grid_pin_4_;
wire [0:0] cby_1__1__125_left_grid_pin_5_;
wire [0:0] cby_1__1__125_left_grid_pin_6_;
wire [0:0] cby_1__1__125_left_grid_pin_7_;
wire [0:0] cby_1__1__125_left_grid_pin_8_;
wire [0:0] cby_1__1__125_left_grid_pin_9_;
wire [0:0] cby_1__1__125_right_grid_pin_52_;
wire [0:0] cby_1__1__126_ccff_tail;
wire [0:19] cby_1__1__126_chany_bottom_out;
wire [0:19] cby_1__1__126_chany_top_out;
wire [0:0] cby_1__1__126_left_grid_pin_0_;
wire [0:0] cby_1__1__126_left_grid_pin_10_;
wire [0:0] cby_1__1__126_left_grid_pin_11_;
wire [0:0] cby_1__1__126_left_grid_pin_12_;
wire [0:0] cby_1__1__126_left_grid_pin_13_;
wire [0:0] cby_1__1__126_left_grid_pin_14_;
wire [0:0] cby_1__1__126_left_grid_pin_15_;
wire [0:0] cby_1__1__126_left_grid_pin_1_;
wire [0:0] cby_1__1__126_left_grid_pin_2_;
wire [0:0] cby_1__1__126_left_grid_pin_3_;
wire [0:0] cby_1__1__126_left_grid_pin_4_;
wire [0:0] cby_1__1__126_left_grid_pin_5_;
wire [0:0] cby_1__1__126_left_grid_pin_6_;
wire [0:0] cby_1__1__126_left_grid_pin_7_;
wire [0:0] cby_1__1__126_left_grid_pin_8_;
wire [0:0] cby_1__1__126_left_grid_pin_9_;
wire [0:0] cby_1__1__126_right_grid_pin_52_;
wire [0:0] cby_1__1__127_ccff_tail;
wire [0:19] cby_1__1__127_chany_bottom_out;
wire [0:19] cby_1__1__127_chany_top_out;
wire [0:0] cby_1__1__127_left_grid_pin_0_;
wire [0:0] cby_1__1__127_left_grid_pin_10_;
wire [0:0] cby_1__1__127_left_grid_pin_11_;
wire [0:0] cby_1__1__127_left_grid_pin_12_;
wire [0:0] cby_1__1__127_left_grid_pin_13_;
wire [0:0] cby_1__1__127_left_grid_pin_14_;
wire [0:0] cby_1__1__127_left_grid_pin_15_;
wire [0:0] cby_1__1__127_left_grid_pin_1_;
wire [0:0] cby_1__1__127_left_grid_pin_2_;
wire [0:0] cby_1__1__127_left_grid_pin_3_;
wire [0:0] cby_1__1__127_left_grid_pin_4_;
wire [0:0] cby_1__1__127_left_grid_pin_5_;
wire [0:0] cby_1__1__127_left_grid_pin_6_;
wire [0:0] cby_1__1__127_left_grid_pin_7_;
wire [0:0] cby_1__1__127_left_grid_pin_8_;
wire [0:0] cby_1__1__127_left_grid_pin_9_;
wire [0:0] cby_1__1__127_right_grid_pin_52_;
wire [0:0] cby_1__1__128_ccff_tail;
wire [0:19] cby_1__1__128_chany_bottom_out;
wire [0:19] cby_1__1__128_chany_top_out;
wire [0:0] cby_1__1__128_left_grid_pin_0_;
wire [0:0] cby_1__1__128_left_grid_pin_10_;
wire [0:0] cby_1__1__128_left_grid_pin_11_;
wire [0:0] cby_1__1__128_left_grid_pin_12_;
wire [0:0] cby_1__1__128_left_grid_pin_13_;
wire [0:0] cby_1__1__128_left_grid_pin_14_;
wire [0:0] cby_1__1__128_left_grid_pin_15_;
wire [0:0] cby_1__1__128_left_grid_pin_1_;
wire [0:0] cby_1__1__128_left_grid_pin_2_;
wire [0:0] cby_1__1__128_left_grid_pin_3_;
wire [0:0] cby_1__1__128_left_grid_pin_4_;
wire [0:0] cby_1__1__128_left_grid_pin_5_;
wire [0:0] cby_1__1__128_left_grid_pin_6_;
wire [0:0] cby_1__1__128_left_grid_pin_7_;
wire [0:0] cby_1__1__128_left_grid_pin_8_;
wire [0:0] cby_1__1__128_left_grid_pin_9_;
wire [0:0] cby_1__1__128_right_grid_pin_52_;
wire [0:0] cby_1__1__129_ccff_tail;
wire [0:19] cby_1__1__129_chany_bottom_out;
wire [0:19] cby_1__1__129_chany_top_out;
wire [0:0] cby_1__1__129_left_grid_pin_0_;
wire [0:0] cby_1__1__129_left_grid_pin_10_;
wire [0:0] cby_1__1__129_left_grid_pin_11_;
wire [0:0] cby_1__1__129_left_grid_pin_12_;
wire [0:0] cby_1__1__129_left_grid_pin_13_;
wire [0:0] cby_1__1__129_left_grid_pin_14_;
wire [0:0] cby_1__1__129_left_grid_pin_15_;
wire [0:0] cby_1__1__129_left_grid_pin_1_;
wire [0:0] cby_1__1__129_left_grid_pin_2_;
wire [0:0] cby_1__1__129_left_grid_pin_3_;
wire [0:0] cby_1__1__129_left_grid_pin_4_;
wire [0:0] cby_1__1__129_left_grid_pin_5_;
wire [0:0] cby_1__1__129_left_grid_pin_6_;
wire [0:0] cby_1__1__129_left_grid_pin_7_;
wire [0:0] cby_1__1__129_left_grid_pin_8_;
wire [0:0] cby_1__1__129_left_grid_pin_9_;
wire [0:0] cby_1__1__129_right_grid_pin_52_;
wire [0:0] cby_1__1__12_ccff_tail;
wire [0:19] cby_1__1__12_chany_bottom_out;
wire [0:19] cby_1__1__12_chany_top_out;
wire [0:0] cby_1__1__12_left_grid_pin_0_;
wire [0:0] cby_1__1__12_left_grid_pin_10_;
wire [0:0] cby_1__1__12_left_grid_pin_11_;
wire [0:0] cby_1__1__12_left_grid_pin_12_;
wire [0:0] cby_1__1__12_left_grid_pin_13_;
wire [0:0] cby_1__1__12_left_grid_pin_14_;
wire [0:0] cby_1__1__12_left_grid_pin_15_;
wire [0:0] cby_1__1__12_left_grid_pin_1_;
wire [0:0] cby_1__1__12_left_grid_pin_2_;
wire [0:0] cby_1__1__12_left_grid_pin_3_;
wire [0:0] cby_1__1__12_left_grid_pin_4_;
wire [0:0] cby_1__1__12_left_grid_pin_5_;
wire [0:0] cby_1__1__12_left_grid_pin_6_;
wire [0:0] cby_1__1__12_left_grid_pin_7_;
wire [0:0] cby_1__1__12_left_grid_pin_8_;
wire [0:0] cby_1__1__12_left_grid_pin_9_;
wire [0:0] cby_1__1__12_right_grid_pin_52_;
wire [0:0] cby_1__1__130_ccff_tail;
wire [0:19] cby_1__1__130_chany_bottom_out;
wire [0:19] cby_1__1__130_chany_top_out;
wire [0:0] cby_1__1__130_left_grid_pin_0_;
wire [0:0] cby_1__1__130_left_grid_pin_10_;
wire [0:0] cby_1__1__130_left_grid_pin_11_;
wire [0:0] cby_1__1__130_left_grid_pin_12_;
wire [0:0] cby_1__1__130_left_grid_pin_13_;
wire [0:0] cby_1__1__130_left_grid_pin_14_;
wire [0:0] cby_1__1__130_left_grid_pin_15_;
wire [0:0] cby_1__1__130_left_grid_pin_1_;
wire [0:0] cby_1__1__130_left_grid_pin_2_;
wire [0:0] cby_1__1__130_left_grid_pin_3_;
wire [0:0] cby_1__1__130_left_grid_pin_4_;
wire [0:0] cby_1__1__130_left_grid_pin_5_;
wire [0:0] cby_1__1__130_left_grid_pin_6_;
wire [0:0] cby_1__1__130_left_grid_pin_7_;
wire [0:0] cby_1__1__130_left_grid_pin_8_;
wire [0:0] cby_1__1__130_left_grid_pin_9_;
wire [0:0] cby_1__1__130_right_grid_pin_52_;
wire [0:0] cby_1__1__131_ccff_tail;
wire [0:19] cby_1__1__131_chany_bottom_out;
wire [0:19] cby_1__1__131_chany_top_out;
wire [0:0] cby_1__1__131_left_grid_pin_0_;
wire [0:0] cby_1__1__131_left_grid_pin_10_;
wire [0:0] cby_1__1__131_left_grid_pin_11_;
wire [0:0] cby_1__1__131_left_grid_pin_12_;
wire [0:0] cby_1__1__131_left_grid_pin_13_;
wire [0:0] cby_1__1__131_left_grid_pin_14_;
wire [0:0] cby_1__1__131_left_grid_pin_15_;
wire [0:0] cby_1__1__131_left_grid_pin_1_;
wire [0:0] cby_1__1__131_left_grid_pin_2_;
wire [0:0] cby_1__1__131_left_grid_pin_3_;
wire [0:0] cby_1__1__131_left_grid_pin_4_;
wire [0:0] cby_1__1__131_left_grid_pin_5_;
wire [0:0] cby_1__1__131_left_grid_pin_6_;
wire [0:0] cby_1__1__131_left_grid_pin_7_;
wire [0:0] cby_1__1__131_left_grid_pin_8_;
wire [0:0] cby_1__1__131_left_grid_pin_9_;
wire [0:0] cby_1__1__131_right_grid_pin_52_;
wire [0:0] cby_1__1__132_ccff_tail;
wire [0:19] cby_1__1__132_chany_bottom_out;
wire [0:19] cby_1__1__132_chany_top_out;
wire [0:0] cby_1__1__132_left_grid_pin_0_;
wire [0:0] cby_1__1__132_left_grid_pin_10_;
wire [0:0] cby_1__1__132_left_grid_pin_11_;
wire [0:0] cby_1__1__132_left_grid_pin_12_;
wire [0:0] cby_1__1__132_left_grid_pin_13_;
wire [0:0] cby_1__1__132_left_grid_pin_14_;
wire [0:0] cby_1__1__132_left_grid_pin_15_;
wire [0:0] cby_1__1__132_left_grid_pin_1_;
wire [0:0] cby_1__1__132_left_grid_pin_2_;
wire [0:0] cby_1__1__132_left_grid_pin_3_;
wire [0:0] cby_1__1__132_left_grid_pin_4_;
wire [0:0] cby_1__1__132_left_grid_pin_5_;
wire [0:0] cby_1__1__132_left_grid_pin_6_;
wire [0:0] cby_1__1__132_left_grid_pin_7_;
wire [0:0] cby_1__1__132_left_grid_pin_8_;
wire [0:0] cby_1__1__132_left_grid_pin_9_;
wire [0:0] cby_1__1__132_right_grid_pin_52_;
wire [0:0] cby_1__1__133_ccff_tail;
wire [0:19] cby_1__1__133_chany_bottom_out;
wire [0:19] cby_1__1__133_chany_top_out;
wire [0:0] cby_1__1__133_left_grid_pin_0_;
wire [0:0] cby_1__1__133_left_grid_pin_10_;
wire [0:0] cby_1__1__133_left_grid_pin_11_;
wire [0:0] cby_1__1__133_left_grid_pin_12_;
wire [0:0] cby_1__1__133_left_grid_pin_13_;
wire [0:0] cby_1__1__133_left_grid_pin_14_;
wire [0:0] cby_1__1__133_left_grid_pin_15_;
wire [0:0] cby_1__1__133_left_grid_pin_1_;
wire [0:0] cby_1__1__133_left_grid_pin_2_;
wire [0:0] cby_1__1__133_left_grid_pin_3_;
wire [0:0] cby_1__1__133_left_grid_pin_4_;
wire [0:0] cby_1__1__133_left_grid_pin_5_;
wire [0:0] cby_1__1__133_left_grid_pin_6_;
wire [0:0] cby_1__1__133_left_grid_pin_7_;
wire [0:0] cby_1__1__133_left_grid_pin_8_;
wire [0:0] cby_1__1__133_left_grid_pin_9_;
wire [0:0] cby_1__1__133_right_grid_pin_52_;
wire [0:0] cby_1__1__134_ccff_tail;
wire [0:19] cby_1__1__134_chany_bottom_out;
wire [0:19] cby_1__1__134_chany_top_out;
wire [0:0] cby_1__1__134_left_grid_pin_0_;
wire [0:0] cby_1__1__134_left_grid_pin_10_;
wire [0:0] cby_1__1__134_left_grid_pin_11_;
wire [0:0] cby_1__1__134_left_grid_pin_12_;
wire [0:0] cby_1__1__134_left_grid_pin_13_;
wire [0:0] cby_1__1__134_left_grid_pin_14_;
wire [0:0] cby_1__1__134_left_grid_pin_15_;
wire [0:0] cby_1__1__134_left_grid_pin_1_;
wire [0:0] cby_1__1__134_left_grid_pin_2_;
wire [0:0] cby_1__1__134_left_grid_pin_3_;
wire [0:0] cby_1__1__134_left_grid_pin_4_;
wire [0:0] cby_1__1__134_left_grid_pin_5_;
wire [0:0] cby_1__1__134_left_grid_pin_6_;
wire [0:0] cby_1__1__134_left_grid_pin_7_;
wire [0:0] cby_1__1__134_left_grid_pin_8_;
wire [0:0] cby_1__1__134_left_grid_pin_9_;
wire [0:0] cby_1__1__134_right_grid_pin_52_;
wire [0:0] cby_1__1__135_ccff_tail;
wire [0:19] cby_1__1__135_chany_bottom_out;
wire [0:19] cby_1__1__135_chany_top_out;
wire [0:0] cby_1__1__135_left_grid_pin_0_;
wire [0:0] cby_1__1__135_left_grid_pin_10_;
wire [0:0] cby_1__1__135_left_grid_pin_11_;
wire [0:0] cby_1__1__135_left_grid_pin_12_;
wire [0:0] cby_1__1__135_left_grid_pin_13_;
wire [0:0] cby_1__1__135_left_grid_pin_14_;
wire [0:0] cby_1__1__135_left_grid_pin_15_;
wire [0:0] cby_1__1__135_left_grid_pin_1_;
wire [0:0] cby_1__1__135_left_grid_pin_2_;
wire [0:0] cby_1__1__135_left_grid_pin_3_;
wire [0:0] cby_1__1__135_left_grid_pin_4_;
wire [0:0] cby_1__1__135_left_grid_pin_5_;
wire [0:0] cby_1__1__135_left_grid_pin_6_;
wire [0:0] cby_1__1__135_left_grid_pin_7_;
wire [0:0] cby_1__1__135_left_grid_pin_8_;
wire [0:0] cby_1__1__135_left_grid_pin_9_;
wire [0:0] cby_1__1__135_right_grid_pin_52_;
wire [0:0] cby_1__1__136_ccff_tail;
wire [0:19] cby_1__1__136_chany_bottom_out;
wire [0:19] cby_1__1__136_chany_top_out;
wire [0:0] cby_1__1__136_left_grid_pin_0_;
wire [0:0] cby_1__1__136_left_grid_pin_10_;
wire [0:0] cby_1__1__136_left_grid_pin_11_;
wire [0:0] cby_1__1__136_left_grid_pin_12_;
wire [0:0] cby_1__1__136_left_grid_pin_13_;
wire [0:0] cby_1__1__136_left_grid_pin_14_;
wire [0:0] cby_1__1__136_left_grid_pin_15_;
wire [0:0] cby_1__1__136_left_grid_pin_1_;
wire [0:0] cby_1__1__136_left_grid_pin_2_;
wire [0:0] cby_1__1__136_left_grid_pin_3_;
wire [0:0] cby_1__1__136_left_grid_pin_4_;
wire [0:0] cby_1__1__136_left_grid_pin_5_;
wire [0:0] cby_1__1__136_left_grid_pin_6_;
wire [0:0] cby_1__1__136_left_grid_pin_7_;
wire [0:0] cby_1__1__136_left_grid_pin_8_;
wire [0:0] cby_1__1__136_left_grid_pin_9_;
wire [0:0] cby_1__1__136_right_grid_pin_52_;
wire [0:0] cby_1__1__137_ccff_tail;
wire [0:19] cby_1__1__137_chany_bottom_out;
wire [0:19] cby_1__1__137_chany_top_out;
wire [0:0] cby_1__1__137_left_grid_pin_0_;
wire [0:0] cby_1__1__137_left_grid_pin_10_;
wire [0:0] cby_1__1__137_left_grid_pin_11_;
wire [0:0] cby_1__1__137_left_grid_pin_12_;
wire [0:0] cby_1__1__137_left_grid_pin_13_;
wire [0:0] cby_1__1__137_left_grid_pin_14_;
wire [0:0] cby_1__1__137_left_grid_pin_15_;
wire [0:0] cby_1__1__137_left_grid_pin_1_;
wire [0:0] cby_1__1__137_left_grid_pin_2_;
wire [0:0] cby_1__1__137_left_grid_pin_3_;
wire [0:0] cby_1__1__137_left_grid_pin_4_;
wire [0:0] cby_1__1__137_left_grid_pin_5_;
wire [0:0] cby_1__1__137_left_grid_pin_6_;
wire [0:0] cby_1__1__137_left_grid_pin_7_;
wire [0:0] cby_1__1__137_left_grid_pin_8_;
wire [0:0] cby_1__1__137_left_grid_pin_9_;
wire [0:0] cby_1__1__137_right_grid_pin_52_;
wire [0:0] cby_1__1__138_ccff_tail;
wire [0:19] cby_1__1__138_chany_bottom_out;
wire [0:19] cby_1__1__138_chany_top_out;
wire [0:0] cby_1__1__138_left_grid_pin_0_;
wire [0:0] cby_1__1__138_left_grid_pin_10_;
wire [0:0] cby_1__1__138_left_grid_pin_11_;
wire [0:0] cby_1__1__138_left_grid_pin_12_;
wire [0:0] cby_1__1__138_left_grid_pin_13_;
wire [0:0] cby_1__1__138_left_grid_pin_14_;
wire [0:0] cby_1__1__138_left_grid_pin_15_;
wire [0:0] cby_1__1__138_left_grid_pin_1_;
wire [0:0] cby_1__1__138_left_grid_pin_2_;
wire [0:0] cby_1__1__138_left_grid_pin_3_;
wire [0:0] cby_1__1__138_left_grid_pin_4_;
wire [0:0] cby_1__1__138_left_grid_pin_5_;
wire [0:0] cby_1__1__138_left_grid_pin_6_;
wire [0:0] cby_1__1__138_left_grid_pin_7_;
wire [0:0] cby_1__1__138_left_grid_pin_8_;
wire [0:0] cby_1__1__138_left_grid_pin_9_;
wire [0:0] cby_1__1__138_right_grid_pin_52_;
wire [0:0] cby_1__1__139_ccff_tail;
wire [0:19] cby_1__1__139_chany_bottom_out;
wire [0:19] cby_1__1__139_chany_top_out;
wire [0:0] cby_1__1__139_left_grid_pin_0_;
wire [0:0] cby_1__1__139_left_grid_pin_10_;
wire [0:0] cby_1__1__139_left_grid_pin_11_;
wire [0:0] cby_1__1__139_left_grid_pin_12_;
wire [0:0] cby_1__1__139_left_grid_pin_13_;
wire [0:0] cby_1__1__139_left_grid_pin_14_;
wire [0:0] cby_1__1__139_left_grid_pin_15_;
wire [0:0] cby_1__1__139_left_grid_pin_1_;
wire [0:0] cby_1__1__139_left_grid_pin_2_;
wire [0:0] cby_1__1__139_left_grid_pin_3_;
wire [0:0] cby_1__1__139_left_grid_pin_4_;
wire [0:0] cby_1__1__139_left_grid_pin_5_;
wire [0:0] cby_1__1__139_left_grid_pin_6_;
wire [0:0] cby_1__1__139_left_grid_pin_7_;
wire [0:0] cby_1__1__139_left_grid_pin_8_;
wire [0:0] cby_1__1__139_left_grid_pin_9_;
wire [0:0] cby_1__1__139_right_grid_pin_52_;
wire [0:0] cby_1__1__13_ccff_tail;
wire [0:19] cby_1__1__13_chany_bottom_out;
wire [0:19] cby_1__1__13_chany_top_out;
wire [0:0] cby_1__1__13_left_grid_pin_0_;
wire [0:0] cby_1__1__13_left_grid_pin_10_;
wire [0:0] cby_1__1__13_left_grid_pin_11_;
wire [0:0] cby_1__1__13_left_grid_pin_12_;
wire [0:0] cby_1__1__13_left_grid_pin_13_;
wire [0:0] cby_1__1__13_left_grid_pin_14_;
wire [0:0] cby_1__1__13_left_grid_pin_15_;
wire [0:0] cby_1__1__13_left_grid_pin_1_;
wire [0:0] cby_1__1__13_left_grid_pin_2_;
wire [0:0] cby_1__1__13_left_grid_pin_3_;
wire [0:0] cby_1__1__13_left_grid_pin_4_;
wire [0:0] cby_1__1__13_left_grid_pin_5_;
wire [0:0] cby_1__1__13_left_grid_pin_6_;
wire [0:0] cby_1__1__13_left_grid_pin_7_;
wire [0:0] cby_1__1__13_left_grid_pin_8_;
wire [0:0] cby_1__1__13_left_grid_pin_9_;
wire [0:0] cby_1__1__13_right_grid_pin_52_;
wire [0:0] cby_1__1__140_ccff_tail;
wire [0:19] cby_1__1__140_chany_bottom_out;
wire [0:19] cby_1__1__140_chany_top_out;
wire [0:0] cby_1__1__140_left_grid_pin_0_;
wire [0:0] cby_1__1__140_left_grid_pin_10_;
wire [0:0] cby_1__1__140_left_grid_pin_11_;
wire [0:0] cby_1__1__140_left_grid_pin_12_;
wire [0:0] cby_1__1__140_left_grid_pin_13_;
wire [0:0] cby_1__1__140_left_grid_pin_14_;
wire [0:0] cby_1__1__140_left_grid_pin_15_;
wire [0:0] cby_1__1__140_left_grid_pin_1_;
wire [0:0] cby_1__1__140_left_grid_pin_2_;
wire [0:0] cby_1__1__140_left_grid_pin_3_;
wire [0:0] cby_1__1__140_left_grid_pin_4_;
wire [0:0] cby_1__1__140_left_grid_pin_5_;
wire [0:0] cby_1__1__140_left_grid_pin_6_;
wire [0:0] cby_1__1__140_left_grid_pin_7_;
wire [0:0] cby_1__1__140_left_grid_pin_8_;
wire [0:0] cby_1__1__140_left_grid_pin_9_;
wire [0:0] cby_1__1__140_right_grid_pin_52_;
wire [0:0] cby_1__1__141_ccff_tail;
wire [0:19] cby_1__1__141_chany_bottom_out;
wire [0:19] cby_1__1__141_chany_top_out;
wire [0:0] cby_1__1__141_left_grid_pin_0_;
wire [0:0] cby_1__1__141_left_grid_pin_10_;
wire [0:0] cby_1__1__141_left_grid_pin_11_;
wire [0:0] cby_1__1__141_left_grid_pin_12_;
wire [0:0] cby_1__1__141_left_grid_pin_13_;
wire [0:0] cby_1__1__141_left_grid_pin_14_;
wire [0:0] cby_1__1__141_left_grid_pin_15_;
wire [0:0] cby_1__1__141_left_grid_pin_1_;
wire [0:0] cby_1__1__141_left_grid_pin_2_;
wire [0:0] cby_1__1__141_left_grid_pin_3_;
wire [0:0] cby_1__1__141_left_grid_pin_4_;
wire [0:0] cby_1__1__141_left_grid_pin_5_;
wire [0:0] cby_1__1__141_left_grid_pin_6_;
wire [0:0] cby_1__1__141_left_grid_pin_7_;
wire [0:0] cby_1__1__141_left_grid_pin_8_;
wire [0:0] cby_1__1__141_left_grid_pin_9_;
wire [0:0] cby_1__1__141_right_grid_pin_52_;
wire [0:0] cby_1__1__142_ccff_tail;
wire [0:19] cby_1__1__142_chany_bottom_out;
wire [0:19] cby_1__1__142_chany_top_out;
wire [0:0] cby_1__1__142_left_grid_pin_0_;
wire [0:0] cby_1__1__142_left_grid_pin_10_;
wire [0:0] cby_1__1__142_left_grid_pin_11_;
wire [0:0] cby_1__1__142_left_grid_pin_12_;
wire [0:0] cby_1__1__142_left_grid_pin_13_;
wire [0:0] cby_1__1__142_left_grid_pin_14_;
wire [0:0] cby_1__1__142_left_grid_pin_15_;
wire [0:0] cby_1__1__142_left_grid_pin_1_;
wire [0:0] cby_1__1__142_left_grid_pin_2_;
wire [0:0] cby_1__1__142_left_grid_pin_3_;
wire [0:0] cby_1__1__142_left_grid_pin_4_;
wire [0:0] cby_1__1__142_left_grid_pin_5_;
wire [0:0] cby_1__1__142_left_grid_pin_6_;
wire [0:0] cby_1__1__142_left_grid_pin_7_;
wire [0:0] cby_1__1__142_left_grid_pin_8_;
wire [0:0] cby_1__1__142_left_grid_pin_9_;
wire [0:0] cby_1__1__142_right_grid_pin_52_;
wire [0:0] cby_1__1__143_ccff_tail;
wire [0:19] cby_1__1__143_chany_bottom_out;
wire [0:19] cby_1__1__143_chany_top_out;
wire [0:0] cby_1__1__143_left_grid_pin_0_;
wire [0:0] cby_1__1__143_left_grid_pin_10_;
wire [0:0] cby_1__1__143_left_grid_pin_11_;
wire [0:0] cby_1__1__143_left_grid_pin_12_;
wire [0:0] cby_1__1__143_left_grid_pin_13_;
wire [0:0] cby_1__1__143_left_grid_pin_14_;
wire [0:0] cby_1__1__143_left_grid_pin_15_;
wire [0:0] cby_1__1__143_left_grid_pin_1_;
wire [0:0] cby_1__1__143_left_grid_pin_2_;
wire [0:0] cby_1__1__143_left_grid_pin_3_;
wire [0:0] cby_1__1__143_left_grid_pin_4_;
wire [0:0] cby_1__1__143_left_grid_pin_5_;
wire [0:0] cby_1__1__143_left_grid_pin_6_;
wire [0:0] cby_1__1__143_left_grid_pin_7_;
wire [0:0] cby_1__1__143_left_grid_pin_8_;
wire [0:0] cby_1__1__143_left_grid_pin_9_;
wire [0:0] cby_1__1__143_right_grid_pin_52_;
wire [0:0] cby_1__1__14_ccff_tail;
wire [0:19] cby_1__1__14_chany_bottom_out;
wire [0:19] cby_1__1__14_chany_top_out;
wire [0:0] cby_1__1__14_left_grid_pin_0_;
wire [0:0] cby_1__1__14_left_grid_pin_10_;
wire [0:0] cby_1__1__14_left_grid_pin_11_;
wire [0:0] cby_1__1__14_left_grid_pin_12_;
wire [0:0] cby_1__1__14_left_grid_pin_13_;
wire [0:0] cby_1__1__14_left_grid_pin_14_;
wire [0:0] cby_1__1__14_left_grid_pin_15_;
wire [0:0] cby_1__1__14_left_grid_pin_1_;
wire [0:0] cby_1__1__14_left_grid_pin_2_;
wire [0:0] cby_1__1__14_left_grid_pin_3_;
wire [0:0] cby_1__1__14_left_grid_pin_4_;
wire [0:0] cby_1__1__14_left_grid_pin_5_;
wire [0:0] cby_1__1__14_left_grid_pin_6_;
wire [0:0] cby_1__1__14_left_grid_pin_7_;
wire [0:0] cby_1__1__14_left_grid_pin_8_;
wire [0:0] cby_1__1__14_left_grid_pin_9_;
wire [0:0] cby_1__1__14_right_grid_pin_52_;
wire [0:0] cby_1__1__15_ccff_tail;
wire [0:19] cby_1__1__15_chany_bottom_out;
wire [0:19] cby_1__1__15_chany_top_out;
wire [0:0] cby_1__1__15_left_grid_pin_0_;
wire [0:0] cby_1__1__15_left_grid_pin_10_;
wire [0:0] cby_1__1__15_left_grid_pin_11_;
wire [0:0] cby_1__1__15_left_grid_pin_12_;
wire [0:0] cby_1__1__15_left_grid_pin_13_;
wire [0:0] cby_1__1__15_left_grid_pin_14_;
wire [0:0] cby_1__1__15_left_grid_pin_15_;
wire [0:0] cby_1__1__15_left_grid_pin_1_;
wire [0:0] cby_1__1__15_left_grid_pin_2_;
wire [0:0] cby_1__1__15_left_grid_pin_3_;
wire [0:0] cby_1__1__15_left_grid_pin_4_;
wire [0:0] cby_1__1__15_left_grid_pin_5_;
wire [0:0] cby_1__1__15_left_grid_pin_6_;
wire [0:0] cby_1__1__15_left_grid_pin_7_;
wire [0:0] cby_1__1__15_left_grid_pin_8_;
wire [0:0] cby_1__1__15_left_grid_pin_9_;
wire [0:0] cby_1__1__15_right_grid_pin_52_;
wire [0:0] cby_1__1__16_ccff_tail;
wire [0:19] cby_1__1__16_chany_bottom_out;
wire [0:19] cby_1__1__16_chany_top_out;
wire [0:0] cby_1__1__16_left_grid_pin_0_;
wire [0:0] cby_1__1__16_left_grid_pin_10_;
wire [0:0] cby_1__1__16_left_grid_pin_11_;
wire [0:0] cby_1__1__16_left_grid_pin_12_;
wire [0:0] cby_1__1__16_left_grid_pin_13_;
wire [0:0] cby_1__1__16_left_grid_pin_14_;
wire [0:0] cby_1__1__16_left_grid_pin_15_;
wire [0:0] cby_1__1__16_left_grid_pin_1_;
wire [0:0] cby_1__1__16_left_grid_pin_2_;
wire [0:0] cby_1__1__16_left_grid_pin_3_;
wire [0:0] cby_1__1__16_left_grid_pin_4_;
wire [0:0] cby_1__1__16_left_grid_pin_5_;
wire [0:0] cby_1__1__16_left_grid_pin_6_;
wire [0:0] cby_1__1__16_left_grid_pin_7_;
wire [0:0] cby_1__1__16_left_grid_pin_8_;
wire [0:0] cby_1__1__16_left_grid_pin_9_;
wire [0:0] cby_1__1__16_right_grid_pin_52_;
wire [0:0] cby_1__1__17_ccff_tail;
wire [0:19] cby_1__1__17_chany_bottom_out;
wire [0:19] cby_1__1__17_chany_top_out;
wire [0:0] cby_1__1__17_left_grid_pin_0_;
wire [0:0] cby_1__1__17_left_grid_pin_10_;
wire [0:0] cby_1__1__17_left_grid_pin_11_;
wire [0:0] cby_1__1__17_left_grid_pin_12_;
wire [0:0] cby_1__1__17_left_grid_pin_13_;
wire [0:0] cby_1__1__17_left_grid_pin_14_;
wire [0:0] cby_1__1__17_left_grid_pin_15_;
wire [0:0] cby_1__1__17_left_grid_pin_1_;
wire [0:0] cby_1__1__17_left_grid_pin_2_;
wire [0:0] cby_1__1__17_left_grid_pin_3_;
wire [0:0] cby_1__1__17_left_grid_pin_4_;
wire [0:0] cby_1__1__17_left_grid_pin_5_;
wire [0:0] cby_1__1__17_left_grid_pin_6_;
wire [0:0] cby_1__1__17_left_grid_pin_7_;
wire [0:0] cby_1__1__17_left_grid_pin_8_;
wire [0:0] cby_1__1__17_left_grid_pin_9_;
wire [0:0] cby_1__1__17_right_grid_pin_52_;
wire [0:0] cby_1__1__18_ccff_tail;
wire [0:19] cby_1__1__18_chany_bottom_out;
wire [0:19] cby_1__1__18_chany_top_out;
wire [0:0] cby_1__1__18_left_grid_pin_0_;
wire [0:0] cby_1__1__18_left_grid_pin_10_;
wire [0:0] cby_1__1__18_left_grid_pin_11_;
wire [0:0] cby_1__1__18_left_grid_pin_12_;
wire [0:0] cby_1__1__18_left_grid_pin_13_;
wire [0:0] cby_1__1__18_left_grid_pin_14_;
wire [0:0] cby_1__1__18_left_grid_pin_15_;
wire [0:0] cby_1__1__18_left_grid_pin_1_;
wire [0:0] cby_1__1__18_left_grid_pin_2_;
wire [0:0] cby_1__1__18_left_grid_pin_3_;
wire [0:0] cby_1__1__18_left_grid_pin_4_;
wire [0:0] cby_1__1__18_left_grid_pin_5_;
wire [0:0] cby_1__1__18_left_grid_pin_6_;
wire [0:0] cby_1__1__18_left_grid_pin_7_;
wire [0:0] cby_1__1__18_left_grid_pin_8_;
wire [0:0] cby_1__1__18_left_grid_pin_9_;
wire [0:0] cby_1__1__18_right_grid_pin_52_;
wire [0:0] cby_1__1__19_ccff_tail;
wire [0:19] cby_1__1__19_chany_bottom_out;
wire [0:19] cby_1__1__19_chany_top_out;
wire [0:0] cby_1__1__19_left_grid_pin_0_;
wire [0:0] cby_1__1__19_left_grid_pin_10_;
wire [0:0] cby_1__1__19_left_grid_pin_11_;
wire [0:0] cby_1__1__19_left_grid_pin_12_;
wire [0:0] cby_1__1__19_left_grid_pin_13_;
wire [0:0] cby_1__1__19_left_grid_pin_14_;
wire [0:0] cby_1__1__19_left_grid_pin_15_;
wire [0:0] cby_1__1__19_left_grid_pin_1_;
wire [0:0] cby_1__1__19_left_grid_pin_2_;
wire [0:0] cby_1__1__19_left_grid_pin_3_;
wire [0:0] cby_1__1__19_left_grid_pin_4_;
wire [0:0] cby_1__1__19_left_grid_pin_5_;
wire [0:0] cby_1__1__19_left_grid_pin_6_;
wire [0:0] cby_1__1__19_left_grid_pin_7_;
wire [0:0] cby_1__1__19_left_grid_pin_8_;
wire [0:0] cby_1__1__19_left_grid_pin_9_;
wire [0:0] cby_1__1__19_right_grid_pin_52_;
wire [0:0] cby_1__1__1_ccff_tail;
wire [0:19] cby_1__1__1_chany_bottom_out;
wire [0:19] cby_1__1__1_chany_top_out;
wire [0:0] cby_1__1__1_left_grid_pin_0_;
wire [0:0] cby_1__1__1_left_grid_pin_10_;
wire [0:0] cby_1__1__1_left_grid_pin_11_;
wire [0:0] cby_1__1__1_left_grid_pin_12_;
wire [0:0] cby_1__1__1_left_grid_pin_13_;
wire [0:0] cby_1__1__1_left_grid_pin_14_;
wire [0:0] cby_1__1__1_left_grid_pin_15_;
wire [0:0] cby_1__1__1_left_grid_pin_1_;
wire [0:0] cby_1__1__1_left_grid_pin_2_;
wire [0:0] cby_1__1__1_left_grid_pin_3_;
wire [0:0] cby_1__1__1_left_grid_pin_4_;
wire [0:0] cby_1__1__1_left_grid_pin_5_;
wire [0:0] cby_1__1__1_left_grid_pin_6_;
wire [0:0] cby_1__1__1_left_grid_pin_7_;
wire [0:0] cby_1__1__1_left_grid_pin_8_;
wire [0:0] cby_1__1__1_left_grid_pin_9_;
wire [0:0] cby_1__1__1_right_grid_pin_52_;
wire [0:0] cby_1__1__20_ccff_tail;
wire [0:19] cby_1__1__20_chany_bottom_out;
wire [0:19] cby_1__1__20_chany_top_out;
wire [0:0] cby_1__1__20_left_grid_pin_0_;
wire [0:0] cby_1__1__20_left_grid_pin_10_;
wire [0:0] cby_1__1__20_left_grid_pin_11_;
wire [0:0] cby_1__1__20_left_grid_pin_12_;
wire [0:0] cby_1__1__20_left_grid_pin_13_;
wire [0:0] cby_1__1__20_left_grid_pin_14_;
wire [0:0] cby_1__1__20_left_grid_pin_15_;
wire [0:0] cby_1__1__20_left_grid_pin_1_;
wire [0:0] cby_1__1__20_left_grid_pin_2_;
wire [0:0] cby_1__1__20_left_grid_pin_3_;
wire [0:0] cby_1__1__20_left_grid_pin_4_;
wire [0:0] cby_1__1__20_left_grid_pin_5_;
wire [0:0] cby_1__1__20_left_grid_pin_6_;
wire [0:0] cby_1__1__20_left_grid_pin_7_;
wire [0:0] cby_1__1__20_left_grid_pin_8_;
wire [0:0] cby_1__1__20_left_grid_pin_9_;
wire [0:0] cby_1__1__20_right_grid_pin_52_;
wire [0:0] cby_1__1__21_ccff_tail;
wire [0:19] cby_1__1__21_chany_bottom_out;
wire [0:19] cby_1__1__21_chany_top_out;
wire [0:0] cby_1__1__21_left_grid_pin_0_;
wire [0:0] cby_1__1__21_left_grid_pin_10_;
wire [0:0] cby_1__1__21_left_grid_pin_11_;
wire [0:0] cby_1__1__21_left_grid_pin_12_;
wire [0:0] cby_1__1__21_left_grid_pin_13_;
wire [0:0] cby_1__1__21_left_grid_pin_14_;
wire [0:0] cby_1__1__21_left_grid_pin_15_;
wire [0:0] cby_1__1__21_left_grid_pin_1_;
wire [0:0] cby_1__1__21_left_grid_pin_2_;
wire [0:0] cby_1__1__21_left_grid_pin_3_;
wire [0:0] cby_1__1__21_left_grid_pin_4_;
wire [0:0] cby_1__1__21_left_grid_pin_5_;
wire [0:0] cby_1__1__21_left_grid_pin_6_;
wire [0:0] cby_1__1__21_left_grid_pin_7_;
wire [0:0] cby_1__1__21_left_grid_pin_8_;
wire [0:0] cby_1__1__21_left_grid_pin_9_;
wire [0:0] cby_1__1__21_right_grid_pin_52_;
wire [0:0] cby_1__1__22_ccff_tail;
wire [0:19] cby_1__1__22_chany_bottom_out;
wire [0:19] cby_1__1__22_chany_top_out;
wire [0:0] cby_1__1__22_left_grid_pin_0_;
wire [0:0] cby_1__1__22_left_grid_pin_10_;
wire [0:0] cby_1__1__22_left_grid_pin_11_;
wire [0:0] cby_1__1__22_left_grid_pin_12_;
wire [0:0] cby_1__1__22_left_grid_pin_13_;
wire [0:0] cby_1__1__22_left_grid_pin_14_;
wire [0:0] cby_1__1__22_left_grid_pin_15_;
wire [0:0] cby_1__1__22_left_grid_pin_1_;
wire [0:0] cby_1__1__22_left_grid_pin_2_;
wire [0:0] cby_1__1__22_left_grid_pin_3_;
wire [0:0] cby_1__1__22_left_grid_pin_4_;
wire [0:0] cby_1__1__22_left_grid_pin_5_;
wire [0:0] cby_1__1__22_left_grid_pin_6_;
wire [0:0] cby_1__1__22_left_grid_pin_7_;
wire [0:0] cby_1__1__22_left_grid_pin_8_;
wire [0:0] cby_1__1__22_left_grid_pin_9_;
wire [0:0] cby_1__1__22_right_grid_pin_52_;
wire [0:0] cby_1__1__23_ccff_tail;
wire [0:19] cby_1__1__23_chany_bottom_out;
wire [0:19] cby_1__1__23_chany_top_out;
wire [0:0] cby_1__1__23_left_grid_pin_0_;
wire [0:0] cby_1__1__23_left_grid_pin_10_;
wire [0:0] cby_1__1__23_left_grid_pin_11_;
wire [0:0] cby_1__1__23_left_grid_pin_12_;
wire [0:0] cby_1__1__23_left_grid_pin_13_;
wire [0:0] cby_1__1__23_left_grid_pin_14_;
wire [0:0] cby_1__1__23_left_grid_pin_15_;
wire [0:0] cby_1__1__23_left_grid_pin_1_;
wire [0:0] cby_1__1__23_left_grid_pin_2_;
wire [0:0] cby_1__1__23_left_grid_pin_3_;
wire [0:0] cby_1__1__23_left_grid_pin_4_;
wire [0:0] cby_1__1__23_left_grid_pin_5_;
wire [0:0] cby_1__1__23_left_grid_pin_6_;
wire [0:0] cby_1__1__23_left_grid_pin_7_;
wire [0:0] cby_1__1__23_left_grid_pin_8_;
wire [0:0] cby_1__1__23_left_grid_pin_9_;
wire [0:0] cby_1__1__23_right_grid_pin_52_;
wire [0:0] cby_1__1__24_ccff_tail;
wire [0:19] cby_1__1__24_chany_bottom_out;
wire [0:19] cby_1__1__24_chany_top_out;
wire [0:0] cby_1__1__24_left_grid_pin_0_;
wire [0:0] cby_1__1__24_left_grid_pin_10_;
wire [0:0] cby_1__1__24_left_grid_pin_11_;
wire [0:0] cby_1__1__24_left_grid_pin_12_;
wire [0:0] cby_1__1__24_left_grid_pin_13_;
wire [0:0] cby_1__1__24_left_grid_pin_14_;
wire [0:0] cby_1__1__24_left_grid_pin_15_;
wire [0:0] cby_1__1__24_left_grid_pin_1_;
wire [0:0] cby_1__1__24_left_grid_pin_2_;
wire [0:0] cby_1__1__24_left_grid_pin_3_;
wire [0:0] cby_1__1__24_left_grid_pin_4_;
wire [0:0] cby_1__1__24_left_grid_pin_5_;
wire [0:0] cby_1__1__24_left_grid_pin_6_;
wire [0:0] cby_1__1__24_left_grid_pin_7_;
wire [0:0] cby_1__1__24_left_grid_pin_8_;
wire [0:0] cby_1__1__24_left_grid_pin_9_;
wire [0:0] cby_1__1__24_right_grid_pin_52_;
wire [0:0] cby_1__1__25_ccff_tail;
wire [0:19] cby_1__1__25_chany_bottom_out;
wire [0:19] cby_1__1__25_chany_top_out;
wire [0:0] cby_1__1__25_left_grid_pin_0_;
wire [0:0] cby_1__1__25_left_grid_pin_10_;
wire [0:0] cby_1__1__25_left_grid_pin_11_;
wire [0:0] cby_1__1__25_left_grid_pin_12_;
wire [0:0] cby_1__1__25_left_grid_pin_13_;
wire [0:0] cby_1__1__25_left_grid_pin_14_;
wire [0:0] cby_1__1__25_left_grid_pin_15_;
wire [0:0] cby_1__1__25_left_grid_pin_1_;
wire [0:0] cby_1__1__25_left_grid_pin_2_;
wire [0:0] cby_1__1__25_left_grid_pin_3_;
wire [0:0] cby_1__1__25_left_grid_pin_4_;
wire [0:0] cby_1__1__25_left_grid_pin_5_;
wire [0:0] cby_1__1__25_left_grid_pin_6_;
wire [0:0] cby_1__1__25_left_grid_pin_7_;
wire [0:0] cby_1__1__25_left_grid_pin_8_;
wire [0:0] cby_1__1__25_left_grid_pin_9_;
wire [0:0] cby_1__1__25_right_grid_pin_52_;
wire [0:0] cby_1__1__26_ccff_tail;
wire [0:19] cby_1__1__26_chany_bottom_out;
wire [0:19] cby_1__1__26_chany_top_out;
wire [0:0] cby_1__1__26_left_grid_pin_0_;
wire [0:0] cby_1__1__26_left_grid_pin_10_;
wire [0:0] cby_1__1__26_left_grid_pin_11_;
wire [0:0] cby_1__1__26_left_grid_pin_12_;
wire [0:0] cby_1__1__26_left_grid_pin_13_;
wire [0:0] cby_1__1__26_left_grid_pin_14_;
wire [0:0] cby_1__1__26_left_grid_pin_15_;
wire [0:0] cby_1__1__26_left_grid_pin_1_;
wire [0:0] cby_1__1__26_left_grid_pin_2_;
wire [0:0] cby_1__1__26_left_grid_pin_3_;
wire [0:0] cby_1__1__26_left_grid_pin_4_;
wire [0:0] cby_1__1__26_left_grid_pin_5_;
wire [0:0] cby_1__1__26_left_grid_pin_6_;
wire [0:0] cby_1__1__26_left_grid_pin_7_;
wire [0:0] cby_1__1__26_left_grid_pin_8_;
wire [0:0] cby_1__1__26_left_grid_pin_9_;
wire [0:0] cby_1__1__26_right_grid_pin_52_;
wire [0:0] cby_1__1__27_ccff_tail;
wire [0:19] cby_1__1__27_chany_bottom_out;
wire [0:19] cby_1__1__27_chany_top_out;
wire [0:0] cby_1__1__27_left_grid_pin_0_;
wire [0:0] cby_1__1__27_left_grid_pin_10_;
wire [0:0] cby_1__1__27_left_grid_pin_11_;
wire [0:0] cby_1__1__27_left_grid_pin_12_;
wire [0:0] cby_1__1__27_left_grid_pin_13_;
wire [0:0] cby_1__1__27_left_grid_pin_14_;
wire [0:0] cby_1__1__27_left_grid_pin_15_;
wire [0:0] cby_1__1__27_left_grid_pin_1_;
wire [0:0] cby_1__1__27_left_grid_pin_2_;
wire [0:0] cby_1__1__27_left_grid_pin_3_;
wire [0:0] cby_1__1__27_left_grid_pin_4_;
wire [0:0] cby_1__1__27_left_grid_pin_5_;
wire [0:0] cby_1__1__27_left_grid_pin_6_;
wire [0:0] cby_1__1__27_left_grid_pin_7_;
wire [0:0] cby_1__1__27_left_grid_pin_8_;
wire [0:0] cby_1__1__27_left_grid_pin_9_;
wire [0:0] cby_1__1__27_right_grid_pin_52_;
wire [0:0] cby_1__1__28_ccff_tail;
wire [0:19] cby_1__1__28_chany_bottom_out;
wire [0:19] cby_1__1__28_chany_top_out;
wire [0:0] cby_1__1__28_left_grid_pin_0_;
wire [0:0] cby_1__1__28_left_grid_pin_10_;
wire [0:0] cby_1__1__28_left_grid_pin_11_;
wire [0:0] cby_1__1__28_left_grid_pin_12_;
wire [0:0] cby_1__1__28_left_grid_pin_13_;
wire [0:0] cby_1__1__28_left_grid_pin_14_;
wire [0:0] cby_1__1__28_left_grid_pin_15_;
wire [0:0] cby_1__1__28_left_grid_pin_1_;
wire [0:0] cby_1__1__28_left_grid_pin_2_;
wire [0:0] cby_1__1__28_left_grid_pin_3_;
wire [0:0] cby_1__1__28_left_grid_pin_4_;
wire [0:0] cby_1__1__28_left_grid_pin_5_;
wire [0:0] cby_1__1__28_left_grid_pin_6_;
wire [0:0] cby_1__1__28_left_grid_pin_7_;
wire [0:0] cby_1__1__28_left_grid_pin_8_;
wire [0:0] cby_1__1__28_left_grid_pin_9_;
wire [0:0] cby_1__1__28_right_grid_pin_52_;
wire [0:0] cby_1__1__29_ccff_tail;
wire [0:19] cby_1__1__29_chany_bottom_out;
wire [0:19] cby_1__1__29_chany_top_out;
wire [0:0] cby_1__1__29_left_grid_pin_0_;
wire [0:0] cby_1__1__29_left_grid_pin_10_;
wire [0:0] cby_1__1__29_left_grid_pin_11_;
wire [0:0] cby_1__1__29_left_grid_pin_12_;
wire [0:0] cby_1__1__29_left_grid_pin_13_;
wire [0:0] cby_1__1__29_left_grid_pin_14_;
wire [0:0] cby_1__1__29_left_grid_pin_15_;
wire [0:0] cby_1__1__29_left_grid_pin_1_;
wire [0:0] cby_1__1__29_left_grid_pin_2_;
wire [0:0] cby_1__1__29_left_grid_pin_3_;
wire [0:0] cby_1__1__29_left_grid_pin_4_;
wire [0:0] cby_1__1__29_left_grid_pin_5_;
wire [0:0] cby_1__1__29_left_grid_pin_6_;
wire [0:0] cby_1__1__29_left_grid_pin_7_;
wire [0:0] cby_1__1__29_left_grid_pin_8_;
wire [0:0] cby_1__1__29_left_grid_pin_9_;
wire [0:0] cby_1__1__29_right_grid_pin_52_;
wire [0:0] cby_1__1__2_ccff_tail;
wire [0:19] cby_1__1__2_chany_bottom_out;
wire [0:19] cby_1__1__2_chany_top_out;
wire [0:0] cby_1__1__2_left_grid_pin_0_;
wire [0:0] cby_1__1__2_left_grid_pin_10_;
wire [0:0] cby_1__1__2_left_grid_pin_11_;
wire [0:0] cby_1__1__2_left_grid_pin_12_;
wire [0:0] cby_1__1__2_left_grid_pin_13_;
wire [0:0] cby_1__1__2_left_grid_pin_14_;
wire [0:0] cby_1__1__2_left_grid_pin_15_;
wire [0:0] cby_1__1__2_left_grid_pin_1_;
wire [0:0] cby_1__1__2_left_grid_pin_2_;
wire [0:0] cby_1__1__2_left_grid_pin_3_;
wire [0:0] cby_1__1__2_left_grid_pin_4_;
wire [0:0] cby_1__1__2_left_grid_pin_5_;
wire [0:0] cby_1__1__2_left_grid_pin_6_;
wire [0:0] cby_1__1__2_left_grid_pin_7_;
wire [0:0] cby_1__1__2_left_grid_pin_8_;
wire [0:0] cby_1__1__2_left_grid_pin_9_;
wire [0:0] cby_1__1__2_right_grid_pin_52_;
wire [0:0] cby_1__1__30_ccff_tail;
wire [0:19] cby_1__1__30_chany_bottom_out;
wire [0:19] cby_1__1__30_chany_top_out;
wire [0:0] cby_1__1__30_left_grid_pin_0_;
wire [0:0] cby_1__1__30_left_grid_pin_10_;
wire [0:0] cby_1__1__30_left_grid_pin_11_;
wire [0:0] cby_1__1__30_left_grid_pin_12_;
wire [0:0] cby_1__1__30_left_grid_pin_13_;
wire [0:0] cby_1__1__30_left_grid_pin_14_;
wire [0:0] cby_1__1__30_left_grid_pin_15_;
wire [0:0] cby_1__1__30_left_grid_pin_1_;
wire [0:0] cby_1__1__30_left_grid_pin_2_;
wire [0:0] cby_1__1__30_left_grid_pin_3_;
wire [0:0] cby_1__1__30_left_grid_pin_4_;
wire [0:0] cby_1__1__30_left_grid_pin_5_;
wire [0:0] cby_1__1__30_left_grid_pin_6_;
wire [0:0] cby_1__1__30_left_grid_pin_7_;
wire [0:0] cby_1__1__30_left_grid_pin_8_;
wire [0:0] cby_1__1__30_left_grid_pin_9_;
wire [0:0] cby_1__1__30_right_grid_pin_52_;
wire [0:0] cby_1__1__31_ccff_tail;
wire [0:19] cby_1__1__31_chany_bottom_out;
wire [0:19] cby_1__1__31_chany_top_out;
wire [0:0] cby_1__1__31_left_grid_pin_0_;
wire [0:0] cby_1__1__31_left_grid_pin_10_;
wire [0:0] cby_1__1__31_left_grid_pin_11_;
wire [0:0] cby_1__1__31_left_grid_pin_12_;
wire [0:0] cby_1__1__31_left_grid_pin_13_;
wire [0:0] cby_1__1__31_left_grid_pin_14_;
wire [0:0] cby_1__1__31_left_grid_pin_15_;
wire [0:0] cby_1__1__31_left_grid_pin_1_;
wire [0:0] cby_1__1__31_left_grid_pin_2_;
wire [0:0] cby_1__1__31_left_grid_pin_3_;
wire [0:0] cby_1__1__31_left_grid_pin_4_;
wire [0:0] cby_1__1__31_left_grid_pin_5_;
wire [0:0] cby_1__1__31_left_grid_pin_6_;
wire [0:0] cby_1__1__31_left_grid_pin_7_;
wire [0:0] cby_1__1__31_left_grid_pin_8_;
wire [0:0] cby_1__1__31_left_grid_pin_9_;
wire [0:0] cby_1__1__31_right_grid_pin_52_;
wire [0:0] cby_1__1__32_ccff_tail;
wire [0:19] cby_1__1__32_chany_bottom_out;
wire [0:19] cby_1__1__32_chany_top_out;
wire [0:0] cby_1__1__32_left_grid_pin_0_;
wire [0:0] cby_1__1__32_left_grid_pin_10_;
wire [0:0] cby_1__1__32_left_grid_pin_11_;
wire [0:0] cby_1__1__32_left_grid_pin_12_;
wire [0:0] cby_1__1__32_left_grid_pin_13_;
wire [0:0] cby_1__1__32_left_grid_pin_14_;
wire [0:0] cby_1__1__32_left_grid_pin_15_;
wire [0:0] cby_1__1__32_left_grid_pin_1_;
wire [0:0] cby_1__1__32_left_grid_pin_2_;
wire [0:0] cby_1__1__32_left_grid_pin_3_;
wire [0:0] cby_1__1__32_left_grid_pin_4_;
wire [0:0] cby_1__1__32_left_grid_pin_5_;
wire [0:0] cby_1__1__32_left_grid_pin_6_;
wire [0:0] cby_1__1__32_left_grid_pin_7_;
wire [0:0] cby_1__1__32_left_grid_pin_8_;
wire [0:0] cby_1__1__32_left_grid_pin_9_;
wire [0:0] cby_1__1__32_right_grid_pin_52_;
wire [0:0] cby_1__1__33_ccff_tail;
wire [0:19] cby_1__1__33_chany_bottom_out;
wire [0:19] cby_1__1__33_chany_top_out;
wire [0:0] cby_1__1__33_left_grid_pin_0_;
wire [0:0] cby_1__1__33_left_grid_pin_10_;
wire [0:0] cby_1__1__33_left_grid_pin_11_;
wire [0:0] cby_1__1__33_left_grid_pin_12_;
wire [0:0] cby_1__1__33_left_grid_pin_13_;
wire [0:0] cby_1__1__33_left_grid_pin_14_;
wire [0:0] cby_1__1__33_left_grid_pin_15_;
wire [0:0] cby_1__1__33_left_grid_pin_1_;
wire [0:0] cby_1__1__33_left_grid_pin_2_;
wire [0:0] cby_1__1__33_left_grid_pin_3_;
wire [0:0] cby_1__1__33_left_grid_pin_4_;
wire [0:0] cby_1__1__33_left_grid_pin_5_;
wire [0:0] cby_1__1__33_left_grid_pin_6_;
wire [0:0] cby_1__1__33_left_grid_pin_7_;
wire [0:0] cby_1__1__33_left_grid_pin_8_;
wire [0:0] cby_1__1__33_left_grid_pin_9_;
wire [0:0] cby_1__1__33_right_grid_pin_52_;
wire [0:0] cby_1__1__34_ccff_tail;
wire [0:19] cby_1__1__34_chany_bottom_out;
wire [0:19] cby_1__1__34_chany_top_out;
wire [0:0] cby_1__1__34_left_grid_pin_0_;
wire [0:0] cby_1__1__34_left_grid_pin_10_;
wire [0:0] cby_1__1__34_left_grid_pin_11_;
wire [0:0] cby_1__1__34_left_grid_pin_12_;
wire [0:0] cby_1__1__34_left_grid_pin_13_;
wire [0:0] cby_1__1__34_left_grid_pin_14_;
wire [0:0] cby_1__1__34_left_grid_pin_15_;
wire [0:0] cby_1__1__34_left_grid_pin_1_;
wire [0:0] cby_1__1__34_left_grid_pin_2_;
wire [0:0] cby_1__1__34_left_grid_pin_3_;
wire [0:0] cby_1__1__34_left_grid_pin_4_;
wire [0:0] cby_1__1__34_left_grid_pin_5_;
wire [0:0] cby_1__1__34_left_grid_pin_6_;
wire [0:0] cby_1__1__34_left_grid_pin_7_;
wire [0:0] cby_1__1__34_left_grid_pin_8_;
wire [0:0] cby_1__1__34_left_grid_pin_9_;
wire [0:0] cby_1__1__34_right_grid_pin_52_;
wire [0:0] cby_1__1__35_ccff_tail;
wire [0:19] cby_1__1__35_chany_bottom_out;
wire [0:19] cby_1__1__35_chany_top_out;
wire [0:0] cby_1__1__35_left_grid_pin_0_;
wire [0:0] cby_1__1__35_left_grid_pin_10_;
wire [0:0] cby_1__1__35_left_grid_pin_11_;
wire [0:0] cby_1__1__35_left_grid_pin_12_;
wire [0:0] cby_1__1__35_left_grid_pin_13_;
wire [0:0] cby_1__1__35_left_grid_pin_14_;
wire [0:0] cby_1__1__35_left_grid_pin_15_;
wire [0:0] cby_1__1__35_left_grid_pin_1_;
wire [0:0] cby_1__1__35_left_grid_pin_2_;
wire [0:0] cby_1__1__35_left_grid_pin_3_;
wire [0:0] cby_1__1__35_left_grid_pin_4_;
wire [0:0] cby_1__1__35_left_grid_pin_5_;
wire [0:0] cby_1__1__35_left_grid_pin_6_;
wire [0:0] cby_1__1__35_left_grid_pin_7_;
wire [0:0] cby_1__1__35_left_grid_pin_8_;
wire [0:0] cby_1__1__35_left_grid_pin_9_;
wire [0:0] cby_1__1__35_right_grid_pin_52_;
wire [0:0] cby_1__1__36_ccff_tail;
wire [0:19] cby_1__1__36_chany_bottom_out;
wire [0:19] cby_1__1__36_chany_top_out;
wire [0:0] cby_1__1__36_left_grid_pin_0_;
wire [0:0] cby_1__1__36_left_grid_pin_10_;
wire [0:0] cby_1__1__36_left_grid_pin_11_;
wire [0:0] cby_1__1__36_left_grid_pin_12_;
wire [0:0] cby_1__1__36_left_grid_pin_13_;
wire [0:0] cby_1__1__36_left_grid_pin_14_;
wire [0:0] cby_1__1__36_left_grid_pin_15_;
wire [0:0] cby_1__1__36_left_grid_pin_1_;
wire [0:0] cby_1__1__36_left_grid_pin_2_;
wire [0:0] cby_1__1__36_left_grid_pin_3_;
wire [0:0] cby_1__1__36_left_grid_pin_4_;
wire [0:0] cby_1__1__36_left_grid_pin_5_;
wire [0:0] cby_1__1__36_left_grid_pin_6_;
wire [0:0] cby_1__1__36_left_grid_pin_7_;
wire [0:0] cby_1__1__36_left_grid_pin_8_;
wire [0:0] cby_1__1__36_left_grid_pin_9_;
wire [0:0] cby_1__1__36_right_grid_pin_52_;
wire [0:0] cby_1__1__37_ccff_tail;
wire [0:19] cby_1__1__37_chany_bottom_out;
wire [0:19] cby_1__1__37_chany_top_out;
wire [0:0] cby_1__1__37_left_grid_pin_0_;
wire [0:0] cby_1__1__37_left_grid_pin_10_;
wire [0:0] cby_1__1__37_left_grid_pin_11_;
wire [0:0] cby_1__1__37_left_grid_pin_12_;
wire [0:0] cby_1__1__37_left_grid_pin_13_;
wire [0:0] cby_1__1__37_left_grid_pin_14_;
wire [0:0] cby_1__1__37_left_grid_pin_15_;
wire [0:0] cby_1__1__37_left_grid_pin_1_;
wire [0:0] cby_1__1__37_left_grid_pin_2_;
wire [0:0] cby_1__1__37_left_grid_pin_3_;
wire [0:0] cby_1__1__37_left_grid_pin_4_;
wire [0:0] cby_1__1__37_left_grid_pin_5_;
wire [0:0] cby_1__1__37_left_grid_pin_6_;
wire [0:0] cby_1__1__37_left_grid_pin_7_;
wire [0:0] cby_1__1__37_left_grid_pin_8_;
wire [0:0] cby_1__1__37_left_grid_pin_9_;
wire [0:0] cby_1__1__37_right_grid_pin_52_;
wire [0:0] cby_1__1__38_ccff_tail;
wire [0:19] cby_1__1__38_chany_bottom_out;
wire [0:19] cby_1__1__38_chany_top_out;
wire [0:0] cby_1__1__38_left_grid_pin_0_;
wire [0:0] cby_1__1__38_left_grid_pin_10_;
wire [0:0] cby_1__1__38_left_grid_pin_11_;
wire [0:0] cby_1__1__38_left_grid_pin_12_;
wire [0:0] cby_1__1__38_left_grid_pin_13_;
wire [0:0] cby_1__1__38_left_grid_pin_14_;
wire [0:0] cby_1__1__38_left_grid_pin_15_;
wire [0:0] cby_1__1__38_left_grid_pin_1_;
wire [0:0] cby_1__1__38_left_grid_pin_2_;
wire [0:0] cby_1__1__38_left_grid_pin_3_;
wire [0:0] cby_1__1__38_left_grid_pin_4_;
wire [0:0] cby_1__1__38_left_grid_pin_5_;
wire [0:0] cby_1__1__38_left_grid_pin_6_;
wire [0:0] cby_1__1__38_left_grid_pin_7_;
wire [0:0] cby_1__1__38_left_grid_pin_8_;
wire [0:0] cby_1__1__38_left_grid_pin_9_;
wire [0:0] cby_1__1__38_right_grid_pin_52_;
wire [0:0] cby_1__1__39_ccff_tail;
wire [0:19] cby_1__1__39_chany_bottom_out;
wire [0:19] cby_1__1__39_chany_top_out;
wire [0:0] cby_1__1__39_left_grid_pin_0_;
wire [0:0] cby_1__1__39_left_grid_pin_10_;
wire [0:0] cby_1__1__39_left_grid_pin_11_;
wire [0:0] cby_1__1__39_left_grid_pin_12_;
wire [0:0] cby_1__1__39_left_grid_pin_13_;
wire [0:0] cby_1__1__39_left_grid_pin_14_;
wire [0:0] cby_1__1__39_left_grid_pin_15_;
wire [0:0] cby_1__1__39_left_grid_pin_1_;
wire [0:0] cby_1__1__39_left_grid_pin_2_;
wire [0:0] cby_1__1__39_left_grid_pin_3_;
wire [0:0] cby_1__1__39_left_grid_pin_4_;
wire [0:0] cby_1__1__39_left_grid_pin_5_;
wire [0:0] cby_1__1__39_left_grid_pin_6_;
wire [0:0] cby_1__1__39_left_grid_pin_7_;
wire [0:0] cby_1__1__39_left_grid_pin_8_;
wire [0:0] cby_1__1__39_left_grid_pin_9_;
wire [0:0] cby_1__1__39_right_grid_pin_52_;
wire [0:0] cby_1__1__3_ccff_tail;
wire [0:19] cby_1__1__3_chany_bottom_out;
wire [0:19] cby_1__1__3_chany_top_out;
wire [0:0] cby_1__1__3_left_grid_pin_0_;
wire [0:0] cby_1__1__3_left_grid_pin_10_;
wire [0:0] cby_1__1__3_left_grid_pin_11_;
wire [0:0] cby_1__1__3_left_grid_pin_12_;
wire [0:0] cby_1__1__3_left_grid_pin_13_;
wire [0:0] cby_1__1__3_left_grid_pin_14_;
wire [0:0] cby_1__1__3_left_grid_pin_15_;
wire [0:0] cby_1__1__3_left_grid_pin_1_;
wire [0:0] cby_1__1__3_left_grid_pin_2_;
wire [0:0] cby_1__1__3_left_grid_pin_3_;
wire [0:0] cby_1__1__3_left_grid_pin_4_;
wire [0:0] cby_1__1__3_left_grid_pin_5_;
wire [0:0] cby_1__1__3_left_grid_pin_6_;
wire [0:0] cby_1__1__3_left_grid_pin_7_;
wire [0:0] cby_1__1__3_left_grid_pin_8_;
wire [0:0] cby_1__1__3_left_grid_pin_9_;
wire [0:0] cby_1__1__3_right_grid_pin_52_;
wire [0:0] cby_1__1__40_ccff_tail;
wire [0:19] cby_1__1__40_chany_bottom_out;
wire [0:19] cby_1__1__40_chany_top_out;
wire [0:0] cby_1__1__40_left_grid_pin_0_;
wire [0:0] cby_1__1__40_left_grid_pin_10_;
wire [0:0] cby_1__1__40_left_grid_pin_11_;
wire [0:0] cby_1__1__40_left_grid_pin_12_;
wire [0:0] cby_1__1__40_left_grid_pin_13_;
wire [0:0] cby_1__1__40_left_grid_pin_14_;
wire [0:0] cby_1__1__40_left_grid_pin_15_;
wire [0:0] cby_1__1__40_left_grid_pin_1_;
wire [0:0] cby_1__1__40_left_grid_pin_2_;
wire [0:0] cby_1__1__40_left_grid_pin_3_;
wire [0:0] cby_1__1__40_left_grid_pin_4_;
wire [0:0] cby_1__1__40_left_grid_pin_5_;
wire [0:0] cby_1__1__40_left_grid_pin_6_;
wire [0:0] cby_1__1__40_left_grid_pin_7_;
wire [0:0] cby_1__1__40_left_grid_pin_8_;
wire [0:0] cby_1__1__40_left_grid_pin_9_;
wire [0:0] cby_1__1__40_right_grid_pin_52_;
wire [0:0] cby_1__1__41_ccff_tail;
wire [0:19] cby_1__1__41_chany_bottom_out;
wire [0:19] cby_1__1__41_chany_top_out;
wire [0:0] cby_1__1__41_left_grid_pin_0_;
wire [0:0] cby_1__1__41_left_grid_pin_10_;
wire [0:0] cby_1__1__41_left_grid_pin_11_;
wire [0:0] cby_1__1__41_left_grid_pin_12_;
wire [0:0] cby_1__1__41_left_grid_pin_13_;
wire [0:0] cby_1__1__41_left_grid_pin_14_;
wire [0:0] cby_1__1__41_left_grid_pin_15_;
wire [0:0] cby_1__1__41_left_grid_pin_1_;
wire [0:0] cby_1__1__41_left_grid_pin_2_;
wire [0:0] cby_1__1__41_left_grid_pin_3_;
wire [0:0] cby_1__1__41_left_grid_pin_4_;
wire [0:0] cby_1__1__41_left_grid_pin_5_;
wire [0:0] cby_1__1__41_left_grid_pin_6_;
wire [0:0] cby_1__1__41_left_grid_pin_7_;
wire [0:0] cby_1__1__41_left_grid_pin_8_;
wire [0:0] cby_1__1__41_left_grid_pin_9_;
wire [0:0] cby_1__1__41_right_grid_pin_52_;
wire [0:0] cby_1__1__42_ccff_tail;
wire [0:19] cby_1__1__42_chany_bottom_out;
wire [0:19] cby_1__1__42_chany_top_out;
wire [0:0] cby_1__1__42_left_grid_pin_0_;
wire [0:0] cby_1__1__42_left_grid_pin_10_;
wire [0:0] cby_1__1__42_left_grid_pin_11_;
wire [0:0] cby_1__1__42_left_grid_pin_12_;
wire [0:0] cby_1__1__42_left_grid_pin_13_;
wire [0:0] cby_1__1__42_left_grid_pin_14_;
wire [0:0] cby_1__1__42_left_grid_pin_15_;
wire [0:0] cby_1__1__42_left_grid_pin_1_;
wire [0:0] cby_1__1__42_left_grid_pin_2_;
wire [0:0] cby_1__1__42_left_grid_pin_3_;
wire [0:0] cby_1__1__42_left_grid_pin_4_;
wire [0:0] cby_1__1__42_left_grid_pin_5_;
wire [0:0] cby_1__1__42_left_grid_pin_6_;
wire [0:0] cby_1__1__42_left_grid_pin_7_;
wire [0:0] cby_1__1__42_left_grid_pin_8_;
wire [0:0] cby_1__1__42_left_grid_pin_9_;
wire [0:0] cby_1__1__42_right_grid_pin_52_;
wire [0:0] cby_1__1__43_ccff_tail;
wire [0:19] cby_1__1__43_chany_bottom_out;
wire [0:19] cby_1__1__43_chany_top_out;
wire [0:0] cby_1__1__43_left_grid_pin_0_;
wire [0:0] cby_1__1__43_left_grid_pin_10_;
wire [0:0] cby_1__1__43_left_grid_pin_11_;
wire [0:0] cby_1__1__43_left_grid_pin_12_;
wire [0:0] cby_1__1__43_left_grid_pin_13_;
wire [0:0] cby_1__1__43_left_grid_pin_14_;
wire [0:0] cby_1__1__43_left_grid_pin_15_;
wire [0:0] cby_1__1__43_left_grid_pin_1_;
wire [0:0] cby_1__1__43_left_grid_pin_2_;
wire [0:0] cby_1__1__43_left_grid_pin_3_;
wire [0:0] cby_1__1__43_left_grid_pin_4_;
wire [0:0] cby_1__1__43_left_grid_pin_5_;
wire [0:0] cby_1__1__43_left_grid_pin_6_;
wire [0:0] cby_1__1__43_left_grid_pin_7_;
wire [0:0] cby_1__1__43_left_grid_pin_8_;
wire [0:0] cby_1__1__43_left_grid_pin_9_;
wire [0:0] cby_1__1__43_right_grid_pin_52_;
wire [0:0] cby_1__1__44_ccff_tail;
wire [0:19] cby_1__1__44_chany_bottom_out;
wire [0:19] cby_1__1__44_chany_top_out;
wire [0:0] cby_1__1__44_left_grid_pin_0_;
wire [0:0] cby_1__1__44_left_grid_pin_10_;
wire [0:0] cby_1__1__44_left_grid_pin_11_;
wire [0:0] cby_1__1__44_left_grid_pin_12_;
wire [0:0] cby_1__1__44_left_grid_pin_13_;
wire [0:0] cby_1__1__44_left_grid_pin_14_;
wire [0:0] cby_1__1__44_left_grid_pin_15_;
wire [0:0] cby_1__1__44_left_grid_pin_1_;
wire [0:0] cby_1__1__44_left_grid_pin_2_;
wire [0:0] cby_1__1__44_left_grid_pin_3_;
wire [0:0] cby_1__1__44_left_grid_pin_4_;
wire [0:0] cby_1__1__44_left_grid_pin_5_;
wire [0:0] cby_1__1__44_left_grid_pin_6_;
wire [0:0] cby_1__1__44_left_grid_pin_7_;
wire [0:0] cby_1__1__44_left_grid_pin_8_;
wire [0:0] cby_1__1__44_left_grid_pin_9_;
wire [0:0] cby_1__1__44_right_grid_pin_52_;
wire [0:0] cby_1__1__45_ccff_tail;
wire [0:19] cby_1__1__45_chany_bottom_out;
wire [0:19] cby_1__1__45_chany_top_out;
wire [0:0] cby_1__1__45_left_grid_pin_0_;
wire [0:0] cby_1__1__45_left_grid_pin_10_;
wire [0:0] cby_1__1__45_left_grid_pin_11_;
wire [0:0] cby_1__1__45_left_grid_pin_12_;
wire [0:0] cby_1__1__45_left_grid_pin_13_;
wire [0:0] cby_1__1__45_left_grid_pin_14_;
wire [0:0] cby_1__1__45_left_grid_pin_15_;
wire [0:0] cby_1__1__45_left_grid_pin_1_;
wire [0:0] cby_1__1__45_left_grid_pin_2_;
wire [0:0] cby_1__1__45_left_grid_pin_3_;
wire [0:0] cby_1__1__45_left_grid_pin_4_;
wire [0:0] cby_1__1__45_left_grid_pin_5_;
wire [0:0] cby_1__1__45_left_grid_pin_6_;
wire [0:0] cby_1__1__45_left_grid_pin_7_;
wire [0:0] cby_1__1__45_left_grid_pin_8_;
wire [0:0] cby_1__1__45_left_grid_pin_9_;
wire [0:0] cby_1__1__45_right_grid_pin_52_;
wire [0:0] cby_1__1__46_ccff_tail;
wire [0:19] cby_1__1__46_chany_bottom_out;
wire [0:19] cby_1__1__46_chany_top_out;
wire [0:0] cby_1__1__46_left_grid_pin_0_;
wire [0:0] cby_1__1__46_left_grid_pin_10_;
wire [0:0] cby_1__1__46_left_grid_pin_11_;
wire [0:0] cby_1__1__46_left_grid_pin_12_;
wire [0:0] cby_1__1__46_left_grid_pin_13_;
wire [0:0] cby_1__1__46_left_grid_pin_14_;
wire [0:0] cby_1__1__46_left_grid_pin_15_;
wire [0:0] cby_1__1__46_left_grid_pin_1_;
wire [0:0] cby_1__1__46_left_grid_pin_2_;
wire [0:0] cby_1__1__46_left_grid_pin_3_;
wire [0:0] cby_1__1__46_left_grid_pin_4_;
wire [0:0] cby_1__1__46_left_grid_pin_5_;
wire [0:0] cby_1__1__46_left_grid_pin_6_;
wire [0:0] cby_1__1__46_left_grid_pin_7_;
wire [0:0] cby_1__1__46_left_grid_pin_8_;
wire [0:0] cby_1__1__46_left_grid_pin_9_;
wire [0:0] cby_1__1__46_right_grid_pin_52_;
wire [0:0] cby_1__1__47_ccff_tail;
wire [0:19] cby_1__1__47_chany_bottom_out;
wire [0:19] cby_1__1__47_chany_top_out;
wire [0:0] cby_1__1__47_left_grid_pin_0_;
wire [0:0] cby_1__1__47_left_grid_pin_10_;
wire [0:0] cby_1__1__47_left_grid_pin_11_;
wire [0:0] cby_1__1__47_left_grid_pin_12_;
wire [0:0] cby_1__1__47_left_grid_pin_13_;
wire [0:0] cby_1__1__47_left_grid_pin_14_;
wire [0:0] cby_1__1__47_left_grid_pin_15_;
wire [0:0] cby_1__1__47_left_grid_pin_1_;
wire [0:0] cby_1__1__47_left_grid_pin_2_;
wire [0:0] cby_1__1__47_left_grid_pin_3_;
wire [0:0] cby_1__1__47_left_grid_pin_4_;
wire [0:0] cby_1__1__47_left_grid_pin_5_;
wire [0:0] cby_1__1__47_left_grid_pin_6_;
wire [0:0] cby_1__1__47_left_grid_pin_7_;
wire [0:0] cby_1__1__47_left_grid_pin_8_;
wire [0:0] cby_1__1__47_left_grid_pin_9_;
wire [0:0] cby_1__1__47_right_grid_pin_52_;
wire [0:0] cby_1__1__48_ccff_tail;
wire [0:19] cby_1__1__48_chany_bottom_out;
wire [0:19] cby_1__1__48_chany_top_out;
wire [0:0] cby_1__1__48_left_grid_pin_0_;
wire [0:0] cby_1__1__48_left_grid_pin_10_;
wire [0:0] cby_1__1__48_left_grid_pin_11_;
wire [0:0] cby_1__1__48_left_grid_pin_12_;
wire [0:0] cby_1__1__48_left_grid_pin_13_;
wire [0:0] cby_1__1__48_left_grid_pin_14_;
wire [0:0] cby_1__1__48_left_grid_pin_15_;
wire [0:0] cby_1__1__48_left_grid_pin_1_;
wire [0:0] cby_1__1__48_left_grid_pin_2_;
wire [0:0] cby_1__1__48_left_grid_pin_3_;
wire [0:0] cby_1__1__48_left_grid_pin_4_;
wire [0:0] cby_1__1__48_left_grid_pin_5_;
wire [0:0] cby_1__1__48_left_grid_pin_6_;
wire [0:0] cby_1__1__48_left_grid_pin_7_;
wire [0:0] cby_1__1__48_left_grid_pin_8_;
wire [0:0] cby_1__1__48_left_grid_pin_9_;
wire [0:0] cby_1__1__48_right_grid_pin_52_;
wire [0:0] cby_1__1__49_ccff_tail;
wire [0:19] cby_1__1__49_chany_bottom_out;
wire [0:19] cby_1__1__49_chany_top_out;
wire [0:0] cby_1__1__49_left_grid_pin_0_;
wire [0:0] cby_1__1__49_left_grid_pin_10_;
wire [0:0] cby_1__1__49_left_grid_pin_11_;
wire [0:0] cby_1__1__49_left_grid_pin_12_;
wire [0:0] cby_1__1__49_left_grid_pin_13_;
wire [0:0] cby_1__1__49_left_grid_pin_14_;
wire [0:0] cby_1__1__49_left_grid_pin_15_;
wire [0:0] cby_1__1__49_left_grid_pin_1_;
wire [0:0] cby_1__1__49_left_grid_pin_2_;
wire [0:0] cby_1__1__49_left_grid_pin_3_;
wire [0:0] cby_1__1__49_left_grid_pin_4_;
wire [0:0] cby_1__1__49_left_grid_pin_5_;
wire [0:0] cby_1__1__49_left_grid_pin_6_;
wire [0:0] cby_1__1__49_left_grid_pin_7_;
wire [0:0] cby_1__1__49_left_grid_pin_8_;
wire [0:0] cby_1__1__49_left_grid_pin_9_;
wire [0:0] cby_1__1__49_right_grid_pin_52_;
wire [0:0] cby_1__1__4_ccff_tail;
wire [0:19] cby_1__1__4_chany_bottom_out;
wire [0:19] cby_1__1__4_chany_top_out;
wire [0:0] cby_1__1__4_left_grid_pin_0_;
wire [0:0] cby_1__1__4_left_grid_pin_10_;
wire [0:0] cby_1__1__4_left_grid_pin_11_;
wire [0:0] cby_1__1__4_left_grid_pin_12_;
wire [0:0] cby_1__1__4_left_grid_pin_13_;
wire [0:0] cby_1__1__4_left_grid_pin_14_;
wire [0:0] cby_1__1__4_left_grid_pin_15_;
wire [0:0] cby_1__1__4_left_grid_pin_1_;
wire [0:0] cby_1__1__4_left_grid_pin_2_;
wire [0:0] cby_1__1__4_left_grid_pin_3_;
wire [0:0] cby_1__1__4_left_grid_pin_4_;
wire [0:0] cby_1__1__4_left_grid_pin_5_;
wire [0:0] cby_1__1__4_left_grid_pin_6_;
wire [0:0] cby_1__1__4_left_grid_pin_7_;
wire [0:0] cby_1__1__4_left_grid_pin_8_;
wire [0:0] cby_1__1__4_left_grid_pin_9_;
wire [0:0] cby_1__1__4_right_grid_pin_52_;
wire [0:0] cby_1__1__50_ccff_tail;
wire [0:19] cby_1__1__50_chany_bottom_out;
wire [0:19] cby_1__1__50_chany_top_out;
wire [0:0] cby_1__1__50_left_grid_pin_0_;
wire [0:0] cby_1__1__50_left_grid_pin_10_;
wire [0:0] cby_1__1__50_left_grid_pin_11_;
wire [0:0] cby_1__1__50_left_grid_pin_12_;
wire [0:0] cby_1__1__50_left_grid_pin_13_;
wire [0:0] cby_1__1__50_left_grid_pin_14_;
wire [0:0] cby_1__1__50_left_grid_pin_15_;
wire [0:0] cby_1__1__50_left_grid_pin_1_;
wire [0:0] cby_1__1__50_left_grid_pin_2_;
wire [0:0] cby_1__1__50_left_grid_pin_3_;
wire [0:0] cby_1__1__50_left_grid_pin_4_;
wire [0:0] cby_1__1__50_left_grid_pin_5_;
wire [0:0] cby_1__1__50_left_grid_pin_6_;
wire [0:0] cby_1__1__50_left_grid_pin_7_;
wire [0:0] cby_1__1__50_left_grid_pin_8_;
wire [0:0] cby_1__1__50_left_grid_pin_9_;
wire [0:0] cby_1__1__50_right_grid_pin_52_;
wire [0:0] cby_1__1__51_ccff_tail;
wire [0:19] cby_1__1__51_chany_bottom_out;
wire [0:19] cby_1__1__51_chany_top_out;
wire [0:0] cby_1__1__51_left_grid_pin_0_;
wire [0:0] cby_1__1__51_left_grid_pin_10_;
wire [0:0] cby_1__1__51_left_grid_pin_11_;
wire [0:0] cby_1__1__51_left_grid_pin_12_;
wire [0:0] cby_1__1__51_left_grid_pin_13_;
wire [0:0] cby_1__1__51_left_grid_pin_14_;
wire [0:0] cby_1__1__51_left_grid_pin_15_;
wire [0:0] cby_1__1__51_left_grid_pin_1_;
wire [0:0] cby_1__1__51_left_grid_pin_2_;
wire [0:0] cby_1__1__51_left_grid_pin_3_;
wire [0:0] cby_1__1__51_left_grid_pin_4_;
wire [0:0] cby_1__1__51_left_grid_pin_5_;
wire [0:0] cby_1__1__51_left_grid_pin_6_;
wire [0:0] cby_1__1__51_left_grid_pin_7_;
wire [0:0] cby_1__1__51_left_grid_pin_8_;
wire [0:0] cby_1__1__51_left_grid_pin_9_;
wire [0:0] cby_1__1__51_right_grid_pin_52_;
wire [0:0] cby_1__1__52_ccff_tail;
wire [0:19] cby_1__1__52_chany_bottom_out;
wire [0:19] cby_1__1__52_chany_top_out;
wire [0:0] cby_1__1__52_left_grid_pin_0_;
wire [0:0] cby_1__1__52_left_grid_pin_10_;
wire [0:0] cby_1__1__52_left_grid_pin_11_;
wire [0:0] cby_1__1__52_left_grid_pin_12_;
wire [0:0] cby_1__1__52_left_grid_pin_13_;
wire [0:0] cby_1__1__52_left_grid_pin_14_;
wire [0:0] cby_1__1__52_left_grid_pin_15_;
wire [0:0] cby_1__1__52_left_grid_pin_1_;
wire [0:0] cby_1__1__52_left_grid_pin_2_;
wire [0:0] cby_1__1__52_left_grid_pin_3_;
wire [0:0] cby_1__1__52_left_grid_pin_4_;
wire [0:0] cby_1__1__52_left_grid_pin_5_;
wire [0:0] cby_1__1__52_left_grid_pin_6_;
wire [0:0] cby_1__1__52_left_grid_pin_7_;
wire [0:0] cby_1__1__52_left_grid_pin_8_;
wire [0:0] cby_1__1__52_left_grid_pin_9_;
wire [0:0] cby_1__1__52_right_grid_pin_52_;
wire [0:0] cby_1__1__53_ccff_tail;
wire [0:19] cby_1__1__53_chany_bottom_out;
wire [0:19] cby_1__1__53_chany_top_out;
wire [0:0] cby_1__1__53_left_grid_pin_0_;
wire [0:0] cby_1__1__53_left_grid_pin_10_;
wire [0:0] cby_1__1__53_left_grid_pin_11_;
wire [0:0] cby_1__1__53_left_grid_pin_12_;
wire [0:0] cby_1__1__53_left_grid_pin_13_;
wire [0:0] cby_1__1__53_left_grid_pin_14_;
wire [0:0] cby_1__1__53_left_grid_pin_15_;
wire [0:0] cby_1__1__53_left_grid_pin_1_;
wire [0:0] cby_1__1__53_left_grid_pin_2_;
wire [0:0] cby_1__1__53_left_grid_pin_3_;
wire [0:0] cby_1__1__53_left_grid_pin_4_;
wire [0:0] cby_1__1__53_left_grid_pin_5_;
wire [0:0] cby_1__1__53_left_grid_pin_6_;
wire [0:0] cby_1__1__53_left_grid_pin_7_;
wire [0:0] cby_1__1__53_left_grid_pin_8_;
wire [0:0] cby_1__1__53_left_grid_pin_9_;
wire [0:0] cby_1__1__53_right_grid_pin_52_;
wire [0:0] cby_1__1__54_ccff_tail;
wire [0:19] cby_1__1__54_chany_bottom_out;
wire [0:19] cby_1__1__54_chany_top_out;
wire [0:0] cby_1__1__54_left_grid_pin_0_;
wire [0:0] cby_1__1__54_left_grid_pin_10_;
wire [0:0] cby_1__1__54_left_grid_pin_11_;
wire [0:0] cby_1__1__54_left_grid_pin_12_;
wire [0:0] cby_1__1__54_left_grid_pin_13_;
wire [0:0] cby_1__1__54_left_grid_pin_14_;
wire [0:0] cby_1__1__54_left_grid_pin_15_;
wire [0:0] cby_1__1__54_left_grid_pin_1_;
wire [0:0] cby_1__1__54_left_grid_pin_2_;
wire [0:0] cby_1__1__54_left_grid_pin_3_;
wire [0:0] cby_1__1__54_left_grid_pin_4_;
wire [0:0] cby_1__1__54_left_grid_pin_5_;
wire [0:0] cby_1__1__54_left_grid_pin_6_;
wire [0:0] cby_1__1__54_left_grid_pin_7_;
wire [0:0] cby_1__1__54_left_grid_pin_8_;
wire [0:0] cby_1__1__54_left_grid_pin_9_;
wire [0:0] cby_1__1__54_right_grid_pin_52_;
wire [0:0] cby_1__1__55_ccff_tail;
wire [0:19] cby_1__1__55_chany_bottom_out;
wire [0:19] cby_1__1__55_chany_top_out;
wire [0:0] cby_1__1__55_left_grid_pin_0_;
wire [0:0] cby_1__1__55_left_grid_pin_10_;
wire [0:0] cby_1__1__55_left_grid_pin_11_;
wire [0:0] cby_1__1__55_left_grid_pin_12_;
wire [0:0] cby_1__1__55_left_grid_pin_13_;
wire [0:0] cby_1__1__55_left_grid_pin_14_;
wire [0:0] cby_1__1__55_left_grid_pin_15_;
wire [0:0] cby_1__1__55_left_grid_pin_1_;
wire [0:0] cby_1__1__55_left_grid_pin_2_;
wire [0:0] cby_1__1__55_left_grid_pin_3_;
wire [0:0] cby_1__1__55_left_grid_pin_4_;
wire [0:0] cby_1__1__55_left_grid_pin_5_;
wire [0:0] cby_1__1__55_left_grid_pin_6_;
wire [0:0] cby_1__1__55_left_grid_pin_7_;
wire [0:0] cby_1__1__55_left_grid_pin_8_;
wire [0:0] cby_1__1__55_left_grid_pin_9_;
wire [0:0] cby_1__1__55_right_grid_pin_52_;
wire [0:0] cby_1__1__56_ccff_tail;
wire [0:19] cby_1__1__56_chany_bottom_out;
wire [0:19] cby_1__1__56_chany_top_out;
wire [0:0] cby_1__1__56_left_grid_pin_0_;
wire [0:0] cby_1__1__56_left_grid_pin_10_;
wire [0:0] cby_1__1__56_left_grid_pin_11_;
wire [0:0] cby_1__1__56_left_grid_pin_12_;
wire [0:0] cby_1__1__56_left_grid_pin_13_;
wire [0:0] cby_1__1__56_left_grid_pin_14_;
wire [0:0] cby_1__1__56_left_grid_pin_15_;
wire [0:0] cby_1__1__56_left_grid_pin_1_;
wire [0:0] cby_1__1__56_left_grid_pin_2_;
wire [0:0] cby_1__1__56_left_grid_pin_3_;
wire [0:0] cby_1__1__56_left_grid_pin_4_;
wire [0:0] cby_1__1__56_left_grid_pin_5_;
wire [0:0] cby_1__1__56_left_grid_pin_6_;
wire [0:0] cby_1__1__56_left_grid_pin_7_;
wire [0:0] cby_1__1__56_left_grid_pin_8_;
wire [0:0] cby_1__1__56_left_grid_pin_9_;
wire [0:0] cby_1__1__56_right_grid_pin_52_;
wire [0:0] cby_1__1__57_ccff_tail;
wire [0:19] cby_1__1__57_chany_bottom_out;
wire [0:19] cby_1__1__57_chany_top_out;
wire [0:0] cby_1__1__57_left_grid_pin_0_;
wire [0:0] cby_1__1__57_left_grid_pin_10_;
wire [0:0] cby_1__1__57_left_grid_pin_11_;
wire [0:0] cby_1__1__57_left_grid_pin_12_;
wire [0:0] cby_1__1__57_left_grid_pin_13_;
wire [0:0] cby_1__1__57_left_grid_pin_14_;
wire [0:0] cby_1__1__57_left_grid_pin_15_;
wire [0:0] cby_1__1__57_left_grid_pin_1_;
wire [0:0] cby_1__1__57_left_grid_pin_2_;
wire [0:0] cby_1__1__57_left_grid_pin_3_;
wire [0:0] cby_1__1__57_left_grid_pin_4_;
wire [0:0] cby_1__1__57_left_grid_pin_5_;
wire [0:0] cby_1__1__57_left_grid_pin_6_;
wire [0:0] cby_1__1__57_left_grid_pin_7_;
wire [0:0] cby_1__1__57_left_grid_pin_8_;
wire [0:0] cby_1__1__57_left_grid_pin_9_;
wire [0:0] cby_1__1__57_right_grid_pin_52_;
wire [0:0] cby_1__1__58_ccff_tail;
wire [0:19] cby_1__1__58_chany_bottom_out;
wire [0:19] cby_1__1__58_chany_top_out;
wire [0:0] cby_1__1__58_left_grid_pin_0_;
wire [0:0] cby_1__1__58_left_grid_pin_10_;
wire [0:0] cby_1__1__58_left_grid_pin_11_;
wire [0:0] cby_1__1__58_left_grid_pin_12_;
wire [0:0] cby_1__1__58_left_grid_pin_13_;
wire [0:0] cby_1__1__58_left_grid_pin_14_;
wire [0:0] cby_1__1__58_left_grid_pin_15_;
wire [0:0] cby_1__1__58_left_grid_pin_1_;
wire [0:0] cby_1__1__58_left_grid_pin_2_;
wire [0:0] cby_1__1__58_left_grid_pin_3_;
wire [0:0] cby_1__1__58_left_grid_pin_4_;
wire [0:0] cby_1__1__58_left_grid_pin_5_;
wire [0:0] cby_1__1__58_left_grid_pin_6_;
wire [0:0] cby_1__1__58_left_grid_pin_7_;
wire [0:0] cby_1__1__58_left_grid_pin_8_;
wire [0:0] cby_1__1__58_left_grid_pin_9_;
wire [0:0] cby_1__1__58_right_grid_pin_52_;
wire [0:0] cby_1__1__59_ccff_tail;
wire [0:19] cby_1__1__59_chany_bottom_out;
wire [0:19] cby_1__1__59_chany_top_out;
wire [0:0] cby_1__1__59_left_grid_pin_0_;
wire [0:0] cby_1__1__59_left_grid_pin_10_;
wire [0:0] cby_1__1__59_left_grid_pin_11_;
wire [0:0] cby_1__1__59_left_grid_pin_12_;
wire [0:0] cby_1__1__59_left_grid_pin_13_;
wire [0:0] cby_1__1__59_left_grid_pin_14_;
wire [0:0] cby_1__1__59_left_grid_pin_15_;
wire [0:0] cby_1__1__59_left_grid_pin_1_;
wire [0:0] cby_1__1__59_left_grid_pin_2_;
wire [0:0] cby_1__1__59_left_grid_pin_3_;
wire [0:0] cby_1__1__59_left_grid_pin_4_;
wire [0:0] cby_1__1__59_left_grid_pin_5_;
wire [0:0] cby_1__1__59_left_grid_pin_6_;
wire [0:0] cby_1__1__59_left_grid_pin_7_;
wire [0:0] cby_1__1__59_left_grid_pin_8_;
wire [0:0] cby_1__1__59_left_grid_pin_9_;
wire [0:0] cby_1__1__59_right_grid_pin_52_;
wire [0:0] cby_1__1__5_ccff_tail;
wire [0:19] cby_1__1__5_chany_bottom_out;
wire [0:19] cby_1__1__5_chany_top_out;
wire [0:0] cby_1__1__5_left_grid_pin_0_;
wire [0:0] cby_1__1__5_left_grid_pin_10_;
wire [0:0] cby_1__1__5_left_grid_pin_11_;
wire [0:0] cby_1__1__5_left_grid_pin_12_;
wire [0:0] cby_1__1__5_left_grid_pin_13_;
wire [0:0] cby_1__1__5_left_grid_pin_14_;
wire [0:0] cby_1__1__5_left_grid_pin_15_;
wire [0:0] cby_1__1__5_left_grid_pin_1_;
wire [0:0] cby_1__1__5_left_grid_pin_2_;
wire [0:0] cby_1__1__5_left_grid_pin_3_;
wire [0:0] cby_1__1__5_left_grid_pin_4_;
wire [0:0] cby_1__1__5_left_grid_pin_5_;
wire [0:0] cby_1__1__5_left_grid_pin_6_;
wire [0:0] cby_1__1__5_left_grid_pin_7_;
wire [0:0] cby_1__1__5_left_grid_pin_8_;
wire [0:0] cby_1__1__5_left_grid_pin_9_;
wire [0:0] cby_1__1__5_right_grid_pin_52_;
wire [0:0] cby_1__1__60_ccff_tail;
wire [0:19] cby_1__1__60_chany_bottom_out;
wire [0:19] cby_1__1__60_chany_top_out;
wire [0:0] cby_1__1__60_left_grid_pin_0_;
wire [0:0] cby_1__1__60_left_grid_pin_10_;
wire [0:0] cby_1__1__60_left_grid_pin_11_;
wire [0:0] cby_1__1__60_left_grid_pin_12_;
wire [0:0] cby_1__1__60_left_grid_pin_13_;
wire [0:0] cby_1__1__60_left_grid_pin_14_;
wire [0:0] cby_1__1__60_left_grid_pin_15_;
wire [0:0] cby_1__1__60_left_grid_pin_1_;
wire [0:0] cby_1__1__60_left_grid_pin_2_;
wire [0:0] cby_1__1__60_left_grid_pin_3_;
wire [0:0] cby_1__1__60_left_grid_pin_4_;
wire [0:0] cby_1__1__60_left_grid_pin_5_;
wire [0:0] cby_1__1__60_left_grid_pin_6_;
wire [0:0] cby_1__1__60_left_grid_pin_7_;
wire [0:0] cby_1__1__60_left_grid_pin_8_;
wire [0:0] cby_1__1__60_left_grid_pin_9_;
wire [0:0] cby_1__1__60_right_grid_pin_52_;
wire [0:0] cby_1__1__61_ccff_tail;
wire [0:19] cby_1__1__61_chany_bottom_out;
wire [0:19] cby_1__1__61_chany_top_out;
wire [0:0] cby_1__1__61_left_grid_pin_0_;
wire [0:0] cby_1__1__61_left_grid_pin_10_;
wire [0:0] cby_1__1__61_left_grid_pin_11_;
wire [0:0] cby_1__1__61_left_grid_pin_12_;
wire [0:0] cby_1__1__61_left_grid_pin_13_;
wire [0:0] cby_1__1__61_left_grid_pin_14_;
wire [0:0] cby_1__1__61_left_grid_pin_15_;
wire [0:0] cby_1__1__61_left_grid_pin_1_;
wire [0:0] cby_1__1__61_left_grid_pin_2_;
wire [0:0] cby_1__1__61_left_grid_pin_3_;
wire [0:0] cby_1__1__61_left_grid_pin_4_;
wire [0:0] cby_1__1__61_left_grid_pin_5_;
wire [0:0] cby_1__1__61_left_grid_pin_6_;
wire [0:0] cby_1__1__61_left_grid_pin_7_;
wire [0:0] cby_1__1__61_left_grid_pin_8_;
wire [0:0] cby_1__1__61_left_grid_pin_9_;
wire [0:0] cby_1__1__61_right_grid_pin_52_;
wire [0:0] cby_1__1__62_ccff_tail;
wire [0:19] cby_1__1__62_chany_bottom_out;
wire [0:19] cby_1__1__62_chany_top_out;
wire [0:0] cby_1__1__62_left_grid_pin_0_;
wire [0:0] cby_1__1__62_left_grid_pin_10_;
wire [0:0] cby_1__1__62_left_grid_pin_11_;
wire [0:0] cby_1__1__62_left_grid_pin_12_;
wire [0:0] cby_1__1__62_left_grid_pin_13_;
wire [0:0] cby_1__1__62_left_grid_pin_14_;
wire [0:0] cby_1__1__62_left_grid_pin_15_;
wire [0:0] cby_1__1__62_left_grid_pin_1_;
wire [0:0] cby_1__1__62_left_grid_pin_2_;
wire [0:0] cby_1__1__62_left_grid_pin_3_;
wire [0:0] cby_1__1__62_left_grid_pin_4_;
wire [0:0] cby_1__1__62_left_grid_pin_5_;
wire [0:0] cby_1__1__62_left_grid_pin_6_;
wire [0:0] cby_1__1__62_left_grid_pin_7_;
wire [0:0] cby_1__1__62_left_grid_pin_8_;
wire [0:0] cby_1__1__62_left_grid_pin_9_;
wire [0:0] cby_1__1__62_right_grid_pin_52_;
wire [0:0] cby_1__1__63_ccff_tail;
wire [0:19] cby_1__1__63_chany_bottom_out;
wire [0:19] cby_1__1__63_chany_top_out;
wire [0:0] cby_1__1__63_left_grid_pin_0_;
wire [0:0] cby_1__1__63_left_grid_pin_10_;
wire [0:0] cby_1__1__63_left_grid_pin_11_;
wire [0:0] cby_1__1__63_left_grid_pin_12_;
wire [0:0] cby_1__1__63_left_grid_pin_13_;
wire [0:0] cby_1__1__63_left_grid_pin_14_;
wire [0:0] cby_1__1__63_left_grid_pin_15_;
wire [0:0] cby_1__1__63_left_grid_pin_1_;
wire [0:0] cby_1__1__63_left_grid_pin_2_;
wire [0:0] cby_1__1__63_left_grid_pin_3_;
wire [0:0] cby_1__1__63_left_grid_pin_4_;
wire [0:0] cby_1__1__63_left_grid_pin_5_;
wire [0:0] cby_1__1__63_left_grid_pin_6_;
wire [0:0] cby_1__1__63_left_grid_pin_7_;
wire [0:0] cby_1__1__63_left_grid_pin_8_;
wire [0:0] cby_1__1__63_left_grid_pin_9_;
wire [0:0] cby_1__1__63_right_grid_pin_52_;
wire [0:0] cby_1__1__64_ccff_tail;
wire [0:19] cby_1__1__64_chany_bottom_out;
wire [0:19] cby_1__1__64_chany_top_out;
wire [0:0] cby_1__1__64_left_grid_pin_0_;
wire [0:0] cby_1__1__64_left_grid_pin_10_;
wire [0:0] cby_1__1__64_left_grid_pin_11_;
wire [0:0] cby_1__1__64_left_grid_pin_12_;
wire [0:0] cby_1__1__64_left_grid_pin_13_;
wire [0:0] cby_1__1__64_left_grid_pin_14_;
wire [0:0] cby_1__1__64_left_grid_pin_15_;
wire [0:0] cby_1__1__64_left_grid_pin_1_;
wire [0:0] cby_1__1__64_left_grid_pin_2_;
wire [0:0] cby_1__1__64_left_grid_pin_3_;
wire [0:0] cby_1__1__64_left_grid_pin_4_;
wire [0:0] cby_1__1__64_left_grid_pin_5_;
wire [0:0] cby_1__1__64_left_grid_pin_6_;
wire [0:0] cby_1__1__64_left_grid_pin_7_;
wire [0:0] cby_1__1__64_left_grid_pin_8_;
wire [0:0] cby_1__1__64_left_grid_pin_9_;
wire [0:0] cby_1__1__64_right_grid_pin_52_;
wire [0:0] cby_1__1__65_ccff_tail;
wire [0:19] cby_1__1__65_chany_bottom_out;
wire [0:19] cby_1__1__65_chany_top_out;
wire [0:0] cby_1__1__65_left_grid_pin_0_;
wire [0:0] cby_1__1__65_left_grid_pin_10_;
wire [0:0] cby_1__1__65_left_grid_pin_11_;
wire [0:0] cby_1__1__65_left_grid_pin_12_;
wire [0:0] cby_1__1__65_left_grid_pin_13_;
wire [0:0] cby_1__1__65_left_grid_pin_14_;
wire [0:0] cby_1__1__65_left_grid_pin_15_;
wire [0:0] cby_1__1__65_left_grid_pin_1_;
wire [0:0] cby_1__1__65_left_grid_pin_2_;
wire [0:0] cby_1__1__65_left_grid_pin_3_;
wire [0:0] cby_1__1__65_left_grid_pin_4_;
wire [0:0] cby_1__1__65_left_grid_pin_5_;
wire [0:0] cby_1__1__65_left_grid_pin_6_;
wire [0:0] cby_1__1__65_left_grid_pin_7_;
wire [0:0] cby_1__1__65_left_grid_pin_8_;
wire [0:0] cby_1__1__65_left_grid_pin_9_;
wire [0:0] cby_1__1__65_right_grid_pin_52_;
wire [0:0] cby_1__1__66_ccff_tail;
wire [0:19] cby_1__1__66_chany_bottom_out;
wire [0:19] cby_1__1__66_chany_top_out;
wire [0:0] cby_1__1__66_left_grid_pin_0_;
wire [0:0] cby_1__1__66_left_grid_pin_10_;
wire [0:0] cby_1__1__66_left_grid_pin_11_;
wire [0:0] cby_1__1__66_left_grid_pin_12_;
wire [0:0] cby_1__1__66_left_grid_pin_13_;
wire [0:0] cby_1__1__66_left_grid_pin_14_;
wire [0:0] cby_1__1__66_left_grid_pin_15_;
wire [0:0] cby_1__1__66_left_grid_pin_1_;
wire [0:0] cby_1__1__66_left_grid_pin_2_;
wire [0:0] cby_1__1__66_left_grid_pin_3_;
wire [0:0] cby_1__1__66_left_grid_pin_4_;
wire [0:0] cby_1__1__66_left_grid_pin_5_;
wire [0:0] cby_1__1__66_left_grid_pin_6_;
wire [0:0] cby_1__1__66_left_grid_pin_7_;
wire [0:0] cby_1__1__66_left_grid_pin_8_;
wire [0:0] cby_1__1__66_left_grid_pin_9_;
wire [0:0] cby_1__1__66_right_grid_pin_52_;
wire [0:0] cby_1__1__67_ccff_tail;
wire [0:19] cby_1__1__67_chany_bottom_out;
wire [0:19] cby_1__1__67_chany_top_out;
wire [0:0] cby_1__1__67_left_grid_pin_0_;
wire [0:0] cby_1__1__67_left_grid_pin_10_;
wire [0:0] cby_1__1__67_left_grid_pin_11_;
wire [0:0] cby_1__1__67_left_grid_pin_12_;
wire [0:0] cby_1__1__67_left_grid_pin_13_;
wire [0:0] cby_1__1__67_left_grid_pin_14_;
wire [0:0] cby_1__1__67_left_grid_pin_15_;
wire [0:0] cby_1__1__67_left_grid_pin_1_;
wire [0:0] cby_1__1__67_left_grid_pin_2_;
wire [0:0] cby_1__1__67_left_grid_pin_3_;
wire [0:0] cby_1__1__67_left_grid_pin_4_;
wire [0:0] cby_1__1__67_left_grid_pin_5_;
wire [0:0] cby_1__1__67_left_grid_pin_6_;
wire [0:0] cby_1__1__67_left_grid_pin_7_;
wire [0:0] cby_1__1__67_left_grid_pin_8_;
wire [0:0] cby_1__1__67_left_grid_pin_9_;
wire [0:0] cby_1__1__67_right_grid_pin_52_;
wire [0:0] cby_1__1__68_ccff_tail;
wire [0:19] cby_1__1__68_chany_bottom_out;
wire [0:19] cby_1__1__68_chany_top_out;
wire [0:0] cby_1__1__68_left_grid_pin_0_;
wire [0:0] cby_1__1__68_left_grid_pin_10_;
wire [0:0] cby_1__1__68_left_grid_pin_11_;
wire [0:0] cby_1__1__68_left_grid_pin_12_;
wire [0:0] cby_1__1__68_left_grid_pin_13_;
wire [0:0] cby_1__1__68_left_grid_pin_14_;
wire [0:0] cby_1__1__68_left_grid_pin_15_;
wire [0:0] cby_1__1__68_left_grid_pin_1_;
wire [0:0] cby_1__1__68_left_grid_pin_2_;
wire [0:0] cby_1__1__68_left_grid_pin_3_;
wire [0:0] cby_1__1__68_left_grid_pin_4_;
wire [0:0] cby_1__1__68_left_grid_pin_5_;
wire [0:0] cby_1__1__68_left_grid_pin_6_;
wire [0:0] cby_1__1__68_left_grid_pin_7_;
wire [0:0] cby_1__1__68_left_grid_pin_8_;
wire [0:0] cby_1__1__68_left_grid_pin_9_;
wire [0:0] cby_1__1__68_right_grid_pin_52_;
wire [0:0] cby_1__1__69_ccff_tail;
wire [0:19] cby_1__1__69_chany_bottom_out;
wire [0:19] cby_1__1__69_chany_top_out;
wire [0:0] cby_1__1__69_left_grid_pin_0_;
wire [0:0] cby_1__1__69_left_grid_pin_10_;
wire [0:0] cby_1__1__69_left_grid_pin_11_;
wire [0:0] cby_1__1__69_left_grid_pin_12_;
wire [0:0] cby_1__1__69_left_grid_pin_13_;
wire [0:0] cby_1__1__69_left_grid_pin_14_;
wire [0:0] cby_1__1__69_left_grid_pin_15_;
wire [0:0] cby_1__1__69_left_grid_pin_1_;
wire [0:0] cby_1__1__69_left_grid_pin_2_;
wire [0:0] cby_1__1__69_left_grid_pin_3_;
wire [0:0] cby_1__1__69_left_grid_pin_4_;
wire [0:0] cby_1__1__69_left_grid_pin_5_;
wire [0:0] cby_1__1__69_left_grid_pin_6_;
wire [0:0] cby_1__1__69_left_grid_pin_7_;
wire [0:0] cby_1__1__69_left_grid_pin_8_;
wire [0:0] cby_1__1__69_left_grid_pin_9_;
wire [0:0] cby_1__1__69_right_grid_pin_52_;
wire [0:0] cby_1__1__6_ccff_tail;
wire [0:19] cby_1__1__6_chany_bottom_out;
wire [0:19] cby_1__1__6_chany_top_out;
wire [0:0] cby_1__1__6_left_grid_pin_0_;
wire [0:0] cby_1__1__6_left_grid_pin_10_;
wire [0:0] cby_1__1__6_left_grid_pin_11_;
wire [0:0] cby_1__1__6_left_grid_pin_12_;
wire [0:0] cby_1__1__6_left_grid_pin_13_;
wire [0:0] cby_1__1__6_left_grid_pin_14_;
wire [0:0] cby_1__1__6_left_grid_pin_15_;
wire [0:0] cby_1__1__6_left_grid_pin_1_;
wire [0:0] cby_1__1__6_left_grid_pin_2_;
wire [0:0] cby_1__1__6_left_grid_pin_3_;
wire [0:0] cby_1__1__6_left_grid_pin_4_;
wire [0:0] cby_1__1__6_left_grid_pin_5_;
wire [0:0] cby_1__1__6_left_grid_pin_6_;
wire [0:0] cby_1__1__6_left_grid_pin_7_;
wire [0:0] cby_1__1__6_left_grid_pin_8_;
wire [0:0] cby_1__1__6_left_grid_pin_9_;
wire [0:0] cby_1__1__6_right_grid_pin_52_;
wire [0:0] cby_1__1__70_ccff_tail;
wire [0:19] cby_1__1__70_chany_bottom_out;
wire [0:19] cby_1__1__70_chany_top_out;
wire [0:0] cby_1__1__70_left_grid_pin_0_;
wire [0:0] cby_1__1__70_left_grid_pin_10_;
wire [0:0] cby_1__1__70_left_grid_pin_11_;
wire [0:0] cby_1__1__70_left_grid_pin_12_;
wire [0:0] cby_1__1__70_left_grid_pin_13_;
wire [0:0] cby_1__1__70_left_grid_pin_14_;
wire [0:0] cby_1__1__70_left_grid_pin_15_;
wire [0:0] cby_1__1__70_left_grid_pin_1_;
wire [0:0] cby_1__1__70_left_grid_pin_2_;
wire [0:0] cby_1__1__70_left_grid_pin_3_;
wire [0:0] cby_1__1__70_left_grid_pin_4_;
wire [0:0] cby_1__1__70_left_grid_pin_5_;
wire [0:0] cby_1__1__70_left_grid_pin_6_;
wire [0:0] cby_1__1__70_left_grid_pin_7_;
wire [0:0] cby_1__1__70_left_grid_pin_8_;
wire [0:0] cby_1__1__70_left_grid_pin_9_;
wire [0:0] cby_1__1__70_right_grid_pin_52_;
wire [0:0] cby_1__1__71_ccff_tail;
wire [0:19] cby_1__1__71_chany_bottom_out;
wire [0:19] cby_1__1__71_chany_top_out;
wire [0:0] cby_1__1__71_left_grid_pin_0_;
wire [0:0] cby_1__1__71_left_grid_pin_10_;
wire [0:0] cby_1__1__71_left_grid_pin_11_;
wire [0:0] cby_1__1__71_left_grid_pin_12_;
wire [0:0] cby_1__1__71_left_grid_pin_13_;
wire [0:0] cby_1__1__71_left_grid_pin_14_;
wire [0:0] cby_1__1__71_left_grid_pin_15_;
wire [0:0] cby_1__1__71_left_grid_pin_1_;
wire [0:0] cby_1__1__71_left_grid_pin_2_;
wire [0:0] cby_1__1__71_left_grid_pin_3_;
wire [0:0] cby_1__1__71_left_grid_pin_4_;
wire [0:0] cby_1__1__71_left_grid_pin_5_;
wire [0:0] cby_1__1__71_left_grid_pin_6_;
wire [0:0] cby_1__1__71_left_grid_pin_7_;
wire [0:0] cby_1__1__71_left_grid_pin_8_;
wire [0:0] cby_1__1__71_left_grid_pin_9_;
wire [0:0] cby_1__1__71_right_grid_pin_52_;
wire [0:0] cby_1__1__72_ccff_tail;
wire [0:19] cby_1__1__72_chany_bottom_out;
wire [0:19] cby_1__1__72_chany_top_out;
wire [0:0] cby_1__1__72_left_grid_pin_0_;
wire [0:0] cby_1__1__72_left_grid_pin_10_;
wire [0:0] cby_1__1__72_left_grid_pin_11_;
wire [0:0] cby_1__1__72_left_grid_pin_12_;
wire [0:0] cby_1__1__72_left_grid_pin_13_;
wire [0:0] cby_1__1__72_left_grid_pin_14_;
wire [0:0] cby_1__1__72_left_grid_pin_15_;
wire [0:0] cby_1__1__72_left_grid_pin_1_;
wire [0:0] cby_1__1__72_left_grid_pin_2_;
wire [0:0] cby_1__1__72_left_grid_pin_3_;
wire [0:0] cby_1__1__72_left_grid_pin_4_;
wire [0:0] cby_1__1__72_left_grid_pin_5_;
wire [0:0] cby_1__1__72_left_grid_pin_6_;
wire [0:0] cby_1__1__72_left_grid_pin_7_;
wire [0:0] cby_1__1__72_left_grid_pin_8_;
wire [0:0] cby_1__1__72_left_grid_pin_9_;
wire [0:0] cby_1__1__72_right_grid_pin_52_;
wire [0:0] cby_1__1__73_ccff_tail;
wire [0:19] cby_1__1__73_chany_bottom_out;
wire [0:19] cby_1__1__73_chany_top_out;
wire [0:0] cby_1__1__73_left_grid_pin_0_;
wire [0:0] cby_1__1__73_left_grid_pin_10_;
wire [0:0] cby_1__1__73_left_grid_pin_11_;
wire [0:0] cby_1__1__73_left_grid_pin_12_;
wire [0:0] cby_1__1__73_left_grid_pin_13_;
wire [0:0] cby_1__1__73_left_grid_pin_14_;
wire [0:0] cby_1__1__73_left_grid_pin_15_;
wire [0:0] cby_1__1__73_left_grid_pin_1_;
wire [0:0] cby_1__1__73_left_grid_pin_2_;
wire [0:0] cby_1__1__73_left_grid_pin_3_;
wire [0:0] cby_1__1__73_left_grid_pin_4_;
wire [0:0] cby_1__1__73_left_grid_pin_5_;
wire [0:0] cby_1__1__73_left_grid_pin_6_;
wire [0:0] cby_1__1__73_left_grid_pin_7_;
wire [0:0] cby_1__1__73_left_grid_pin_8_;
wire [0:0] cby_1__1__73_left_grid_pin_9_;
wire [0:0] cby_1__1__73_right_grid_pin_52_;
wire [0:0] cby_1__1__74_ccff_tail;
wire [0:19] cby_1__1__74_chany_bottom_out;
wire [0:19] cby_1__1__74_chany_top_out;
wire [0:0] cby_1__1__74_left_grid_pin_0_;
wire [0:0] cby_1__1__74_left_grid_pin_10_;
wire [0:0] cby_1__1__74_left_grid_pin_11_;
wire [0:0] cby_1__1__74_left_grid_pin_12_;
wire [0:0] cby_1__1__74_left_grid_pin_13_;
wire [0:0] cby_1__1__74_left_grid_pin_14_;
wire [0:0] cby_1__1__74_left_grid_pin_15_;
wire [0:0] cby_1__1__74_left_grid_pin_1_;
wire [0:0] cby_1__1__74_left_grid_pin_2_;
wire [0:0] cby_1__1__74_left_grid_pin_3_;
wire [0:0] cby_1__1__74_left_grid_pin_4_;
wire [0:0] cby_1__1__74_left_grid_pin_5_;
wire [0:0] cby_1__1__74_left_grid_pin_6_;
wire [0:0] cby_1__1__74_left_grid_pin_7_;
wire [0:0] cby_1__1__74_left_grid_pin_8_;
wire [0:0] cby_1__1__74_left_grid_pin_9_;
wire [0:0] cby_1__1__74_right_grid_pin_52_;
wire [0:0] cby_1__1__75_ccff_tail;
wire [0:19] cby_1__1__75_chany_bottom_out;
wire [0:19] cby_1__1__75_chany_top_out;
wire [0:0] cby_1__1__75_left_grid_pin_0_;
wire [0:0] cby_1__1__75_left_grid_pin_10_;
wire [0:0] cby_1__1__75_left_grid_pin_11_;
wire [0:0] cby_1__1__75_left_grid_pin_12_;
wire [0:0] cby_1__1__75_left_grid_pin_13_;
wire [0:0] cby_1__1__75_left_grid_pin_14_;
wire [0:0] cby_1__1__75_left_grid_pin_15_;
wire [0:0] cby_1__1__75_left_grid_pin_1_;
wire [0:0] cby_1__1__75_left_grid_pin_2_;
wire [0:0] cby_1__1__75_left_grid_pin_3_;
wire [0:0] cby_1__1__75_left_grid_pin_4_;
wire [0:0] cby_1__1__75_left_grid_pin_5_;
wire [0:0] cby_1__1__75_left_grid_pin_6_;
wire [0:0] cby_1__1__75_left_grid_pin_7_;
wire [0:0] cby_1__1__75_left_grid_pin_8_;
wire [0:0] cby_1__1__75_left_grid_pin_9_;
wire [0:0] cby_1__1__75_right_grid_pin_52_;
wire [0:0] cby_1__1__76_ccff_tail;
wire [0:19] cby_1__1__76_chany_bottom_out;
wire [0:19] cby_1__1__76_chany_top_out;
wire [0:0] cby_1__1__76_left_grid_pin_0_;
wire [0:0] cby_1__1__76_left_grid_pin_10_;
wire [0:0] cby_1__1__76_left_grid_pin_11_;
wire [0:0] cby_1__1__76_left_grid_pin_12_;
wire [0:0] cby_1__1__76_left_grid_pin_13_;
wire [0:0] cby_1__1__76_left_grid_pin_14_;
wire [0:0] cby_1__1__76_left_grid_pin_15_;
wire [0:0] cby_1__1__76_left_grid_pin_1_;
wire [0:0] cby_1__1__76_left_grid_pin_2_;
wire [0:0] cby_1__1__76_left_grid_pin_3_;
wire [0:0] cby_1__1__76_left_grid_pin_4_;
wire [0:0] cby_1__1__76_left_grid_pin_5_;
wire [0:0] cby_1__1__76_left_grid_pin_6_;
wire [0:0] cby_1__1__76_left_grid_pin_7_;
wire [0:0] cby_1__1__76_left_grid_pin_8_;
wire [0:0] cby_1__1__76_left_grid_pin_9_;
wire [0:0] cby_1__1__76_right_grid_pin_52_;
wire [0:0] cby_1__1__77_ccff_tail;
wire [0:19] cby_1__1__77_chany_bottom_out;
wire [0:19] cby_1__1__77_chany_top_out;
wire [0:0] cby_1__1__77_left_grid_pin_0_;
wire [0:0] cby_1__1__77_left_grid_pin_10_;
wire [0:0] cby_1__1__77_left_grid_pin_11_;
wire [0:0] cby_1__1__77_left_grid_pin_12_;
wire [0:0] cby_1__1__77_left_grid_pin_13_;
wire [0:0] cby_1__1__77_left_grid_pin_14_;
wire [0:0] cby_1__1__77_left_grid_pin_15_;
wire [0:0] cby_1__1__77_left_grid_pin_1_;
wire [0:0] cby_1__1__77_left_grid_pin_2_;
wire [0:0] cby_1__1__77_left_grid_pin_3_;
wire [0:0] cby_1__1__77_left_grid_pin_4_;
wire [0:0] cby_1__1__77_left_grid_pin_5_;
wire [0:0] cby_1__1__77_left_grid_pin_6_;
wire [0:0] cby_1__1__77_left_grid_pin_7_;
wire [0:0] cby_1__1__77_left_grid_pin_8_;
wire [0:0] cby_1__1__77_left_grid_pin_9_;
wire [0:0] cby_1__1__77_right_grid_pin_52_;
wire [0:0] cby_1__1__78_ccff_tail;
wire [0:19] cby_1__1__78_chany_bottom_out;
wire [0:19] cby_1__1__78_chany_top_out;
wire [0:0] cby_1__1__78_left_grid_pin_0_;
wire [0:0] cby_1__1__78_left_grid_pin_10_;
wire [0:0] cby_1__1__78_left_grid_pin_11_;
wire [0:0] cby_1__1__78_left_grid_pin_12_;
wire [0:0] cby_1__1__78_left_grid_pin_13_;
wire [0:0] cby_1__1__78_left_grid_pin_14_;
wire [0:0] cby_1__1__78_left_grid_pin_15_;
wire [0:0] cby_1__1__78_left_grid_pin_1_;
wire [0:0] cby_1__1__78_left_grid_pin_2_;
wire [0:0] cby_1__1__78_left_grid_pin_3_;
wire [0:0] cby_1__1__78_left_grid_pin_4_;
wire [0:0] cby_1__1__78_left_grid_pin_5_;
wire [0:0] cby_1__1__78_left_grid_pin_6_;
wire [0:0] cby_1__1__78_left_grid_pin_7_;
wire [0:0] cby_1__1__78_left_grid_pin_8_;
wire [0:0] cby_1__1__78_left_grid_pin_9_;
wire [0:0] cby_1__1__78_right_grid_pin_52_;
wire [0:0] cby_1__1__79_ccff_tail;
wire [0:19] cby_1__1__79_chany_bottom_out;
wire [0:19] cby_1__1__79_chany_top_out;
wire [0:0] cby_1__1__79_left_grid_pin_0_;
wire [0:0] cby_1__1__79_left_grid_pin_10_;
wire [0:0] cby_1__1__79_left_grid_pin_11_;
wire [0:0] cby_1__1__79_left_grid_pin_12_;
wire [0:0] cby_1__1__79_left_grid_pin_13_;
wire [0:0] cby_1__1__79_left_grid_pin_14_;
wire [0:0] cby_1__1__79_left_grid_pin_15_;
wire [0:0] cby_1__1__79_left_grid_pin_1_;
wire [0:0] cby_1__1__79_left_grid_pin_2_;
wire [0:0] cby_1__1__79_left_grid_pin_3_;
wire [0:0] cby_1__1__79_left_grid_pin_4_;
wire [0:0] cby_1__1__79_left_grid_pin_5_;
wire [0:0] cby_1__1__79_left_grid_pin_6_;
wire [0:0] cby_1__1__79_left_grid_pin_7_;
wire [0:0] cby_1__1__79_left_grid_pin_8_;
wire [0:0] cby_1__1__79_left_grid_pin_9_;
wire [0:0] cby_1__1__79_right_grid_pin_52_;
wire [0:0] cby_1__1__7_ccff_tail;
wire [0:19] cby_1__1__7_chany_bottom_out;
wire [0:19] cby_1__1__7_chany_top_out;
wire [0:0] cby_1__1__7_left_grid_pin_0_;
wire [0:0] cby_1__1__7_left_grid_pin_10_;
wire [0:0] cby_1__1__7_left_grid_pin_11_;
wire [0:0] cby_1__1__7_left_grid_pin_12_;
wire [0:0] cby_1__1__7_left_grid_pin_13_;
wire [0:0] cby_1__1__7_left_grid_pin_14_;
wire [0:0] cby_1__1__7_left_grid_pin_15_;
wire [0:0] cby_1__1__7_left_grid_pin_1_;
wire [0:0] cby_1__1__7_left_grid_pin_2_;
wire [0:0] cby_1__1__7_left_grid_pin_3_;
wire [0:0] cby_1__1__7_left_grid_pin_4_;
wire [0:0] cby_1__1__7_left_grid_pin_5_;
wire [0:0] cby_1__1__7_left_grid_pin_6_;
wire [0:0] cby_1__1__7_left_grid_pin_7_;
wire [0:0] cby_1__1__7_left_grid_pin_8_;
wire [0:0] cby_1__1__7_left_grid_pin_9_;
wire [0:0] cby_1__1__7_right_grid_pin_52_;
wire [0:0] cby_1__1__80_ccff_tail;
wire [0:19] cby_1__1__80_chany_bottom_out;
wire [0:19] cby_1__1__80_chany_top_out;
wire [0:0] cby_1__1__80_left_grid_pin_0_;
wire [0:0] cby_1__1__80_left_grid_pin_10_;
wire [0:0] cby_1__1__80_left_grid_pin_11_;
wire [0:0] cby_1__1__80_left_grid_pin_12_;
wire [0:0] cby_1__1__80_left_grid_pin_13_;
wire [0:0] cby_1__1__80_left_grid_pin_14_;
wire [0:0] cby_1__1__80_left_grid_pin_15_;
wire [0:0] cby_1__1__80_left_grid_pin_1_;
wire [0:0] cby_1__1__80_left_grid_pin_2_;
wire [0:0] cby_1__1__80_left_grid_pin_3_;
wire [0:0] cby_1__1__80_left_grid_pin_4_;
wire [0:0] cby_1__1__80_left_grid_pin_5_;
wire [0:0] cby_1__1__80_left_grid_pin_6_;
wire [0:0] cby_1__1__80_left_grid_pin_7_;
wire [0:0] cby_1__1__80_left_grid_pin_8_;
wire [0:0] cby_1__1__80_left_grid_pin_9_;
wire [0:0] cby_1__1__80_right_grid_pin_52_;
wire [0:0] cby_1__1__81_ccff_tail;
wire [0:19] cby_1__1__81_chany_bottom_out;
wire [0:19] cby_1__1__81_chany_top_out;
wire [0:0] cby_1__1__81_left_grid_pin_0_;
wire [0:0] cby_1__1__81_left_grid_pin_10_;
wire [0:0] cby_1__1__81_left_grid_pin_11_;
wire [0:0] cby_1__1__81_left_grid_pin_12_;
wire [0:0] cby_1__1__81_left_grid_pin_13_;
wire [0:0] cby_1__1__81_left_grid_pin_14_;
wire [0:0] cby_1__1__81_left_grid_pin_15_;
wire [0:0] cby_1__1__81_left_grid_pin_1_;
wire [0:0] cby_1__1__81_left_grid_pin_2_;
wire [0:0] cby_1__1__81_left_grid_pin_3_;
wire [0:0] cby_1__1__81_left_grid_pin_4_;
wire [0:0] cby_1__1__81_left_grid_pin_5_;
wire [0:0] cby_1__1__81_left_grid_pin_6_;
wire [0:0] cby_1__1__81_left_grid_pin_7_;
wire [0:0] cby_1__1__81_left_grid_pin_8_;
wire [0:0] cby_1__1__81_left_grid_pin_9_;
wire [0:0] cby_1__1__81_right_grid_pin_52_;
wire [0:0] cby_1__1__82_ccff_tail;
wire [0:19] cby_1__1__82_chany_bottom_out;
wire [0:19] cby_1__1__82_chany_top_out;
wire [0:0] cby_1__1__82_left_grid_pin_0_;
wire [0:0] cby_1__1__82_left_grid_pin_10_;
wire [0:0] cby_1__1__82_left_grid_pin_11_;
wire [0:0] cby_1__1__82_left_grid_pin_12_;
wire [0:0] cby_1__1__82_left_grid_pin_13_;
wire [0:0] cby_1__1__82_left_grid_pin_14_;
wire [0:0] cby_1__1__82_left_grid_pin_15_;
wire [0:0] cby_1__1__82_left_grid_pin_1_;
wire [0:0] cby_1__1__82_left_grid_pin_2_;
wire [0:0] cby_1__1__82_left_grid_pin_3_;
wire [0:0] cby_1__1__82_left_grid_pin_4_;
wire [0:0] cby_1__1__82_left_grid_pin_5_;
wire [0:0] cby_1__1__82_left_grid_pin_6_;
wire [0:0] cby_1__1__82_left_grid_pin_7_;
wire [0:0] cby_1__1__82_left_grid_pin_8_;
wire [0:0] cby_1__1__82_left_grid_pin_9_;
wire [0:0] cby_1__1__82_right_grid_pin_52_;
wire [0:0] cby_1__1__83_ccff_tail;
wire [0:19] cby_1__1__83_chany_bottom_out;
wire [0:19] cby_1__1__83_chany_top_out;
wire [0:0] cby_1__1__83_left_grid_pin_0_;
wire [0:0] cby_1__1__83_left_grid_pin_10_;
wire [0:0] cby_1__1__83_left_grid_pin_11_;
wire [0:0] cby_1__1__83_left_grid_pin_12_;
wire [0:0] cby_1__1__83_left_grid_pin_13_;
wire [0:0] cby_1__1__83_left_grid_pin_14_;
wire [0:0] cby_1__1__83_left_grid_pin_15_;
wire [0:0] cby_1__1__83_left_grid_pin_1_;
wire [0:0] cby_1__1__83_left_grid_pin_2_;
wire [0:0] cby_1__1__83_left_grid_pin_3_;
wire [0:0] cby_1__1__83_left_grid_pin_4_;
wire [0:0] cby_1__1__83_left_grid_pin_5_;
wire [0:0] cby_1__1__83_left_grid_pin_6_;
wire [0:0] cby_1__1__83_left_grid_pin_7_;
wire [0:0] cby_1__1__83_left_grid_pin_8_;
wire [0:0] cby_1__1__83_left_grid_pin_9_;
wire [0:0] cby_1__1__83_right_grid_pin_52_;
wire [0:0] cby_1__1__84_ccff_tail;
wire [0:19] cby_1__1__84_chany_bottom_out;
wire [0:19] cby_1__1__84_chany_top_out;
wire [0:0] cby_1__1__84_left_grid_pin_0_;
wire [0:0] cby_1__1__84_left_grid_pin_10_;
wire [0:0] cby_1__1__84_left_grid_pin_11_;
wire [0:0] cby_1__1__84_left_grid_pin_12_;
wire [0:0] cby_1__1__84_left_grid_pin_13_;
wire [0:0] cby_1__1__84_left_grid_pin_14_;
wire [0:0] cby_1__1__84_left_grid_pin_15_;
wire [0:0] cby_1__1__84_left_grid_pin_1_;
wire [0:0] cby_1__1__84_left_grid_pin_2_;
wire [0:0] cby_1__1__84_left_grid_pin_3_;
wire [0:0] cby_1__1__84_left_grid_pin_4_;
wire [0:0] cby_1__1__84_left_grid_pin_5_;
wire [0:0] cby_1__1__84_left_grid_pin_6_;
wire [0:0] cby_1__1__84_left_grid_pin_7_;
wire [0:0] cby_1__1__84_left_grid_pin_8_;
wire [0:0] cby_1__1__84_left_grid_pin_9_;
wire [0:0] cby_1__1__84_right_grid_pin_52_;
wire [0:0] cby_1__1__85_ccff_tail;
wire [0:19] cby_1__1__85_chany_bottom_out;
wire [0:19] cby_1__1__85_chany_top_out;
wire [0:0] cby_1__1__85_left_grid_pin_0_;
wire [0:0] cby_1__1__85_left_grid_pin_10_;
wire [0:0] cby_1__1__85_left_grid_pin_11_;
wire [0:0] cby_1__1__85_left_grid_pin_12_;
wire [0:0] cby_1__1__85_left_grid_pin_13_;
wire [0:0] cby_1__1__85_left_grid_pin_14_;
wire [0:0] cby_1__1__85_left_grid_pin_15_;
wire [0:0] cby_1__1__85_left_grid_pin_1_;
wire [0:0] cby_1__1__85_left_grid_pin_2_;
wire [0:0] cby_1__1__85_left_grid_pin_3_;
wire [0:0] cby_1__1__85_left_grid_pin_4_;
wire [0:0] cby_1__1__85_left_grid_pin_5_;
wire [0:0] cby_1__1__85_left_grid_pin_6_;
wire [0:0] cby_1__1__85_left_grid_pin_7_;
wire [0:0] cby_1__1__85_left_grid_pin_8_;
wire [0:0] cby_1__1__85_left_grid_pin_9_;
wire [0:0] cby_1__1__85_right_grid_pin_52_;
wire [0:0] cby_1__1__86_ccff_tail;
wire [0:19] cby_1__1__86_chany_bottom_out;
wire [0:19] cby_1__1__86_chany_top_out;
wire [0:0] cby_1__1__86_left_grid_pin_0_;
wire [0:0] cby_1__1__86_left_grid_pin_10_;
wire [0:0] cby_1__1__86_left_grid_pin_11_;
wire [0:0] cby_1__1__86_left_grid_pin_12_;
wire [0:0] cby_1__1__86_left_grid_pin_13_;
wire [0:0] cby_1__1__86_left_grid_pin_14_;
wire [0:0] cby_1__1__86_left_grid_pin_15_;
wire [0:0] cby_1__1__86_left_grid_pin_1_;
wire [0:0] cby_1__1__86_left_grid_pin_2_;
wire [0:0] cby_1__1__86_left_grid_pin_3_;
wire [0:0] cby_1__1__86_left_grid_pin_4_;
wire [0:0] cby_1__1__86_left_grid_pin_5_;
wire [0:0] cby_1__1__86_left_grid_pin_6_;
wire [0:0] cby_1__1__86_left_grid_pin_7_;
wire [0:0] cby_1__1__86_left_grid_pin_8_;
wire [0:0] cby_1__1__86_left_grid_pin_9_;
wire [0:0] cby_1__1__86_right_grid_pin_52_;
wire [0:0] cby_1__1__87_ccff_tail;
wire [0:19] cby_1__1__87_chany_bottom_out;
wire [0:19] cby_1__1__87_chany_top_out;
wire [0:0] cby_1__1__87_left_grid_pin_0_;
wire [0:0] cby_1__1__87_left_grid_pin_10_;
wire [0:0] cby_1__1__87_left_grid_pin_11_;
wire [0:0] cby_1__1__87_left_grid_pin_12_;
wire [0:0] cby_1__1__87_left_grid_pin_13_;
wire [0:0] cby_1__1__87_left_grid_pin_14_;
wire [0:0] cby_1__1__87_left_grid_pin_15_;
wire [0:0] cby_1__1__87_left_grid_pin_1_;
wire [0:0] cby_1__1__87_left_grid_pin_2_;
wire [0:0] cby_1__1__87_left_grid_pin_3_;
wire [0:0] cby_1__1__87_left_grid_pin_4_;
wire [0:0] cby_1__1__87_left_grid_pin_5_;
wire [0:0] cby_1__1__87_left_grid_pin_6_;
wire [0:0] cby_1__1__87_left_grid_pin_7_;
wire [0:0] cby_1__1__87_left_grid_pin_8_;
wire [0:0] cby_1__1__87_left_grid_pin_9_;
wire [0:0] cby_1__1__87_right_grid_pin_52_;
wire [0:0] cby_1__1__88_ccff_tail;
wire [0:19] cby_1__1__88_chany_bottom_out;
wire [0:19] cby_1__1__88_chany_top_out;
wire [0:0] cby_1__1__88_left_grid_pin_0_;
wire [0:0] cby_1__1__88_left_grid_pin_10_;
wire [0:0] cby_1__1__88_left_grid_pin_11_;
wire [0:0] cby_1__1__88_left_grid_pin_12_;
wire [0:0] cby_1__1__88_left_grid_pin_13_;
wire [0:0] cby_1__1__88_left_grid_pin_14_;
wire [0:0] cby_1__1__88_left_grid_pin_15_;
wire [0:0] cby_1__1__88_left_grid_pin_1_;
wire [0:0] cby_1__1__88_left_grid_pin_2_;
wire [0:0] cby_1__1__88_left_grid_pin_3_;
wire [0:0] cby_1__1__88_left_grid_pin_4_;
wire [0:0] cby_1__1__88_left_grid_pin_5_;
wire [0:0] cby_1__1__88_left_grid_pin_6_;
wire [0:0] cby_1__1__88_left_grid_pin_7_;
wire [0:0] cby_1__1__88_left_grid_pin_8_;
wire [0:0] cby_1__1__88_left_grid_pin_9_;
wire [0:0] cby_1__1__88_right_grid_pin_52_;
wire [0:0] cby_1__1__89_ccff_tail;
wire [0:19] cby_1__1__89_chany_bottom_out;
wire [0:19] cby_1__1__89_chany_top_out;
wire [0:0] cby_1__1__89_left_grid_pin_0_;
wire [0:0] cby_1__1__89_left_grid_pin_10_;
wire [0:0] cby_1__1__89_left_grid_pin_11_;
wire [0:0] cby_1__1__89_left_grid_pin_12_;
wire [0:0] cby_1__1__89_left_grid_pin_13_;
wire [0:0] cby_1__1__89_left_grid_pin_14_;
wire [0:0] cby_1__1__89_left_grid_pin_15_;
wire [0:0] cby_1__1__89_left_grid_pin_1_;
wire [0:0] cby_1__1__89_left_grid_pin_2_;
wire [0:0] cby_1__1__89_left_grid_pin_3_;
wire [0:0] cby_1__1__89_left_grid_pin_4_;
wire [0:0] cby_1__1__89_left_grid_pin_5_;
wire [0:0] cby_1__1__89_left_grid_pin_6_;
wire [0:0] cby_1__1__89_left_grid_pin_7_;
wire [0:0] cby_1__1__89_left_grid_pin_8_;
wire [0:0] cby_1__1__89_left_grid_pin_9_;
wire [0:0] cby_1__1__89_right_grid_pin_52_;
wire [0:0] cby_1__1__8_ccff_tail;
wire [0:19] cby_1__1__8_chany_bottom_out;
wire [0:19] cby_1__1__8_chany_top_out;
wire [0:0] cby_1__1__8_left_grid_pin_0_;
wire [0:0] cby_1__1__8_left_grid_pin_10_;
wire [0:0] cby_1__1__8_left_grid_pin_11_;
wire [0:0] cby_1__1__8_left_grid_pin_12_;
wire [0:0] cby_1__1__8_left_grid_pin_13_;
wire [0:0] cby_1__1__8_left_grid_pin_14_;
wire [0:0] cby_1__1__8_left_grid_pin_15_;
wire [0:0] cby_1__1__8_left_grid_pin_1_;
wire [0:0] cby_1__1__8_left_grid_pin_2_;
wire [0:0] cby_1__1__8_left_grid_pin_3_;
wire [0:0] cby_1__1__8_left_grid_pin_4_;
wire [0:0] cby_1__1__8_left_grid_pin_5_;
wire [0:0] cby_1__1__8_left_grid_pin_6_;
wire [0:0] cby_1__1__8_left_grid_pin_7_;
wire [0:0] cby_1__1__8_left_grid_pin_8_;
wire [0:0] cby_1__1__8_left_grid_pin_9_;
wire [0:0] cby_1__1__8_right_grid_pin_52_;
wire [0:0] cby_1__1__90_ccff_tail;
wire [0:19] cby_1__1__90_chany_bottom_out;
wire [0:19] cby_1__1__90_chany_top_out;
wire [0:0] cby_1__1__90_left_grid_pin_0_;
wire [0:0] cby_1__1__90_left_grid_pin_10_;
wire [0:0] cby_1__1__90_left_grid_pin_11_;
wire [0:0] cby_1__1__90_left_grid_pin_12_;
wire [0:0] cby_1__1__90_left_grid_pin_13_;
wire [0:0] cby_1__1__90_left_grid_pin_14_;
wire [0:0] cby_1__1__90_left_grid_pin_15_;
wire [0:0] cby_1__1__90_left_grid_pin_1_;
wire [0:0] cby_1__1__90_left_grid_pin_2_;
wire [0:0] cby_1__1__90_left_grid_pin_3_;
wire [0:0] cby_1__1__90_left_grid_pin_4_;
wire [0:0] cby_1__1__90_left_grid_pin_5_;
wire [0:0] cby_1__1__90_left_grid_pin_6_;
wire [0:0] cby_1__1__90_left_grid_pin_7_;
wire [0:0] cby_1__1__90_left_grid_pin_8_;
wire [0:0] cby_1__1__90_left_grid_pin_9_;
wire [0:0] cby_1__1__90_right_grid_pin_52_;
wire [0:0] cby_1__1__91_ccff_tail;
wire [0:19] cby_1__1__91_chany_bottom_out;
wire [0:19] cby_1__1__91_chany_top_out;
wire [0:0] cby_1__1__91_left_grid_pin_0_;
wire [0:0] cby_1__1__91_left_grid_pin_10_;
wire [0:0] cby_1__1__91_left_grid_pin_11_;
wire [0:0] cby_1__1__91_left_grid_pin_12_;
wire [0:0] cby_1__1__91_left_grid_pin_13_;
wire [0:0] cby_1__1__91_left_grid_pin_14_;
wire [0:0] cby_1__1__91_left_grid_pin_15_;
wire [0:0] cby_1__1__91_left_grid_pin_1_;
wire [0:0] cby_1__1__91_left_grid_pin_2_;
wire [0:0] cby_1__1__91_left_grid_pin_3_;
wire [0:0] cby_1__1__91_left_grid_pin_4_;
wire [0:0] cby_1__1__91_left_grid_pin_5_;
wire [0:0] cby_1__1__91_left_grid_pin_6_;
wire [0:0] cby_1__1__91_left_grid_pin_7_;
wire [0:0] cby_1__1__91_left_grid_pin_8_;
wire [0:0] cby_1__1__91_left_grid_pin_9_;
wire [0:0] cby_1__1__91_right_grid_pin_52_;
wire [0:0] cby_1__1__92_ccff_tail;
wire [0:19] cby_1__1__92_chany_bottom_out;
wire [0:19] cby_1__1__92_chany_top_out;
wire [0:0] cby_1__1__92_left_grid_pin_0_;
wire [0:0] cby_1__1__92_left_grid_pin_10_;
wire [0:0] cby_1__1__92_left_grid_pin_11_;
wire [0:0] cby_1__1__92_left_grid_pin_12_;
wire [0:0] cby_1__1__92_left_grid_pin_13_;
wire [0:0] cby_1__1__92_left_grid_pin_14_;
wire [0:0] cby_1__1__92_left_grid_pin_15_;
wire [0:0] cby_1__1__92_left_grid_pin_1_;
wire [0:0] cby_1__1__92_left_grid_pin_2_;
wire [0:0] cby_1__1__92_left_grid_pin_3_;
wire [0:0] cby_1__1__92_left_grid_pin_4_;
wire [0:0] cby_1__1__92_left_grid_pin_5_;
wire [0:0] cby_1__1__92_left_grid_pin_6_;
wire [0:0] cby_1__1__92_left_grid_pin_7_;
wire [0:0] cby_1__1__92_left_grid_pin_8_;
wire [0:0] cby_1__1__92_left_grid_pin_9_;
wire [0:0] cby_1__1__92_right_grid_pin_52_;
wire [0:0] cby_1__1__93_ccff_tail;
wire [0:19] cby_1__1__93_chany_bottom_out;
wire [0:19] cby_1__1__93_chany_top_out;
wire [0:0] cby_1__1__93_left_grid_pin_0_;
wire [0:0] cby_1__1__93_left_grid_pin_10_;
wire [0:0] cby_1__1__93_left_grid_pin_11_;
wire [0:0] cby_1__1__93_left_grid_pin_12_;
wire [0:0] cby_1__1__93_left_grid_pin_13_;
wire [0:0] cby_1__1__93_left_grid_pin_14_;
wire [0:0] cby_1__1__93_left_grid_pin_15_;
wire [0:0] cby_1__1__93_left_grid_pin_1_;
wire [0:0] cby_1__1__93_left_grid_pin_2_;
wire [0:0] cby_1__1__93_left_grid_pin_3_;
wire [0:0] cby_1__1__93_left_grid_pin_4_;
wire [0:0] cby_1__1__93_left_grid_pin_5_;
wire [0:0] cby_1__1__93_left_grid_pin_6_;
wire [0:0] cby_1__1__93_left_grid_pin_7_;
wire [0:0] cby_1__1__93_left_grid_pin_8_;
wire [0:0] cby_1__1__93_left_grid_pin_9_;
wire [0:0] cby_1__1__93_right_grid_pin_52_;
wire [0:0] cby_1__1__94_ccff_tail;
wire [0:19] cby_1__1__94_chany_bottom_out;
wire [0:19] cby_1__1__94_chany_top_out;
wire [0:0] cby_1__1__94_left_grid_pin_0_;
wire [0:0] cby_1__1__94_left_grid_pin_10_;
wire [0:0] cby_1__1__94_left_grid_pin_11_;
wire [0:0] cby_1__1__94_left_grid_pin_12_;
wire [0:0] cby_1__1__94_left_grid_pin_13_;
wire [0:0] cby_1__1__94_left_grid_pin_14_;
wire [0:0] cby_1__1__94_left_grid_pin_15_;
wire [0:0] cby_1__1__94_left_grid_pin_1_;
wire [0:0] cby_1__1__94_left_grid_pin_2_;
wire [0:0] cby_1__1__94_left_grid_pin_3_;
wire [0:0] cby_1__1__94_left_grid_pin_4_;
wire [0:0] cby_1__1__94_left_grid_pin_5_;
wire [0:0] cby_1__1__94_left_grid_pin_6_;
wire [0:0] cby_1__1__94_left_grid_pin_7_;
wire [0:0] cby_1__1__94_left_grid_pin_8_;
wire [0:0] cby_1__1__94_left_grid_pin_9_;
wire [0:0] cby_1__1__94_right_grid_pin_52_;
wire [0:0] cby_1__1__95_ccff_tail;
wire [0:19] cby_1__1__95_chany_bottom_out;
wire [0:19] cby_1__1__95_chany_top_out;
wire [0:0] cby_1__1__95_left_grid_pin_0_;
wire [0:0] cby_1__1__95_left_grid_pin_10_;
wire [0:0] cby_1__1__95_left_grid_pin_11_;
wire [0:0] cby_1__1__95_left_grid_pin_12_;
wire [0:0] cby_1__1__95_left_grid_pin_13_;
wire [0:0] cby_1__1__95_left_grid_pin_14_;
wire [0:0] cby_1__1__95_left_grid_pin_15_;
wire [0:0] cby_1__1__95_left_grid_pin_1_;
wire [0:0] cby_1__1__95_left_grid_pin_2_;
wire [0:0] cby_1__1__95_left_grid_pin_3_;
wire [0:0] cby_1__1__95_left_grid_pin_4_;
wire [0:0] cby_1__1__95_left_grid_pin_5_;
wire [0:0] cby_1__1__95_left_grid_pin_6_;
wire [0:0] cby_1__1__95_left_grid_pin_7_;
wire [0:0] cby_1__1__95_left_grid_pin_8_;
wire [0:0] cby_1__1__95_left_grid_pin_9_;
wire [0:0] cby_1__1__95_right_grid_pin_52_;
wire [0:0] cby_1__1__96_ccff_tail;
wire [0:19] cby_1__1__96_chany_bottom_out;
wire [0:19] cby_1__1__96_chany_top_out;
wire [0:0] cby_1__1__96_left_grid_pin_0_;
wire [0:0] cby_1__1__96_left_grid_pin_10_;
wire [0:0] cby_1__1__96_left_grid_pin_11_;
wire [0:0] cby_1__1__96_left_grid_pin_12_;
wire [0:0] cby_1__1__96_left_grid_pin_13_;
wire [0:0] cby_1__1__96_left_grid_pin_14_;
wire [0:0] cby_1__1__96_left_grid_pin_15_;
wire [0:0] cby_1__1__96_left_grid_pin_1_;
wire [0:0] cby_1__1__96_left_grid_pin_2_;
wire [0:0] cby_1__1__96_left_grid_pin_3_;
wire [0:0] cby_1__1__96_left_grid_pin_4_;
wire [0:0] cby_1__1__96_left_grid_pin_5_;
wire [0:0] cby_1__1__96_left_grid_pin_6_;
wire [0:0] cby_1__1__96_left_grid_pin_7_;
wire [0:0] cby_1__1__96_left_grid_pin_8_;
wire [0:0] cby_1__1__96_left_grid_pin_9_;
wire [0:0] cby_1__1__96_right_grid_pin_52_;
wire [0:0] cby_1__1__97_ccff_tail;
wire [0:19] cby_1__1__97_chany_bottom_out;
wire [0:19] cby_1__1__97_chany_top_out;
wire [0:0] cby_1__1__97_left_grid_pin_0_;
wire [0:0] cby_1__1__97_left_grid_pin_10_;
wire [0:0] cby_1__1__97_left_grid_pin_11_;
wire [0:0] cby_1__1__97_left_grid_pin_12_;
wire [0:0] cby_1__1__97_left_grid_pin_13_;
wire [0:0] cby_1__1__97_left_grid_pin_14_;
wire [0:0] cby_1__1__97_left_grid_pin_15_;
wire [0:0] cby_1__1__97_left_grid_pin_1_;
wire [0:0] cby_1__1__97_left_grid_pin_2_;
wire [0:0] cby_1__1__97_left_grid_pin_3_;
wire [0:0] cby_1__1__97_left_grid_pin_4_;
wire [0:0] cby_1__1__97_left_grid_pin_5_;
wire [0:0] cby_1__1__97_left_grid_pin_6_;
wire [0:0] cby_1__1__97_left_grid_pin_7_;
wire [0:0] cby_1__1__97_left_grid_pin_8_;
wire [0:0] cby_1__1__97_left_grid_pin_9_;
wire [0:0] cby_1__1__97_right_grid_pin_52_;
wire [0:0] cby_1__1__98_ccff_tail;
wire [0:19] cby_1__1__98_chany_bottom_out;
wire [0:19] cby_1__1__98_chany_top_out;
wire [0:0] cby_1__1__98_left_grid_pin_0_;
wire [0:0] cby_1__1__98_left_grid_pin_10_;
wire [0:0] cby_1__1__98_left_grid_pin_11_;
wire [0:0] cby_1__1__98_left_grid_pin_12_;
wire [0:0] cby_1__1__98_left_grid_pin_13_;
wire [0:0] cby_1__1__98_left_grid_pin_14_;
wire [0:0] cby_1__1__98_left_grid_pin_15_;
wire [0:0] cby_1__1__98_left_grid_pin_1_;
wire [0:0] cby_1__1__98_left_grid_pin_2_;
wire [0:0] cby_1__1__98_left_grid_pin_3_;
wire [0:0] cby_1__1__98_left_grid_pin_4_;
wire [0:0] cby_1__1__98_left_grid_pin_5_;
wire [0:0] cby_1__1__98_left_grid_pin_6_;
wire [0:0] cby_1__1__98_left_grid_pin_7_;
wire [0:0] cby_1__1__98_left_grid_pin_8_;
wire [0:0] cby_1__1__98_left_grid_pin_9_;
wire [0:0] cby_1__1__98_right_grid_pin_52_;
wire [0:0] cby_1__1__99_ccff_tail;
wire [0:19] cby_1__1__99_chany_bottom_out;
wire [0:19] cby_1__1__99_chany_top_out;
wire [0:0] cby_1__1__99_left_grid_pin_0_;
wire [0:0] cby_1__1__99_left_grid_pin_10_;
wire [0:0] cby_1__1__99_left_grid_pin_11_;
wire [0:0] cby_1__1__99_left_grid_pin_12_;
wire [0:0] cby_1__1__99_left_grid_pin_13_;
wire [0:0] cby_1__1__99_left_grid_pin_14_;
wire [0:0] cby_1__1__99_left_grid_pin_15_;
wire [0:0] cby_1__1__99_left_grid_pin_1_;
wire [0:0] cby_1__1__99_left_grid_pin_2_;
wire [0:0] cby_1__1__99_left_grid_pin_3_;
wire [0:0] cby_1__1__99_left_grid_pin_4_;
wire [0:0] cby_1__1__99_left_grid_pin_5_;
wire [0:0] cby_1__1__99_left_grid_pin_6_;
wire [0:0] cby_1__1__99_left_grid_pin_7_;
wire [0:0] cby_1__1__99_left_grid_pin_8_;
wire [0:0] cby_1__1__99_left_grid_pin_9_;
wire [0:0] cby_1__1__99_right_grid_pin_52_;
wire [0:0] cby_1__1__9_ccff_tail;
wire [0:19] cby_1__1__9_chany_bottom_out;
wire [0:19] cby_1__1__9_chany_top_out;
wire [0:0] cby_1__1__9_left_grid_pin_0_;
wire [0:0] cby_1__1__9_left_grid_pin_10_;
wire [0:0] cby_1__1__9_left_grid_pin_11_;
wire [0:0] cby_1__1__9_left_grid_pin_12_;
wire [0:0] cby_1__1__9_left_grid_pin_13_;
wire [0:0] cby_1__1__9_left_grid_pin_14_;
wire [0:0] cby_1__1__9_left_grid_pin_15_;
wire [0:0] cby_1__1__9_left_grid_pin_1_;
wire [0:0] cby_1__1__9_left_grid_pin_2_;
wire [0:0] cby_1__1__9_left_grid_pin_3_;
wire [0:0] cby_1__1__9_left_grid_pin_4_;
wire [0:0] cby_1__1__9_left_grid_pin_5_;
wire [0:0] cby_1__1__9_left_grid_pin_6_;
wire [0:0] cby_1__1__9_left_grid_pin_7_;
wire [0:0] cby_1__1__9_left_grid_pin_8_;
wire [0:0] cby_1__1__9_left_grid_pin_9_;
wire [0:0] cby_1__1__9_right_grid_pin_52_;
wire [0:0] direct_interc_0_out;
wire [0:0] direct_interc_100_out;
wire [0:0] direct_interc_101_out;
wire [0:0] direct_interc_102_out;
wire [0:0] direct_interc_103_out;
wire [0:0] direct_interc_104_out;
wire [0:0] direct_interc_105_out;
wire [0:0] direct_interc_106_out;
wire [0:0] direct_interc_107_out;
wire [0:0] direct_interc_108_out;
wire [0:0] direct_interc_109_out;
wire [0:0] direct_interc_10_out;
wire [0:0] direct_interc_110_out;
wire [0:0] direct_interc_111_out;
wire [0:0] direct_interc_112_out;
wire [0:0] direct_interc_113_out;
wire [0:0] direct_interc_114_out;
wire [0:0] direct_interc_115_out;
wire [0:0] direct_interc_116_out;
wire [0:0] direct_interc_117_out;
wire [0:0] direct_interc_118_out;
wire [0:0] direct_interc_119_out;
wire [0:0] direct_interc_11_out;
wire [0:0] direct_interc_120_out;
wire [0:0] direct_interc_121_out;
wire [0:0] direct_interc_122_out;
wire [0:0] direct_interc_123_out;
wire [0:0] direct_interc_124_out;
wire [0:0] direct_interc_125_out;
wire [0:0] direct_interc_126_out;
wire [0:0] direct_interc_127_out;
wire [0:0] direct_interc_128_out;
wire [0:0] direct_interc_129_out;
wire [0:0] direct_interc_12_out;
wire [0:0] direct_interc_130_out;
wire [0:0] direct_interc_131_out;
wire [0:0] direct_interc_132_out;
wire [0:0] direct_interc_133_out;
wire [0:0] direct_interc_134_out;
wire [0:0] direct_interc_135_out;
wire [0:0] direct_interc_136_out;
wire [0:0] direct_interc_137_out;
wire [0:0] direct_interc_138_out;
wire [0:0] direct_interc_139_out;
wire [0:0] direct_interc_13_out;
wire [0:0] direct_interc_140_out;
wire [0:0] direct_interc_141_out;
wire [0:0] direct_interc_142_out;
wire [0:0] direct_interc_143_out;
wire [0:0] direct_interc_144_out;
wire [0:0] direct_interc_145_out;
wire [0:0] direct_interc_146_out;
wire [0:0] direct_interc_147_out;
wire [0:0] direct_interc_148_out;
wire [0:0] direct_interc_149_out;
wire [0:0] direct_interc_14_out;
wire [0:0] direct_interc_150_out;
wire [0:0] direct_interc_151_out;
wire [0:0] direct_interc_152_out;
wire [0:0] direct_interc_153_out;
wire [0:0] direct_interc_154_out;
wire [0:0] direct_interc_155_out;
wire [0:0] direct_interc_156_out;
wire [0:0] direct_interc_157_out;
wire [0:0] direct_interc_158_out;
wire [0:0] direct_interc_159_out;
wire [0:0] direct_interc_15_out;
wire [0:0] direct_interc_160_out;
wire [0:0] direct_interc_161_out;
wire [0:0] direct_interc_162_out;
wire [0:0] direct_interc_163_out;
wire [0:0] direct_interc_164_out;
wire [0:0] direct_interc_165_out;
wire [0:0] direct_interc_166_out;
wire [0:0] direct_interc_167_out;
wire [0:0] direct_interc_168_out;
wire [0:0] direct_interc_169_out;
wire [0:0] direct_interc_16_out;
wire [0:0] direct_interc_170_out;
wire [0:0] direct_interc_171_out;
wire [0:0] direct_interc_172_out;
wire [0:0] direct_interc_173_out;
wire [0:0] direct_interc_174_out;
wire [0:0] direct_interc_175_out;
wire [0:0] direct_interc_176_out;
wire [0:0] direct_interc_177_out;
wire [0:0] direct_interc_178_out;
wire [0:0] direct_interc_179_out;
wire [0:0] direct_interc_17_out;
wire [0:0] direct_interc_180_out;
wire [0:0] direct_interc_181_out;
wire [0:0] direct_interc_182_out;
wire [0:0] direct_interc_183_out;
wire [0:0] direct_interc_184_out;
wire [0:0] direct_interc_185_out;
wire [0:0] direct_interc_186_out;
wire [0:0] direct_interc_187_out;
wire [0:0] direct_interc_188_out;
wire [0:0] direct_interc_189_out;
wire [0:0] direct_interc_18_out;
wire [0:0] direct_interc_190_out;
wire [0:0] direct_interc_191_out;
wire [0:0] direct_interc_192_out;
wire [0:0] direct_interc_193_out;
wire [0:0] direct_interc_194_out;
wire [0:0] direct_interc_195_out;
wire [0:0] direct_interc_196_out;
wire [0:0] direct_interc_197_out;
wire [0:0] direct_interc_198_out;
wire [0:0] direct_interc_199_out;
wire [0:0] direct_interc_19_out;
wire [0:0] direct_interc_1_out;
wire [0:0] direct_interc_200_out;
wire [0:0] direct_interc_201_out;
wire [0:0] direct_interc_202_out;
wire [0:0] direct_interc_203_out;
wire [0:0] direct_interc_204_out;
wire [0:0] direct_interc_205_out;
wire [0:0] direct_interc_206_out;
wire [0:0] direct_interc_207_out;
wire [0:0] direct_interc_208_out;
wire [0:0] direct_interc_209_out;
wire [0:0] direct_interc_20_out;
wire [0:0] direct_interc_210_out;
wire [0:0] direct_interc_211_out;
wire [0:0] direct_interc_212_out;
wire [0:0] direct_interc_213_out;
wire [0:0] direct_interc_214_out;
wire [0:0] direct_interc_215_out;
wire [0:0] direct_interc_216_out;
wire [0:0] direct_interc_217_out;
wire [0:0] direct_interc_218_out;
wire [0:0] direct_interc_219_out;
wire [0:0] direct_interc_21_out;
wire [0:0] direct_interc_220_out;
wire [0:0] direct_interc_221_out;
wire [0:0] direct_interc_222_out;
wire [0:0] direct_interc_223_out;
wire [0:0] direct_interc_224_out;
wire [0:0] direct_interc_225_out;
wire [0:0] direct_interc_226_out;
wire [0:0] direct_interc_227_out;
wire [0:0] direct_interc_228_out;
wire [0:0] direct_interc_229_out;
wire [0:0] direct_interc_22_out;
wire [0:0] direct_interc_230_out;
wire [0:0] direct_interc_231_out;
wire [0:0] direct_interc_232_out;
wire [0:0] direct_interc_233_out;
wire [0:0] direct_interc_234_out;
wire [0:0] direct_interc_235_out;
wire [0:0] direct_interc_236_out;
wire [0:0] direct_interc_237_out;
wire [0:0] direct_interc_238_out;
wire [0:0] direct_interc_239_out;
wire [0:0] direct_interc_23_out;
wire [0:0] direct_interc_240_out;
wire [0:0] direct_interc_241_out;
wire [0:0] direct_interc_242_out;
wire [0:0] direct_interc_243_out;
wire [0:0] direct_interc_244_out;
wire [0:0] direct_interc_245_out;
wire [0:0] direct_interc_246_out;
wire [0:0] direct_interc_247_out;
wire [0:0] direct_interc_248_out;
wire [0:0] direct_interc_249_out;
wire [0:0] direct_interc_24_out;
wire [0:0] direct_interc_250_out;
wire [0:0] direct_interc_251_out;
wire [0:0] direct_interc_252_out;
wire [0:0] direct_interc_253_out;
wire [0:0] direct_interc_254_out;
wire [0:0] direct_interc_255_out;
wire [0:0] direct_interc_256_out;
wire [0:0] direct_interc_257_out;
wire [0:0] direct_interc_258_out;
wire [0:0] direct_interc_259_out;
wire [0:0] direct_interc_25_out;
wire [0:0] direct_interc_260_out;
wire [0:0] direct_interc_261_out;
wire [0:0] direct_interc_262_out;
wire [0:0] direct_interc_263_out;
wire [0:0] direct_interc_264_out;
wire [0:0] direct_interc_265_out;
wire [0:0] direct_interc_266_out;
wire [0:0] direct_interc_267_out;
wire [0:0] direct_interc_268_out;
wire [0:0] direct_interc_269_out;
wire [0:0] direct_interc_26_out;
wire [0:0] direct_interc_270_out;
wire [0:0] direct_interc_271_out;
wire [0:0] direct_interc_272_out;
wire [0:0] direct_interc_273_out;
wire [0:0] direct_interc_274_out;
wire [0:0] direct_interc_275_out;
wire [0:0] direct_interc_276_out;
wire [0:0] direct_interc_277_out;
wire [0:0] direct_interc_278_out;
wire [0:0] direct_interc_279_out;
wire [0:0] direct_interc_27_out;
wire [0:0] direct_interc_280_out;
wire [0:0] direct_interc_281_out;
wire [0:0] direct_interc_282_out;
wire [0:0] direct_interc_283_out;
wire [0:0] direct_interc_284_out;
wire [0:0] direct_interc_285_out;
wire [0:0] direct_interc_28_out;
wire [0:0] direct_interc_29_out;
wire [0:0] direct_interc_2_out;
wire [0:0] direct_interc_30_out;
wire [0:0] direct_interc_31_out;
wire [0:0] direct_interc_32_out;
wire [0:0] direct_interc_33_out;
wire [0:0] direct_interc_34_out;
wire [0:0] direct_interc_35_out;
wire [0:0] direct_interc_36_out;
wire [0:0] direct_interc_37_out;
wire [0:0] direct_interc_38_out;
wire [0:0] direct_interc_39_out;
wire [0:0] direct_interc_3_out;
wire [0:0] direct_interc_40_out;
wire [0:0] direct_interc_41_out;
wire [0:0] direct_interc_42_out;
wire [0:0] direct_interc_43_out;
wire [0:0] direct_interc_44_out;
wire [0:0] direct_interc_45_out;
wire [0:0] direct_interc_46_out;
wire [0:0] direct_interc_47_out;
wire [0:0] direct_interc_48_out;
wire [0:0] direct_interc_49_out;
wire [0:0] direct_interc_4_out;
wire [0:0] direct_interc_50_out;
wire [0:0] direct_interc_51_out;
wire [0:0] direct_interc_52_out;
wire [0:0] direct_interc_53_out;
wire [0:0] direct_interc_54_out;
wire [0:0] direct_interc_55_out;
wire [0:0] direct_interc_56_out;
wire [0:0] direct_interc_57_out;
wire [0:0] direct_interc_58_out;
wire [0:0] direct_interc_59_out;
wire [0:0] direct_interc_5_out;
wire [0:0] direct_interc_60_out;
wire [0:0] direct_interc_61_out;
wire [0:0] direct_interc_62_out;
wire [0:0] direct_interc_63_out;
wire [0:0] direct_interc_64_out;
wire [0:0] direct_interc_65_out;
wire [0:0] direct_interc_66_out;
wire [0:0] direct_interc_67_out;
wire [0:0] direct_interc_68_out;
wire [0:0] direct_interc_69_out;
wire [0:0] direct_interc_6_out;
wire [0:0] direct_interc_70_out;
wire [0:0] direct_interc_71_out;
wire [0:0] direct_interc_72_out;
wire [0:0] direct_interc_73_out;
wire [0:0] direct_interc_74_out;
wire [0:0] direct_interc_75_out;
wire [0:0] direct_interc_76_out;
wire [0:0] direct_interc_77_out;
wire [0:0] direct_interc_78_out;
wire [0:0] direct_interc_79_out;
wire [0:0] direct_interc_7_out;
wire [0:0] direct_interc_80_out;
wire [0:0] direct_interc_81_out;
wire [0:0] direct_interc_82_out;
wire [0:0] direct_interc_83_out;
wire [0:0] direct_interc_84_out;
wire [0:0] direct_interc_85_out;
wire [0:0] direct_interc_86_out;
wire [0:0] direct_interc_87_out;
wire [0:0] direct_interc_88_out;
wire [0:0] direct_interc_89_out;
wire [0:0] direct_interc_8_out;
wire [0:0] direct_interc_90_out;
wire [0:0] direct_interc_91_out;
wire [0:0] direct_interc_92_out;
wire [0:0] direct_interc_93_out;
wire [0:0] direct_interc_94_out;
wire [0:0] direct_interc_95_out;
wire [0:0] direct_interc_96_out;
wire [0:0] direct_interc_97_out;
wire [0:0] direct_interc_98_out;
wire [0:0] direct_interc_99_out;
wire [0:0] direct_interc_9_out;
wire [0:0] grid_clb_0_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_0_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_0_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_0_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_0_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_0_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_0_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_0_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_0_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_0_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_0_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_0_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_0_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_0_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_0_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_0_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_0_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_0_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_0_ccff_tail;
wire [0:0] grid_clb_0_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_0_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_0_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_0_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_0_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_0_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_0_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_0_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_0_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_0_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_0_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_0_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_0_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_0_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_0_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_0_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_100_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_100_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_100_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_100_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_100_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_100_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_100_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_100_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_100_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_100_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_100_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_100_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_100_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_100_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_100_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_100_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_100_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_100_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_100_ccff_tail;
wire [0:0] grid_clb_100_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_100_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_100_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_100_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_100_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_100_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_100_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_100_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_100_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_100_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_100_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_100_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_100_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_100_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_100_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_100_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_101_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_101_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_101_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_101_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_101_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_101_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_101_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_101_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_101_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_101_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_101_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_101_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_101_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_101_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_101_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_101_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_101_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_101_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_101_ccff_tail;
wire [0:0] grid_clb_101_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_101_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_101_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_101_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_101_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_101_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_101_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_101_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_101_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_101_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_101_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_101_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_101_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_101_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_101_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_101_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_102_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_102_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_102_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_102_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_102_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_102_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_102_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_102_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_102_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_102_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_102_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_102_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_102_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_102_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_102_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_102_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_102_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_102_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_102_ccff_tail;
wire [0:0] grid_clb_102_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_102_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_102_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_102_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_102_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_102_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_102_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_102_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_102_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_102_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_102_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_102_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_102_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_102_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_102_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_102_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_103_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_103_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_103_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_103_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_103_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_103_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_103_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_103_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_103_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_103_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_103_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_103_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_103_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_103_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_103_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_103_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_103_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_103_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_103_ccff_tail;
wire [0:0] grid_clb_103_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_103_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_103_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_103_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_103_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_103_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_103_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_103_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_103_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_103_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_103_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_103_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_103_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_103_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_103_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_103_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_104_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_104_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_104_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_104_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_104_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_104_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_104_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_104_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_104_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_104_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_104_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_104_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_104_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_104_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_104_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_104_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_104_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_104_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_104_ccff_tail;
wire [0:0] grid_clb_104_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_104_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_104_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_104_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_104_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_104_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_104_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_104_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_104_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_104_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_104_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_104_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_104_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_104_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_104_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_104_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_105_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_105_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_105_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_105_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_105_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_105_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_105_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_105_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_105_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_105_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_105_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_105_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_105_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_105_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_105_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_105_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_105_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_105_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_105_ccff_tail;
wire [0:0] grid_clb_105_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_105_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_105_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_105_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_105_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_105_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_105_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_105_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_105_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_105_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_105_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_105_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_105_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_105_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_105_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_105_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_106_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_106_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_106_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_106_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_106_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_106_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_106_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_106_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_106_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_106_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_106_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_106_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_106_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_106_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_106_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_106_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_106_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_106_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_106_ccff_tail;
wire [0:0] grid_clb_106_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_106_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_106_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_106_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_106_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_106_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_106_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_106_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_106_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_106_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_106_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_106_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_106_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_106_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_106_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_106_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_107_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_107_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_107_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_107_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_107_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_107_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_107_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_107_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_107_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_107_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_107_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_107_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_107_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_107_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_107_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_107_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_107_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_107_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_107_ccff_tail;
wire [0:0] grid_clb_107_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_107_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_107_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_107_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_107_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_107_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_107_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_107_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_107_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_107_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_107_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_107_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_107_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_107_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_107_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_107_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_108_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_108_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_108_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_108_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_108_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_108_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_108_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_108_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_108_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_108_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_108_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_108_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_108_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_108_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_108_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_108_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_108_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_108_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_108_ccff_tail;
wire [0:0] grid_clb_108_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_108_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_108_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_108_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_108_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_108_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_108_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_108_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_108_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_108_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_108_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_108_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_108_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_108_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_108_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_108_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_109_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_109_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_109_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_109_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_109_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_109_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_109_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_109_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_109_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_109_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_109_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_109_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_109_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_109_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_109_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_109_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_109_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_109_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_109_ccff_tail;
wire [0:0] grid_clb_109_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_109_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_109_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_109_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_109_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_109_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_109_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_109_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_109_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_109_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_109_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_109_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_109_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_109_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_109_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_109_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_10_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_10_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_10_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_10_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_10_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_10_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_10_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_10_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_10_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_10_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_10_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_10_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_10_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_10_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_10_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_10_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_10_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_10_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_10_ccff_tail;
wire [0:0] grid_clb_10_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_10_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_10_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_10_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_10_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_10_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_10_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_10_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_10_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_10_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_10_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_10_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_10_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_10_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_10_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_10_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_110_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_110_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_110_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_110_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_110_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_110_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_110_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_110_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_110_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_110_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_110_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_110_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_110_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_110_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_110_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_110_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_110_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_110_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_110_ccff_tail;
wire [0:0] grid_clb_110_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_110_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_110_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_110_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_110_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_110_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_110_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_110_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_110_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_110_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_110_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_110_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_110_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_110_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_110_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_110_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_111_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_111_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_111_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_111_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_111_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_111_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_111_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_111_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_111_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_111_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_111_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_111_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_111_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_111_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_111_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_111_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_111_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_111_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_111_ccff_tail;
wire [0:0] grid_clb_111_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_111_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_111_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_111_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_111_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_111_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_111_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_111_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_111_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_111_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_111_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_111_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_111_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_111_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_111_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_111_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_112_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_112_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_112_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_112_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_112_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_112_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_112_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_112_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_112_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_112_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_112_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_112_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_112_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_112_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_112_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_112_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_112_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_112_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_112_ccff_tail;
wire [0:0] grid_clb_112_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_112_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_112_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_112_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_112_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_112_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_112_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_112_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_112_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_112_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_112_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_112_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_112_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_112_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_112_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_112_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_113_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_113_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_113_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_113_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_113_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_113_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_113_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_113_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_113_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_113_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_113_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_113_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_113_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_113_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_113_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_113_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_113_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_113_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_113_ccff_tail;
wire [0:0] grid_clb_113_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_113_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_113_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_113_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_113_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_113_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_113_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_113_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_113_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_113_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_113_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_113_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_113_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_113_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_113_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_113_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_114_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_114_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_114_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_114_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_114_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_114_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_114_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_114_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_114_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_114_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_114_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_114_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_114_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_114_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_114_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_114_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_114_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_114_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_114_ccff_tail;
wire [0:0] grid_clb_114_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_114_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_114_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_114_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_114_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_114_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_114_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_114_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_114_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_114_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_114_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_114_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_114_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_114_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_114_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_114_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_115_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_115_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_115_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_115_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_115_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_115_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_115_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_115_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_115_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_115_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_115_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_115_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_115_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_115_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_115_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_115_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_115_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_115_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_115_ccff_tail;
wire [0:0] grid_clb_115_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_115_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_115_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_115_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_115_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_115_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_115_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_115_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_115_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_115_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_115_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_115_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_115_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_115_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_115_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_115_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_116_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_116_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_116_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_116_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_116_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_116_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_116_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_116_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_116_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_116_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_116_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_116_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_116_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_116_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_116_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_116_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_116_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_116_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_116_ccff_tail;
wire [0:0] grid_clb_116_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_116_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_116_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_116_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_116_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_116_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_116_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_116_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_116_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_116_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_116_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_116_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_116_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_116_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_116_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_116_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_117_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_117_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_117_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_117_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_117_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_117_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_117_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_117_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_117_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_117_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_117_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_117_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_117_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_117_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_117_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_117_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_117_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_117_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_117_ccff_tail;
wire [0:0] grid_clb_117_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_117_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_117_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_117_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_117_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_117_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_117_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_117_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_117_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_117_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_117_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_117_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_117_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_117_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_117_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_117_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_118_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_118_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_118_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_118_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_118_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_118_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_118_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_118_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_118_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_118_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_118_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_118_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_118_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_118_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_118_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_118_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_118_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_118_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_118_ccff_tail;
wire [0:0] grid_clb_118_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_118_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_118_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_118_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_118_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_118_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_118_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_118_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_118_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_118_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_118_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_118_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_118_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_118_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_118_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_118_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_119_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_119_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_119_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_119_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_119_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_119_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_119_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_119_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_119_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_119_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_119_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_119_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_119_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_119_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_119_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_119_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_119_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_119_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_119_ccff_tail;
wire [0:0] grid_clb_119_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_119_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_119_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_119_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_119_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_119_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_119_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_119_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_119_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_119_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_119_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_119_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_119_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_119_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_119_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_119_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_11_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_11_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_11_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_11_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_11_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_11_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_11_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_11_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_11_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_11_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_11_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_11_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_11_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_11_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_11_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_11_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_11_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_11_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_11_ccff_tail;
wire [0:0] grid_clb_11_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_11_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_11_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_11_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_11_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_11_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_11_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_11_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_11_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_11_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_11_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_11_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_11_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_11_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_11_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_11_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_120_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_120_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_120_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_120_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_120_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_120_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_120_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_120_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_120_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_120_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_120_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_120_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_120_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_120_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_120_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_120_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_120_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_120_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_120_ccff_tail;
wire [0:0] grid_clb_120_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_120_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_120_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_120_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_120_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_120_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_120_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_120_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_120_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_120_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_120_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_120_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_120_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_120_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_120_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_120_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_121_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_121_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_121_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_121_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_121_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_121_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_121_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_121_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_121_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_121_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_121_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_121_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_121_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_121_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_121_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_121_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_121_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_121_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_121_ccff_tail;
wire [0:0] grid_clb_121_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_121_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_121_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_121_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_121_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_121_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_121_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_121_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_121_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_121_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_121_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_121_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_121_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_121_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_121_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_121_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_122_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_122_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_122_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_122_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_122_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_122_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_122_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_122_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_122_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_122_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_122_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_122_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_122_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_122_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_122_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_122_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_122_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_122_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_122_ccff_tail;
wire [0:0] grid_clb_122_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_122_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_122_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_122_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_122_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_122_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_122_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_122_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_122_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_122_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_122_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_122_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_122_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_122_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_122_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_122_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_123_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_123_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_123_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_123_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_123_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_123_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_123_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_123_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_123_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_123_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_123_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_123_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_123_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_123_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_123_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_123_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_123_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_123_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_123_ccff_tail;
wire [0:0] grid_clb_123_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_123_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_123_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_123_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_123_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_123_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_123_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_123_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_123_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_123_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_123_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_123_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_123_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_123_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_123_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_123_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_124_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_124_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_124_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_124_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_124_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_124_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_124_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_124_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_124_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_124_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_124_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_124_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_124_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_124_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_124_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_124_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_124_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_124_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_124_ccff_tail;
wire [0:0] grid_clb_124_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_124_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_124_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_124_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_124_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_124_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_124_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_124_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_124_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_124_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_124_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_124_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_124_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_124_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_124_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_124_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_125_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_125_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_125_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_125_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_125_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_125_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_125_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_125_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_125_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_125_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_125_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_125_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_125_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_125_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_125_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_125_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_125_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_125_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_125_ccff_tail;
wire [0:0] grid_clb_125_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_125_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_125_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_125_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_125_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_125_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_125_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_125_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_125_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_125_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_125_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_125_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_125_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_125_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_125_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_125_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_126_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_126_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_126_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_126_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_126_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_126_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_126_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_126_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_126_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_126_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_126_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_126_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_126_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_126_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_126_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_126_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_126_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_126_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_126_ccff_tail;
wire [0:0] grid_clb_126_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_126_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_126_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_126_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_126_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_126_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_126_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_126_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_126_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_126_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_126_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_126_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_126_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_126_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_126_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_126_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_127_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_127_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_127_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_127_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_127_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_127_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_127_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_127_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_127_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_127_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_127_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_127_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_127_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_127_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_127_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_127_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_127_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_127_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_127_ccff_tail;
wire [0:0] grid_clb_127_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_127_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_127_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_127_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_127_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_127_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_127_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_127_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_127_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_127_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_127_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_127_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_127_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_127_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_127_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_127_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_128_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_128_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_128_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_128_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_128_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_128_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_128_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_128_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_128_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_128_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_128_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_128_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_128_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_128_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_128_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_128_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_128_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_128_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_128_ccff_tail;
wire [0:0] grid_clb_128_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_128_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_128_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_128_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_128_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_128_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_128_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_128_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_128_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_128_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_128_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_128_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_128_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_128_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_128_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_128_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_129_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_129_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_129_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_129_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_129_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_129_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_129_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_129_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_129_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_129_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_129_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_129_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_129_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_129_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_129_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_129_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_129_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_129_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_129_ccff_tail;
wire [0:0] grid_clb_129_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_129_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_129_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_129_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_129_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_129_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_129_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_129_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_129_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_129_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_129_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_129_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_129_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_129_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_129_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_129_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_12__1__undriven_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_12__1__undriven_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_12_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_12_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_12_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_12_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_12_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_12_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_12_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_12_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_12_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_12_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_12_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_12_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_12_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_12_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_12_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_12_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_12_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_12_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_12_ccff_tail;
wire [0:0] grid_clb_12_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_12_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_12_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_12_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_12_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_12_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_12_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_12_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_12_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_12_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_12_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_12_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_12_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_12_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_12_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_12_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_130_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_130_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_130_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_130_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_130_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_130_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_130_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_130_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_130_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_130_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_130_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_130_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_130_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_130_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_130_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_130_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_130_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_130_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_130_ccff_tail;
wire [0:0] grid_clb_130_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_130_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_130_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_130_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_130_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_130_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_130_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_130_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_130_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_130_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_130_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_130_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_130_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_130_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_130_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_130_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_131_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_131_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_131_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_131_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_131_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_131_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_131_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_131_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_131_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_131_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_131_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_131_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_131_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_131_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_131_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_131_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_131_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_131_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_131_ccff_tail;
wire [0:0] grid_clb_131_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_131_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_131_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_131_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_131_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_131_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_131_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_131_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_131_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_131_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_131_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_131_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_131_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_131_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_131_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_131_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_132_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_132_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_132_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_132_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_132_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_132_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_132_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_132_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_132_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_132_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_132_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_132_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_132_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_132_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_132_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_132_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_132_ccff_tail;
wire [0:0] grid_clb_132_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_132_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_132_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_132_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_132_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_132_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_132_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_132_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_132_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_132_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_132_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_132_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_132_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_132_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_132_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_132_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_133_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_133_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_133_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_133_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_133_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_133_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_133_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_133_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_133_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_133_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_133_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_133_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_133_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_133_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_133_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_133_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_133_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_133_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_133_ccff_tail;
wire [0:0] grid_clb_133_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_133_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_133_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_133_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_133_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_133_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_133_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_133_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_133_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_133_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_133_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_133_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_133_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_133_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_133_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_133_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_134_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_134_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_134_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_134_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_134_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_134_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_134_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_134_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_134_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_134_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_134_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_134_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_134_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_134_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_134_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_134_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_134_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_134_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_134_ccff_tail;
wire [0:0] grid_clb_134_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_134_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_134_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_134_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_134_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_134_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_134_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_134_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_134_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_134_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_134_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_134_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_134_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_134_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_134_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_134_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_135_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_135_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_135_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_135_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_135_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_135_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_135_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_135_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_135_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_135_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_135_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_135_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_135_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_135_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_135_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_135_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_135_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_135_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_135_ccff_tail;
wire [0:0] grid_clb_135_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_135_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_135_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_135_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_135_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_135_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_135_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_135_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_135_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_135_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_135_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_135_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_135_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_135_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_135_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_135_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_136_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_136_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_136_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_136_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_136_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_136_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_136_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_136_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_136_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_136_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_136_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_136_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_136_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_136_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_136_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_136_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_136_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_136_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_136_ccff_tail;
wire [0:0] grid_clb_136_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_136_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_136_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_136_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_136_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_136_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_136_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_136_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_136_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_136_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_136_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_136_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_136_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_136_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_136_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_136_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_137_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_137_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_137_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_137_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_137_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_137_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_137_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_137_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_137_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_137_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_137_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_137_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_137_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_137_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_137_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_137_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_137_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_137_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_137_ccff_tail;
wire [0:0] grid_clb_137_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_137_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_137_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_137_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_137_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_137_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_137_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_137_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_137_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_137_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_137_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_137_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_137_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_137_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_137_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_137_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_138_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_138_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_138_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_138_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_138_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_138_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_138_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_138_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_138_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_138_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_138_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_138_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_138_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_138_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_138_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_138_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_138_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_138_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_138_ccff_tail;
wire [0:0] grid_clb_138_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_138_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_138_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_138_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_138_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_138_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_138_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_138_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_138_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_138_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_138_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_138_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_138_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_138_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_138_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_138_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_139_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_139_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_139_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_139_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_139_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_139_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_139_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_139_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_139_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_139_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_139_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_139_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_139_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_139_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_139_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_139_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_139_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_139_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_139_ccff_tail;
wire [0:0] grid_clb_139_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_139_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_139_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_139_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_139_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_139_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_139_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_139_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_139_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_139_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_139_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_139_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_139_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_139_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_139_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_139_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_13_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_13_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_13_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_13_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_13_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_13_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_13_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_13_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_13_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_13_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_13_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_13_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_13_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_13_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_13_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_13_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_13_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_13_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_13_ccff_tail;
wire [0:0] grid_clb_13_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_13_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_13_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_13_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_13_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_13_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_13_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_13_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_13_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_13_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_13_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_13_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_13_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_13_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_13_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_13_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_140_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_140_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_140_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_140_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_140_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_140_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_140_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_140_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_140_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_140_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_140_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_140_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_140_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_140_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_140_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_140_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_140_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_140_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_140_ccff_tail;
wire [0:0] grid_clb_140_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_140_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_140_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_140_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_140_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_140_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_140_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_140_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_140_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_140_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_140_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_140_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_140_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_140_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_140_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_140_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_141_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_141_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_141_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_141_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_141_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_141_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_141_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_141_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_141_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_141_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_141_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_141_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_141_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_141_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_141_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_141_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_141_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_141_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_141_ccff_tail;
wire [0:0] grid_clb_141_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_141_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_141_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_141_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_141_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_141_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_141_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_141_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_141_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_141_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_141_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_141_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_141_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_141_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_141_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_141_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_142_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_142_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_142_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_142_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_142_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_142_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_142_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_142_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_142_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_142_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_142_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_142_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_142_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_142_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_142_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_142_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_142_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_142_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_142_ccff_tail;
wire [0:0] grid_clb_142_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_142_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_142_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_142_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_142_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_142_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_142_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_142_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_142_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_142_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_142_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_142_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_142_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_142_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_142_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_142_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_143_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_143_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_143_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_143_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_143_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_143_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_143_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_143_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_143_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_143_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_143_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_143_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_143_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_143_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_143_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_143_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_143_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_143_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_143_ccff_tail;
wire [0:0] grid_clb_143_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_143_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_143_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_143_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_143_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_143_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_143_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_143_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_143_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_143_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_143_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_143_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_143_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_143_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_143_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_143_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_14_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_14_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_14_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_14_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_14_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_14_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_14_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_14_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_14_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_14_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_14_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_14_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_14_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_14_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_14_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_14_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_14_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_14_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_14_ccff_tail;
wire [0:0] grid_clb_14_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_14_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_14_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_14_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_14_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_14_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_14_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_14_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_14_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_14_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_14_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_14_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_14_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_14_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_14_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_14_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_15_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_15_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_15_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_15_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_15_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_15_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_15_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_15_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_15_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_15_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_15_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_15_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_15_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_15_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_15_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_15_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_15_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_15_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_15_ccff_tail;
wire [0:0] grid_clb_15_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_15_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_15_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_15_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_15_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_15_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_15_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_15_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_15_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_15_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_15_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_15_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_15_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_15_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_15_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_15_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_16_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_16_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_16_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_16_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_16_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_16_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_16_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_16_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_16_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_16_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_16_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_16_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_16_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_16_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_16_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_16_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_16_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_16_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_16_ccff_tail;
wire [0:0] grid_clb_16_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_16_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_16_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_16_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_16_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_16_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_16_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_16_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_16_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_16_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_16_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_16_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_16_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_16_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_16_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_16_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_17_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_17_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_17_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_17_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_17_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_17_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_17_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_17_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_17_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_17_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_17_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_17_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_17_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_17_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_17_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_17_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_17_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_17_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_17_ccff_tail;
wire [0:0] grid_clb_17_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_17_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_17_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_17_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_17_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_17_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_17_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_17_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_17_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_17_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_17_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_17_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_17_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_17_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_17_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_17_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_18_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_18_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_18_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_18_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_18_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_18_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_18_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_18_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_18_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_18_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_18_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_18_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_18_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_18_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_18_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_18_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_18_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_18_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_18_ccff_tail;
wire [0:0] grid_clb_18_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_18_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_18_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_18_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_18_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_18_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_18_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_18_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_18_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_18_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_18_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_18_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_18_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_18_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_18_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_18_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_19_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_19_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_19_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_19_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_19_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_19_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_19_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_19_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_19_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_19_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_19_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_19_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_19_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_19_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_19_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_19_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_19_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_19_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_19_ccff_tail;
wire [0:0] grid_clb_19_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_19_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_19_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_19_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_19_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_19_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_19_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_19_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_19_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_19_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_19_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_19_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_19_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_19_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_19_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_19_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_1__12__undriven_top_width_0_height_0__pin_32_;
wire [0:0] grid_clb_1__12__undriven_top_width_0_height_0__pin_33_;
wire [0:0] grid_clb_1_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_1_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_1_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_1_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_1_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_1_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_1_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_1_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_1_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_1_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_1_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_1_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_1_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_1_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_1_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_1_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_1_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_1_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_1_ccff_tail;
wire [0:0] grid_clb_1_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_1_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_1_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_1_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_1_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_1_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_1_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_1_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_1_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_1_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_1_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_1_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_1_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_1_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_1_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_1_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_20_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_20_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_20_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_20_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_20_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_20_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_20_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_20_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_20_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_20_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_20_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_20_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_20_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_20_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_20_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_20_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_20_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_20_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_20_ccff_tail;
wire [0:0] grid_clb_20_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_20_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_20_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_20_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_20_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_20_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_20_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_20_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_20_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_20_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_20_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_20_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_20_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_20_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_20_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_20_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_21_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_21_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_21_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_21_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_21_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_21_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_21_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_21_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_21_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_21_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_21_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_21_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_21_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_21_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_21_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_21_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_21_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_21_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_21_ccff_tail;
wire [0:0] grid_clb_21_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_21_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_21_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_21_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_21_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_21_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_21_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_21_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_21_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_21_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_21_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_21_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_21_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_21_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_21_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_21_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_22_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_22_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_22_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_22_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_22_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_22_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_22_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_22_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_22_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_22_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_22_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_22_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_22_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_22_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_22_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_22_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_22_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_22_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_22_ccff_tail;
wire [0:0] grid_clb_22_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_22_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_22_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_22_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_22_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_22_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_22_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_22_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_22_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_22_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_22_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_22_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_22_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_22_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_22_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_22_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_23_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_23_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_23_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_23_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_23_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_23_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_23_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_23_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_23_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_23_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_23_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_23_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_23_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_23_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_23_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_23_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_23_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_23_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_23_ccff_tail;
wire [0:0] grid_clb_23_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_23_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_23_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_23_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_23_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_23_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_23_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_23_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_23_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_23_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_23_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_23_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_23_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_23_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_23_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_23_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_24_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_24_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_24_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_24_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_24_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_24_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_24_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_24_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_24_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_24_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_24_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_24_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_24_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_24_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_24_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_24_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_24_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_24_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_24_ccff_tail;
wire [0:0] grid_clb_24_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_24_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_24_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_24_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_24_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_24_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_24_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_24_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_24_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_24_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_24_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_24_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_24_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_24_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_24_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_24_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_25_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_25_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_25_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_25_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_25_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_25_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_25_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_25_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_25_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_25_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_25_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_25_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_25_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_25_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_25_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_25_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_25_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_25_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_25_ccff_tail;
wire [0:0] grid_clb_25_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_25_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_25_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_25_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_25_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_25_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_25_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_25_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_25_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_25_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_25_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_25_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_25_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_25_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_25_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_25_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_26_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_26_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_26_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_26_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_26_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_26_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_26_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_26_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_26_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_26_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_26_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_26_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_26_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_26_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_26_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_26_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_26_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_26_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_26_ccff_tail;
wire [0:0] grid_clb_26_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_26_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_26_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_26_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_26_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_26_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_26_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_26_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_26_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_26_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_26_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_26_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_26_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_26_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_26_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_26_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_27_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_27_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_27_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_27_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_27_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_27_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_27_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_27_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_27_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_27_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_27_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_27_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_27_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_27_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_27_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_27_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_27_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_27_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_27_ccff_tail;
wire [0:0] grid_clb_27_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_27_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_27_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_27_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_27_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_27_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_27_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_27_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_27_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_27_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_27_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_27_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_27_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_27_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_27_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_27_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_28_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_28_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_28_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_28_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_28_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_28_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_28_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_28_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_28_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_28_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_28_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_28_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_28_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_28_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_28_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_28_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_28_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_28_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_28_ccff_tail;
wire [0:0] grid_clb_28_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_28_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_28_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_28_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_28_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_28_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_28_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_28_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_28_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_28_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_28_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_28_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_28_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_28_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_28_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_28_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_29_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_29_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_29_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_29_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_29_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_29_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_29_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_29_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_29_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_29_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_29_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_29_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_29_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_29_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_29_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_29_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_29_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_29_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_29_ccff_tail;
wire [0:0] grid_clb_29_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_29_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_29_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_29_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_29_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_29_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_29_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_29_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_29_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_29_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_29_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_29_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_29_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_29_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_29_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_29_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_2_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_2_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_2_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_2_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_2_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_2_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_2_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_2_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_2_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_2_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_2_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_2_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_2_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_2_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_2_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_2_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_2_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_2_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_2_ccff_tail;
wire [0:0] grid_clb_2_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_2_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_2_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_2_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_2_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_2_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_2_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_2_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_2_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_2_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_2_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_2_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_2_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_2_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_2_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_2_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_30_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_30_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_30_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_30_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_30_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_30_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_30_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_30_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_30_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_30_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_30_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_30_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_30_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_30_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_30_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_30_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_30_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_30_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_30_ccff_tail;
wire [0:0] grid_clb_30_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_30_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_30_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_30_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_30_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_30_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_30_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_30_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_30_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_30_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_30_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_30_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_30_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_30_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_30_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_30_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_31_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_31_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_31_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_31_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_31_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_31_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_31_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_31_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_31_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_31_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_31_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_31_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_31_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_31_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_31_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_31_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_31_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_31_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_31_ccff_tail;
wire [0:0] grid_clb_31_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_31_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_31_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_31_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_31_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_31_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_31_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_31_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_31_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_31_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_31_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_31_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_31_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_31_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_31_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_31_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_32_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_32_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_32_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_32_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_32_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_32_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_32_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_32_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_32_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_32_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_32_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_32_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_32_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_32_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_32_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_32_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_32_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_32_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_32_ccff_tail;
wire [0:0] grid_clb_32_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_32_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_32_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_32_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_32_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_32_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_32_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_32_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_32_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_32_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_32_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_32_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_32_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_32_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_32_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_32_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_33_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_33_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_33_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_33_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_33_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_33_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_33_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_33_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_33_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_33_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_33_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_33_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_33_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_33_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_33_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_33_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_33_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_33_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_33_ccff_tail;
wire [0:0] grid_clb_33_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_33_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_33_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_33_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_33_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_33_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_33_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_33_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_33_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_33_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_33_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_33_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_33_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_33_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_33_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_33_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_34_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_34_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_34_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_34_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_34_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_34_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_34_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_34_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_34_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_34_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_34_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_34_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_34_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_34_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_34_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_34_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_34_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_34_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_34_ccff_tail;
wire [0:0] grid_clb_34_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_34_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_34_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_34_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_34_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_34_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_34_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_34_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_34_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_34_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_34_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_34_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_34_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_34_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_34_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_34_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_35_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_35_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_35_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_35_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_35_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_35_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_35_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_35_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_35_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_35_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_35_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_35_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_35_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_35_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_35_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_35_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_35_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_35_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_35_ccff_tail;
wire [0:0] grid_clb_35_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_35_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_35_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_35_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_35_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_35_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_35_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_35_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_35_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_35_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_35_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_35_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_35_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_35_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_35_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_35_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_36_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_36_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_36_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_36_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_36_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_36_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_36_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_36_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_36_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_36_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_36_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_36_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_36_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_36_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_36_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_36_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_36_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_36_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_36_ccff_tail;
wire [0:0] grid_clb_36_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_36_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_36_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_36_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_36_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_36_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_36_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_36_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_36_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_36_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_36_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_36_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_36_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_36_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_36_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_36_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_37_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_37_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_37_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_37_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_37_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_37_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_37_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_37_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_37_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_37_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_37_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_37_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_37_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_37_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_37_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_37_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_37_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_37_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_37_ccff_tail;
wire [0:0] grid_clb_37_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_37_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_37_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_37_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_37_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_37_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_37_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_37_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_37_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_37_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_37_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_37_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_37_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_37_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_37_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_37_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_38_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_38_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_38_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_38_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_38_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_38_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_38_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_38_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_38_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_38_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_38_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_38_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_38_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_38_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_38_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_38_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_38_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_38_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_38_ccff_tail;
wire [0:0] grid_clb_38_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_38_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_38_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_38_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_38_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_38_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_38_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_38_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_38_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_38_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_38_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_38_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_38_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_38_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_38_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_38_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_39_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_39_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_39_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_39_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_39_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_39_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_39_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_39_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_39_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_39_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_39_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_39_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_39_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_39_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_39_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_39_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_39_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_39_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_39_ccff_tail;
wire [0:0] grid_clb_39_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_39_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_39_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_39_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_39_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_39_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_39_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_39_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_39_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_39_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_39_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_39_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_39_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_39_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_39_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_39_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_3_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_3_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_3_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_3_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_3_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_3_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_3_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_3_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_3_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_3_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_3_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_3_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_3_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_3_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_3_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_3_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_3_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_3_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_3_ccff_tail;
wire [0:0] grid_clb_3_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_3_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_3_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_3_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_3_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_3_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_3_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_3_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_3_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_3_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_3_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_3_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_3_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_3_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_3_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_3_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_40_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_40_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_40_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_40_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_40_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_40_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_40_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_40_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_40_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_40_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_40_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_40_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_40_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_40_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_40_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_40_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_40_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_40_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_40_ccff_tail;
wire [0:0] grid_clb_40_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_40_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_40_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_40_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_40_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_40_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_40_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_40_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_40_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_40_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_40_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_40_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_40_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_40_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_40_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_40_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_41_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_41_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_41_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_41_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_41_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_41_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_41_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_41_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_41_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_41_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_41_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_41_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_41_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_41_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_41_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_41_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_41_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_41_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_41_ccff_tail;
wire [0:0] grid_clb_41_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_41_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_41_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_41_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_41_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_41_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_41_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_41_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_41_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_41_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_41_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_41_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_41_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_41_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_41_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_41_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_42_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_42_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_42_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_42_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_42_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_42_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_42_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_42_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_42_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_42_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_42_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_42_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_42_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_42_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_42_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_42_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_42_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_42_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_42_ccff_tail;
wire [0:0] grid_clb_42_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_42_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_42_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_42_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_42_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_42_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_42_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_42_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_42_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_42_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_42_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_42_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_42_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_42_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_42_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_42_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_43_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_43_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_43_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_43_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_43_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_43_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_43_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_43_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_43_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_43_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_43_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_43_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_43_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_43_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_43_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_43_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_43_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_43_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_43_ccff_tail;
wire [0:0] grid_clb_43_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_43_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_43_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_43_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_43_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_43_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_43_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_43_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_43_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_43_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_43_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_43_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_43_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_43_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_43_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_43_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_44_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_44_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_44_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_44_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_44_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_44_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_44_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_44_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_44_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_44_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_44_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_44_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_44_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_44_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_44_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_44_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_44_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_44_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_44_ccff_tail;
wire [0:0] grid_clb_44_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_44_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_44_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_44_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_44_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_44_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_44_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_44_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_44_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_44_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_44_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_44_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_44_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_44_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_44_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_44_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_45_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_45_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_45_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_45_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_45_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_45_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_45_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_45_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_45_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_45_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_45_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_45_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_45_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_45_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_45_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_45_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_45_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_45_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_45_ccff_tail;
wire [0:0] grid_clb_45_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_45_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_45_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_45_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_45_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_45_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_45_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_45_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_45_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_45_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_45_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_45_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_45_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_45_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_45_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_45_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_46_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_46_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_46_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_46_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_46_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_46_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_46_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_46_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_46_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_46_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_46_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_46_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_46_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_46_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_46_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_46_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_46_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_46_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_46_ccff_tail;
wire [0:0] grid_clb_46_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_46_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_46_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_46_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_46_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_46_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_46_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_46_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_46_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_46_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_46_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_46_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_46_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_46_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_46_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_46_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_47_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_47_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_47_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_47_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_47_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_47_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_47_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_47_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_47_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_47_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_47_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_47_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_47_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_47_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_47_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_47_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_47_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_47_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_47_ccff_tail;
wire [0:0] grid_clb_47_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_47_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_47_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_47_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_47_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_47_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_47_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_47_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_47_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_47_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_47_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_47_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_47_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_47_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_47_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_47_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_48_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_48_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_48_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_48_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_48_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_48_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_48_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_48_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_48_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_48_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_48_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_48_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_48_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_48_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_48_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_48_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_48_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_48_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_48_ccff_tail;
wire [0:0] grid_clb_48_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_48_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_48_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_48_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_48_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_48_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_48_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_48_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_48_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_48_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_48_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_48_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_48_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_48_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_48_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_48_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_49_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_49_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_49_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_49_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_49_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_49_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_49_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_49_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_49_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_49_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_49_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_49_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_49_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_49_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_49_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_49_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_49_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_49_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_49_ccff_tail;
wire [0:0] grid_clb_49_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_49_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_49_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_49_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_49_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_49_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_49_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_49_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_49_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_49_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_49_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_49_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_49_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_49_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_49_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_49_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_4_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_4_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_4_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_4_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_4_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_4_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_4_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_4_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_4_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_4_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_4_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_4_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_4_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_4_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_4_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_4_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_4_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_4_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_4_ccff_tail;
wire [0:0] grid_clb_4_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_4_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_4_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_4_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_4_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_4_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_4_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_4_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_4_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_4_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_4_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_4_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_4_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_4_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_4_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_4_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_50_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_50_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_50_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_50_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_50_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_50_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_50_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_50_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_50_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_50_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_50_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_50_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_50_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_50_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_50_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_50_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_50_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_50_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_50_ccff_tail;
wire [0:0] grid_clb_50_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_50_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_50_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_50_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_50_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_50_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_50_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_50_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_50_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_50_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_50_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_50_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_50_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_50_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_50_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_50_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_51_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_51_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_51_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_51_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_51_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_51_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_51_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_51_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_51_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_51_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_51_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_51_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_51_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_51_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_51_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_51_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_51_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_51_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_51_ccff_tail;
wire [0:0] grid_clb_51_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_51_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_51_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_51_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_51_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_51_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_51_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_51_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_51_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_51_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_51_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_51_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_51_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_51_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_51_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_51_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_52_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_52_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_52_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_52_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_52_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_52_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_52_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_52_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_52_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_52_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_52_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_52_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_52_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_52_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_52_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_52_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_52_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_52_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_52_ccff_tail;
wire [0:0] grid_clb_52_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_52_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_52_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_52_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_52_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_52_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_52_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_52_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_52_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_52_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_52_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_52_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_52_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_52_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_52_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_52_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_53_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_53_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_53_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_53_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_53_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_53_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_53_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_53_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_53_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_53_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_53_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_53_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_53_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_53_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_53_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_53_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_53_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_53_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_53_ccff_tail;
wire [0:0] grid_clb_53_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_53_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_53_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_53_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_53_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_53_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_53_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_53_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_53_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_53_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_53_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_53_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_53_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_53_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_53_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_53_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_54_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_54_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_54_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_54_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_54_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_54_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_54_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_54_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_54_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_54_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_54_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_54_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_54_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_54_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_54_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_54_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_54_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_54_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_54_ccff_tail;
wire [0:0] grid_clb_54_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_54_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_54_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_54_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_54_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_54_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_54_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_54_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_54_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_54_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_54_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_54_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_54_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_54_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_54_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_54_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_55_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_55_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_55_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_55_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_55_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_55_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_55_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_55_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_55_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_55_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_55_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_55_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_55_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_55_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_55_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_55_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_55_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_55_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_55_ccff_tail;
wire [0:0] grid_clb_55_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_55_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_55_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_55_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_55_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_55_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_55_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_55_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_55_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_55_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_55_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_55_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_55_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_55_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_55_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_55_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_56_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_56_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_56_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_56_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_56_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_56_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_56_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_56_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_56_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_56_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_56_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_56_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_56_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_56_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_56_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_56_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_56_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_56_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_56_ccff_tail;
wire [0:0] grid_clb_56_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_56_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_56_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_56_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_56_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_56_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_56_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_56_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_56_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_56_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_56_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_56_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_56_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_56_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_56_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_56_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_57_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_57_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_57_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_57_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_57_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_57_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_57_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_57_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_57_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_57_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_57_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_57_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_57_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_57_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_57_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_57_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_57_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_57_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_57_ccff_tail;
wire [0:0] grid_clb_57_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_57_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_57_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_57_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_57_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_57_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_57_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_57_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_57_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_57_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_57_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_57_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_57_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_57_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_57_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_57_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_58_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_58_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_58_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_58_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_58_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_58_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_58_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_58_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_58_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_58_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_58_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_58_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_58_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_58_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_58_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_58_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_58_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_58_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_58_ccff_tail;
wire [0:0] grid_clb_58_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_58_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_58_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_58_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_58_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_58_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_58_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_58_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_58_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_58_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_58_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_58_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_58_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_58_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_58_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_58_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_59_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_59_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_59_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_59_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_59_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_59_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_59_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_59_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_59_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_59_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_59_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_59_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_59_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_59_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_59_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_59_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_59_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_59_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_59_ccff_tail;
wire [0:0] grid_clb_59_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_59_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_59_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_59_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_59_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_59_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_59_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_59_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_59_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_59_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_59_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_59_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_59_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_59_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_59_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_59_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_5_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_5_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_5_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_5_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_5_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_5_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_5_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_5_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_5_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_5_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_5_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_5_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_5_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_5_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_5_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_5_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_5_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_5_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_5_ccff_tail;
wire [0:0] grid_clb_5_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_5_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_5_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_5_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_5_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_5_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_5_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_5_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_5_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_5_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_5_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_5_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_5_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_5_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_5_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_5_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_60_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_60_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_60_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_60_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_60_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_60_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_60_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_60_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_60_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_60_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_60_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_60_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_60_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_60_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_60_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_60_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_60_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_60_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_60_ccff_tail;
wire [0:0] grid_clb_60_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_60_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_60_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_60_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_60_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_60_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_60_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_60_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_60_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_60_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_60_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_60_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_60_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_60_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_60_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_60_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_61_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_61_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_61_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_61_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_61_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_61_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_61_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_61_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_61_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_61_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_61_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_61_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_61_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_61_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_61_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_61_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_61_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_61_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_61_ccff_tail;
wire [0:0] grid_clb_61_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_61_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_61_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_61_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_61_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_61_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_61_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_61_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_61_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_61_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_61_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_61_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_61_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_61_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_61_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_61_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_62_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_62_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_62_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_62_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_62_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_62_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_62_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_62_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_62_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_62_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_62_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_62_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_62_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_62_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_62_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_62_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_62_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_62_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_62_ccff_tail;
wire [0:0] grid_clb_62_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_62_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_62_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_62_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_62_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_62_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_62_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_62_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_62_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_62_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_62_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_62_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_62_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_62_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_62_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_62_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_63_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_63_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_63_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_63_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_63_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_63_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_63_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_63_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_63_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_63_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_63_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_63_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_63_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_63_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_63_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_63_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_63_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_63_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_63_ccff_tail;
wire [0:0] grid_clb_63_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_63_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_63_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_63_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_63_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_63_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_63_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_63_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_63_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_63_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_63_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_63_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_63_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_63_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_63_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_63_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_64_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_64_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_64_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_64_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_64_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_64_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_64_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_64_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_64_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_64_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_64_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_64_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_64_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_64_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_64_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_64_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_64_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_64_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_64_ccff_tail;
wire [0:0] grid_clb_64_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_64_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_64_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_64_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_64_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_64_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_64_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_64_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_64_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_64_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_64_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_64_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_64_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_64_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_64_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_64_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_65_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_65_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_65_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_65_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_65_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_65_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_65_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_65_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_65_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_65_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_65_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_65_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_65_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_65_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_65_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_65_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_65_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_65_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_65_ccff_tail;
wire [0:0] grid_clb_65_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_65_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_65_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_65_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_65_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_65_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_65_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_65_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_65_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_65_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_65_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_65_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_65_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_65_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_65_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_65_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_66_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_66_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_66_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_66_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_66_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_66_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_66_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_66_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_66_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_66_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_66_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_66_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_66_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_66_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_66_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_66_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_66_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_66_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_66_ccff_tail;
wire [0:0] grid_clb_66_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_66_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_66_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_66_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_66_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_66_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_66_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_66_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_66_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_66_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_66_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_66_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_66_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_66_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_66_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_66_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_67_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_67_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_67_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_67_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_67_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_67_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_67_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_67_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_67_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_67_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_67_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_67_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_67_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_67_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_67_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_67_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_67_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_67_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_67_ccff_tail;
wire [0:0] grid_clb_67_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_67_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_67_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_67_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_67_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_67_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_67_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_67_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_67_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_67_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_67_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_67_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_67_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_67_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_67_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_67_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_68_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_68_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_68_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_68_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_68_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_68_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_68_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_68_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_68_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_68_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_68_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_68_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_68_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_68_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_68_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_68_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_68_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_68_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_68_ccff_tail;
wire [0:0] grid_clb_68_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_68_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_68_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_68_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_68_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_68_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_68_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_68_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_68_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_68_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_68_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_68_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_68_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_68_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_68_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_68_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_69_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_69_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_69_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_69_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_69_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_69_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_69_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_69_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_69_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_69_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_69_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_69_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_69_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_69_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_69_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_69_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_69_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_69_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_69_ccff_tail;
wire [0:0] grid_clb_69_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_69_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_69_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_69_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_69_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_69_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_69_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_69_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_69_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_69_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_69_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_69_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_69_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_69_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_69_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_69_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_6_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_6_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_6_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_6_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_6_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_6_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_6_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_6_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_6_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_6_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_6_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_6_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_6_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_6_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_6_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_6_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_6_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_6_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_6_ccff_tail;
wire [0:0] grid_clb_6_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_6_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_6_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_6_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_6_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_6_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_6_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_6_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_6_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_6_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_6_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_6_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_6_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_6_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_6_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_6_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_70_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_70_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_70_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_70_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_70_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_70_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_70_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_70_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_70_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_70_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_70_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_70_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_70_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_70_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_70_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_70_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_70_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_70_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_70_ccff_tail;
wire [0:0] grid_clb_70_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_70_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_70_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_70_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_70_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_70_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_70_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_70_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_70_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_70_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_70_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_70_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_70_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_70_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_70_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_70_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_71_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_71_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_71_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_71_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_71_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_71_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_71_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_71_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_71_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_71_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_71_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_71_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_71_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_71_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_71_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_71_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_71_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_71_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_71_ccff_tail;
wire [0:0] grid_clb_71_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_71_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_71_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_71_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_71_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_71_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_71_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_71_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_71_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_71_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_71_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_71_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_71_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_71_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_71_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_71_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_72_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_72_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_72_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_72_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_72_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_72_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_72_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_72_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_72_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_72_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_72_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_72_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_72_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_72_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_72_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_72_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_72_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_72_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_72_ccff_tail;
wire [0:0] grid_clb_72_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_72_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_72_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_72_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_72_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_72_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_72_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_72_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_72_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_72_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_72_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_72_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_72_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_72_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_72_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_72_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_73_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_73_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_73_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_73_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_73_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_73_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_73_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_73_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_73_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_73_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_73_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_73_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_73_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_73_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_73_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_73_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_73_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_73_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_73_ccff_tail;
wire [0:0] grid_clb_73_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_73_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_73_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_73_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_73_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_73_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_73_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_73_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_73_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_73_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_73_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_73_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_73_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_73_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_73_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_73_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_74_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_74_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_74_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_74_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_74_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_74_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_74_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_74_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_74_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_74_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_74_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_74_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_74_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_74_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_74_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_74_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_74_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_74_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_74_ccff_tail;
wire [0:0] grid_clb_74_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_74_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_74_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_74_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_74_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_74_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_74_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_74_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_74_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_74_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_74_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_74_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_74_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_74_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_74_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_74_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_75_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_75_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_75_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_75_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_75_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_75_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_75_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_75_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_75_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_75_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_75_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_75_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_75_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_75_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_75_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_75_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_75_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_75_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_75_ccff_tail;
wire [0:0] grid_clb_75_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_75_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_75_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_75_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_75_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_75_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_75_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_75_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_75_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_75_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_75_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_75_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_75_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_75_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_75_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_75_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_76_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_76_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_76_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_76_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_76_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_76_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_76_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_76_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_76_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_76_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_76_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_76_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_76_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_76_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_76_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_76_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_76_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_76_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_76_ccff_tail;
wire [0:0] grid_clb_76_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_76_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_76_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_76_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_76_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_76_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_76_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_76_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_76_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_76_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_76_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_76_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_76_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_76_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_76_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_76_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_77_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_77_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_77_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_77_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_77_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_77_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_77_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_77_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_77_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_77_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_77_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_77_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_77_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_77_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_77_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_77_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_77_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_77_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_77_ccff_tail;
wire [0:0] grid_clb_77_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_77_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_77_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_77_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_77_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_77_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_77_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_77_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_77_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_77_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_77_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_77_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_77_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_77_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_77_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_77_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_78_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_78_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_78_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_78_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_78_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_78_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_78_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_78_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_78_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_78_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_78_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_78_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_78_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_78_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_78_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_78_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_78_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_78_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_78_ccff_tail;
wire [0:0] grid_clb_78_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_78_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_78_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_78_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_78_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_78_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_78_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_78_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_78_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_78_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_78_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_78_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_78_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_78_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_78_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_78_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_79_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_79_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_79_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_79_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_79_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_79_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_79_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_79_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_79_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_79_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_79_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_79_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_79_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_79_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_79_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_79_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_79_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_79_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_79_ccff_tail;
wire [0:0] grid_clb_79_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_79_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_79_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_79_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_79_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_79_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_79_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_79_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_79_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_79_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_79_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_79_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_79_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_79_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_79_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_79_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_7_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_7_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_7_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_7_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_7_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_7_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_7_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_7_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_7_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_7_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_7_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_7_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_7_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_7_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_7_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_7_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_7_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_7_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_7_ccff_tail;
wire [0:0] grid_clb_7_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_7_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_7_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_7_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_7_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_7_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_7_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_7_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_7_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_7_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_7_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_7_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_7_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_7_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_7_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_7_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_80_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_80_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_80_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_80_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_80_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_80_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_80_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_80_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_80_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_80_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_80_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_80_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_80_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_80_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_80_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_80_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_80_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_80_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_80_ccff_tail;
wire [0:0] grid_clb_80_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_80_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_80_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_80_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_80_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_80_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_80_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_80_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_80_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_80_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_80_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_80_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_80_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_80_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_80_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_80_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_81_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_81_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_81_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_81_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_81_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_81_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_81_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_81_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_81_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_81_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_81_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_81_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_81_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_81_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_81_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_81_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_81_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_81_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_81_ccff_tail;
wire [0:0] grid_clb_81_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_81_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_81_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_81_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_81_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_81_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_81_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_81_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_81_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_81_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_81_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_81_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_81_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_81_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_81_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_81_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_82_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_82_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_82_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_82_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_82_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_82_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_82_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_82_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_82_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_82_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_82_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_82_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_82_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_82_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_82_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_82_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_82_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_82_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_82_ccff_tail;
wire [0:0] grid_clb_82_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_82_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_82_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_82_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_82_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_82_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_82_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_82_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_82_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_82_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_82_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_82_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_82_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_82_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_82_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_82_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_83_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_83_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_83_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_83_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_83_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_83_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_83_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_83_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_83_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_83_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_83_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_83_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_83_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_83_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_83_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_83_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_83_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_83_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_83_ccff_tail;
wire [0:0] grid_clb_83_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_83_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_83_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_83_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_83_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_83_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_83_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_83_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_83_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_83_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_83_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_83_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_83_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_83_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_83_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_83_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_84_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_84_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_84_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_84_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_84_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_84_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_84_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_84_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_84_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_84_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_84_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_84_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_84_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_84_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_84_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_84_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_84_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_84_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_84_ccff_tail;
wire [0:0] grid_clb_84_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_84_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_84_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_84_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_84_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_84_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_84_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_84_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_84_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_84_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_84_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_84_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_84_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_84_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_84_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_84_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_85_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_85_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_85_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_85_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_85_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_85_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_85_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_85_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_85_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_85_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_85_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_85_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_85_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_85_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_85_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_85_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_85_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_85_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_85_ccff_tail;
wire [0:0] grid_clb_85_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_85_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_85_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_85_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_85_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_85_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_85_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_85_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_85_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_85_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_85_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_85_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_85_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_85_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_85_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_85_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_86_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_86_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_86_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_86_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_86_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_86_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_86_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_86_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_86_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_86_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_86_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_86_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_86_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_86_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_86_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_86_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_86_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_86_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_86_ccff_tail;
wire [0:0] grid_clb_86_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_86_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_86_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_86_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_86_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_86_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_86_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_86_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_86_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_86_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_86_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_86_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_86_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_86_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_86_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_86_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_87_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_87_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_87_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_87_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_87_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_87_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_87_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_87_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_87_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_87_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_87_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_87_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_87_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_87_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_87_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_87_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_87_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_87_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_87_ccff_tail;
wire [0:0] grid_clb_87_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_87_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_87_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_87_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_87_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_87_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_87_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_87_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_87_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_87_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_87_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_87_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_87_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_87_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_87_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_87_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_88_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_88_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_88_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_88_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_88_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_88_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_88_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_88_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_88_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_88_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_88_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_88_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_88_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_88_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_88_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_88_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_88_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_88_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_88_ccff_tail;
wire [0:0] grid_clb_88_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_88_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_88_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_88_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_88_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_88_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_88_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_88_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_88_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_88_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_88_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_88_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_88_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_88_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_88_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_88_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_89_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_89_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_89_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_89_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_89_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_89_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_89_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_89_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_89_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_89_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_89_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_89_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_89_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_89_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_89_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_89_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_89_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_89_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_89_ccff_tail;
wire [0:0] grid_clb_89_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_89_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_89_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_89_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_89_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_89_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_89_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_89_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_89_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_89_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_89_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_89_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_89_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_89_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_89_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_89_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_8_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_8_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_8_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_8_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_8_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_8_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_8_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_8_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_8_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_8_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_8_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_8_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_8_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_8_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_8_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_8_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_8_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_8_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_8_ccff_tail;
wire [0:0] grid_clb_8_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_8_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_8_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_8_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_8_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_8_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_8_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_8_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_8_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_8_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_8_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_8_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_8_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_8_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_8_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_8_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_90_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_90_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_90_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_90_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_90_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_90_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_90_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_90_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_90_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_90_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_90_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_90_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_90_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_90_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_90_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_90_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_90_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_90_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_90_ccff_tail;
wire [0:0] grid_clb_90_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_90_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_90_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_90_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_90_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_90_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_90_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_90_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_90_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_90_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_90_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_90_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_90_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_90_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_90_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_90_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_91_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_91_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_91_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_91_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_91_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_91_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_91_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_91_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_91_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_91_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_91_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_91_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_91_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_91_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_91_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_91_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_91_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_91_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_91_ccff_tail;
wire [0:0] grid_clb_91_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_91_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_91_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_91_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_91_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_91_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_91_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_91_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_91_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_91_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_91_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_91_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_91_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_91_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_91_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_91_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_92_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_92_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_92_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_92_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_92_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_92_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_92_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_92_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_92_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_92_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_92_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_92_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_92_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_92_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_92_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_92_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_92_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_92_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_92_ccff_tail;
wire [0:0] grid_clb_92_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_92_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_92_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_92_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_92_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_92_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_92_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_92_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_92_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_92_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_92_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_92_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_92_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_92_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_92_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_92_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_93_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_93_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_93_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_93_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_93_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_93_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_93_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_93_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_93_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_93_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_93_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_93_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_93_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_93_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_93_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_93_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_93_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_93_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_93_ccff_tail;
wire [0:0] grid_clb_93_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_93_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_93_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_93_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_93_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_93_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_93_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_93_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_93_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_93_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_93_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_93_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_93_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_93_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_93_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_93_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_94_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_94_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_94_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_94_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_94_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_94_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_94_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_94_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_94_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_94_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_94_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_94_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_94_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_94_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_94_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_94_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_94_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_94_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_94_ccff_tail;
wire [0:0] grid_clb_94_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_94_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_94_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_94_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_94_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_94_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_94_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_94_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_94_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_94_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_94_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_94_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_94_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_94_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_94_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_94_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_95_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_95_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_95_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_95_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_95_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_95_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_95_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_95_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_95_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_95_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_95_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_95_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_95_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_95_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_95_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_95_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_95_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_95_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_95_ccff_tail;
wire [0:0] grid_clb_95_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_95_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_95_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_95_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_95_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_95_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_95_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_95_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_95_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_95_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_95_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_95_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_95_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_95_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_95_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_95_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_96_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_96_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_96_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_96_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_96_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_96_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_96_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_96_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_96_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_96_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_96_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_96_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_96_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_96_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_96_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_96_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_96_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_96_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_96_ccff_tail;
wire [0:0] grid_clb_96_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_96_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_96_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_96_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_96_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_96_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_96_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_96_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_96_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_96_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_96_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_96_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_96_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_96_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_96_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_96_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_97_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_97_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_97_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_97_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_97_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_97_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_97_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_97_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_97_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_97_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_97_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_97_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_97_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_97_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_97_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_97_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_97_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_97_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_97_ccff_tail;
wire [0:0] grid_clb_97_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_97_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_97_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_97_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_97_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_97_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_97_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_97_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_97_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_97_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_97_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_97_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_97_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_97_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_97_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_97_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_98_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_98_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_98_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_98_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_98_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_98_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_98_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_98_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_98_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_98_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_98_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_98_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_98_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_98_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_98_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_98_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_98_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_98_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_98_ccff_tail;
wire [0:0] grid_clb_98_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_98_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_98_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_98_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_98_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_98_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_98_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_98_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_98_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_98_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_98_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_98_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_98_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_98_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_98_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_98_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_99_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_99_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_99_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_99_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_99_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_99_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_99_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_99_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_99_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_99_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_99_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_99_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_99_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_99_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_99_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_99_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_99_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_99_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_99_ccff_tail;
wire [0:0] grid_clb_99_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_99_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_99_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_99_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_99_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_99_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_99_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_99_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_99_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_99_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_99_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_99_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_99_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_99_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_99_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_99_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_clb_9_bottom_width_0_height_0__pin_42_lower;
wire [0:0] grid_clb_9_bottom_width_0_height_0__pin_42_upper;
wire [0:0] grid_clb_9_bottom_width_0_height_0__pin_43_lower;
wire [0:0] grid_clb_9_bottom_width_0_height_0__pin_43_upper;
wire [0:0] grid_clb_9_bottom_width_0_height_0__pin_44_lower;
wire [0:0] grid_clb_9_bottom_width_0_height_0__pin_44_upper;
wire [0:0] grid_clb_9_bottom_width_0_height_0__pin_45_lower;
wire [0:0] grid_clb_9_bottom_width_0_height_0__pin_45_upper;
wire [0:0] grid_clb_9_bottom_width_0_height_0__pin_46_lower;
wire [0:0] grid_clb_9_bottom_width_0_height_0__pin_46_upper;
wire [0:0] grid_clb_9_bottom_width_0_height_0__pin_47_lower;
wire [0:0] grid_clb_9_bottom_width_0_height_0__pin_47_upper;
wire [0:0] grid_clb_9_bottom_width_0_height_0__pin_48_lower;
wire [0:0] grid_clb_9_bottom_width_0_height_0__pin_48_upper;
wire [0:0] grid_clb_9_bottom_width_0_height_0__pin_49_lower;
wire [0:0] grid_clb_9_bottom_width_0_height_0__pin_49_upper;
wire [0:0] grid_clb_9_bottom_width_0_height_0__pin_50_;
wire [0:0] grid_clb_9_bottom_width_0_height_0__pin_51_;
wire [0:0] grid_clb_9_ccff_tail;
wire [0:0] grid_clb_9_right_width_0_height_0__pin_34_lower;
wire [0:0] grid_clb_9_right_width_0_height_0__pin_34_upper;
wire [0:0] grid_clb_9_right_width_0_height_0__pin_35_lower;
wire [0:0] grid_clb_9_right_width_0_height_0__pin_35_upper;
wire [0:0] grid_clb_9_right_width_0_height_0__pin_36_lower;
wire [0:0] grid_clb_9_right_width_0_height_0__pin_36_upper;
wire [0:0] grid_clb_9_right_width_0_height_0__pin_37_lower;
wire [0:0] grid_clb_9_right_width_0_height_0__pin_37_upper;
wire [0:0] grid_clb_9_right_width_0_height_0__pin_38_lower;
wire [0:0] grid_clb_9_right_width_0_height_0__pin_38_upper;
wire [0:0] grid_clb_9_right_width_0_height_0__pin_39_lower;
wire [0:0] grid_clb_9_right_width_0_height_0__pin_39_upper;
wire [0:0] grid_clb_9_right_width_0_height_0__pin_40_lower;
wire [0:0] grid_clb_9_right_width_0_height_0__pin_40_upper;
wire [0:0] grid_clb_9_right_width_0_height_0__pin_41_lower;
wire [0:0] grid_clb_9_right_width_0_height_0__pin_41_upper;
wire [0:0] grid_io_bottom_0_ccff_tail;
wire [0:0] grid_io_bottom_0_top_width_0_height_0__pin_1_lower;
wire [0:0] grid_io_bottom_0_top_width_0_height_0__pin_1_upper;
wire [0:0] grid_io_bottom_10_ccff_tail;
wire [0:0] grid_io_bottom_10_top_width_0_height_0__pin_1_lower;
wire [0:0] grid_io_bottom_10_top_width_0_height_0__pin_1_upper;
wire [0:0] grid_io_bottom_11_ccff_tail;
wire [0:0] grid_io_bottom_11_top_width_0_height_0__pin_1_lower;
wire [0:0] grid_io_bottom_11_top_width_0_height_0__pin_1_upper;
wire [0:0] grid_io_bottom_1_ccff_tail;
wire [0:0] grid_io_bottom_1_top_width_0_height_0__pin_1_lower;
wire [0:0] grid_io_bottom_1_top_width_0_height_0__pin_1_upper;
wire [0:0] grid_io_bottom_2_ccff_tail;
wire [0:0] grid_io_bottom_2_top_width_0_height_0__pin_1_lower;
wire [0:0] grid_io_bottom_2_top_width_0_height_0__pin_1_upper;
wire [0:0] grid_io_bottom_3_ccff_tail;
wire [0:0] grid_io_bottom_3_top_width_0_height_0__pin_1_lower;
wire [0:0] grid_io_bottom_3_top_width_0_height_0__pin_1_upper;
wire [0:0] grid_io_bottom_4_ccff_tail;
wire [0:0] grid_io_bottom_4_top_width_0_height_0__pin_1_lower;
wire [0:0] grid_io_bottom_4_top_width_0_height_0__pin_1_upper;
wire [0:0] grid_io_bottom_5_ccff_tail;
wire [0:0] grid_io_bottom_5_top_width_0_height_0__pin_1_lower;
wire [0:0] grid_io_bottom_5_top_width_0_height_0__pin_1_upper;
wire [0:0] grid_io_bottom_6_ccff_tail;
wire [0:0] grid_io_bottom_6_top_width_0_height_0__pin_1_lower;
wire [0:0] grid_io_bottom_6_top_width_0_height_0__pin_1_upper;
wire [0:0] grid_io_bottom_7_ccff_tail;
wire [0:0] grid_io_bottom_7_top_width_0_height_0__pin_1_lower;
wire [0:0] grid_io_bottom_7_top_width_0_height_0__pin_1_upper;
wire [0:0] grid_io_bottom_8_ccff_tail;
wire [0:0] grid_io_bottom_8_top_width_0_height_0__pin_1_lower;
wire [0:0] grid_io_bottom_8_top_width_0_height_0__pin_1_upper;
wire [0:0] grid_io_bottom_9_ccff_tail;
wire [0:0] grid_io_bottom_9_top_width_0_height_0__pin_1_lower;
wire [0:0] grid_io_bottom_9_top_width_0_height_0__pin_1_upper;
wire [0:0] grid_io_left_0_ccff_tail;
wire [0:0] grid_io_left_0_right_width_0_height_0__pin_1_lower;
wire [0:0] grid_io_left_0_right_width_0_height_0__pin_1_upper;
wire [0:0] grid_io_left_10_ccff_tail;
wire [0:0] grid_io_left_10_right_width_0_height_0__pin_1_lower;
wire [0:0] grid_io_left_10_right_width_0_height_0__pin_1_upper;
wire [0:0] grid_io_left_11_ccff_tail;
wire [0:0] grid_io_left_11_right_width_0_height_0__pin_1_lower;
wire [0:0] grid_io_left_11_right_width_0_height_0__pin_1_upper;
wire [0:0] grid_io_left_1_ccff_tail;
wire [0:0] grid_io_left_1_right_width_0_height_0__pin_1_lower;
wire [0:0] grid_io_left_1_right_width_0_height_0__pin_1_upper;
wire [0:0] grid_io_left_2_ccff_tail;
wire [0:0] grid_io_left_2_right_width_0_height_0__pin_1_lower;
wire [0:0] grid_io_left_2_right_width_0_height_0__pin_1_upper;
wire [0:0] grid_io_left_3_ccff_tail;
wire [0:0] grid_io_left_3_right_width_0_height_0__pin_1_lower;
wire [0:0] grid_io_left_3_right_width_0_height_0__pin_1_upper;
wire [0:0] grid_io_left_4_ccff_tail;
wire [0:0] grid_io_left_4_right_width_0_height_0__pin_1_lower;
wire [0:0] grid_io_left_4_right_width_0_height_0__pin_1_upper;
wire [0:0] grid_io_left_5_ccff_tail;
wire [0:0] grid_io_left_5_right_width_0_height_0__pin_1_lower;
wire [0:0] grid_io_left_5_right_width_0_height_0__pin_1_upper;
wire [0:0] grid_io_left_6_ccff_tail;
wire [0:0] grid_io_left_6_right_width_0_height_0__pin_1_lower;
wire [0:0] grid_io_left_6_right_width_0_height_0__pin_1_upper;
wire [0:0] grid_io_left_7_ccff_tail;
wire [0:0] grid_io_left_7_right_width_0_height_0__pin_1_lower;
wire [0:0] grid_io_left_7_right_width_0_height_0__pin_1_upper;
wire [0:0] grid_io_left_8_ccff_tail;
wire [0:0] grid_io_left_8_right_width_0_height_0__pin_1_lower;
wire [0:0] grid_io_left_8_right_width_0_height_0__pin_1_upper;
wire [0:0] grid_io_left_9_ccff_tail;
wire [0:0] grid_io_left_9_right_width_0_height_0__pin_1_lower;
wire [0:0] grid_io_left_9_right_width_0_height_0__pin_1_upper;
wire [0:0] grid_io_right_0_ccff_tail;
wire [0:0] grid_io_right_0_left_width_0_height_0__pin_1_lower;
wire [0:0] grid_io_right_0_left_width_0_height_0__pin_1_upper;
wire [0:0] grid_io_right_10_ccff_tail;
wire [0:0] grid_io_right_10_left_width_0_height_0__pin_1_lower;
wire [0:0] grid_io_right_10_left_width_0_height_0__pin_1_upper;
wire [0:0] grid_io_right_11_ccff_tail;
wire [0:0] grid_io_right_11_left_width_0_height_0__pin_1_lower;
wire [0:0] grid_io_right_11_left_width_0_height_0__pin_1_upper;
wire [0:0] grid_io_right_1_ccff_tail;
wire [0:0] grid_io_right_1_left_width_0_height_0__pin_1_lower;
wire [0:0] grid_io_right_1_left_width_0_height_0__pin_1_upper;
wire [0:0] grid_io_right_2_ccff_tail;
wire [0:0] grid_io_right_2_left_width_0_height_0__pin_1_lower;
wire [0:0] grid_io_right_2_left_width_0_height_0__pin_1_upper;
wire [0:0] grid_io_right_3_ccff_tail;
wire [0:0] grid_io_right_3_left_width_0_height_0__pin_1_lower;
wire [0:0] grid_io_right_3_left_width_0_height_0__pin_1_upper;
wire [0:0] grid_io_right_4_ccff_tail;
wire [0:0] grid_io_right_4_left_width_0_height_0__pin_1_lower;
wire [0:0] grid_io_right_4_left_width_0_height_0__pin_1_upper;
wire [0:0] grid_io_right_5_ccff_tail;
wire [0:0] grid_io_right_5_left_width_0_height_0__pin_1_lower;
wire [0:0] grid_io_right_5_left_width_0_height_0__pin_1_upper;
wire [0:0] grid_io_right_6_ccff_tail;
wire [0:0] grid_io_right_6_left_width_0_height_0__pin_1_lower;
wire [0:0] grid_io_right_6_left_width_0_height_0__pin_1_upper;
wire [0:0] grid_io_right_7_ccff_tail;
wire [0:0] grid_io_right_7_left_width_0_height_0__pin_1_lower;
wire [0:0] grid_io_right_7_left_width_0_height_0__pin_1_upper;
wire [0:0] grid_io_right_8_ccff_tail;
wire [0:0] grid_io_right_8_left_width_0_height_0__pin_1_lower;
wire [0:0] grid_io_right_8_left_width_0_height_0__pin_1_upper;
wire [0:0] grid_io_right_9_ccff_tail;
wire [0:0] grid_io_right_9_left_width_0_height_0__pin_1_lower;
wire [0:0] grid_io_right_9_left_width_0_height_0__pin_1_upper;
wire [0:0] grid_io_top_0_bottom_width_0_height_0__pin_1_lower;
wire [0:0] grid_io_top_0_bottom_width_0_height_0__pin_1_upper;
wire [0:0] grid_io_top_0_ccff_tail;
wire [0:0] grid_io_top_10_bottom_width_0_height_0__pin_1_lower;
wire [0:0] grid_io_top_10_bottom_width_0_height_0__pin_1_upper;
wire [0:0] grid_io_top_10_ccff_tail;
wire [0:0] grid_io_top_11_bottom_width_0_height_0__pin_1_lower;
wire [0:0] grid_io_top_11_bottom_width_0_height_0__pin_1_upper;
wire [0:0] grid_io_top_11_ccff_tail;
wire [0:0] grid_io_top_1_bottom_width_0_height_0__pin_1_lower;
wire [0:0] grid_io_top_1_bottom_width_0_height_0__pin_1_upper;
wire [0:0] grid_io_top_1_ccff_tail;
wire [0:0] grid_io_top_2_bottom_width_0_height_0__pin_1_lower;
wire [0:0] grid_io_top_2_bottom_width_0_height_0__pin_1_upper;
wire [0:0] grid_io_top_2_ccff_tail;
wire [0:0] grid_io_top_3_bottom_width_0_height_0__pin_1_lower;
wire [0:0] grid_io_top_3_bottom_width_0_height_0__pin_1_upper;
wire [0:0] grid_io_top_3_ccff_tail;
wire [0:0] grid_io_top_4_bottom_width_0_height_0__pin_1_lower;
wire [0:0] grid_io_top_4_bottom_width_0_height_0__pin_1_upper;
wire [0:0] grid_io_top_4_ccff_tail;
wire [0:0] grid_io_top_5_bottom_width_0_height_0__pin_1_lower;
wire [0:0] grid_io_top_5_bottom_width_0_height_0__pin_1_upper;
wire [0:0] grid_io_top_5_ccff_tail;
wire [0:0] grid_io_top_6_bottom_width_0_height_0__pin_1_lower;
wire [0:0] grid_io_top_6_bottom_width_0_height_0__pin_1_upper;
wire [0:0] grid_io_top_6_ccff_tail;
wire [0:0] grid_io_top_7_bottom_width_0_height_0__pin_1_lower;
wire [0:0] grid_io_top_7_bottom_width_0_height_0__pin_1_upper;
wire [0:0] grid_io_top_7_ccff_tail;
wire [0:0] grid_io_top_8_bottom_width_0_height_0__pin_1_lower;
wire [0:0] grid_io_top_8_bottom_width_0_height_0__pin_1_upper;
wire [0:0] grid_io_top_8_ccff_tail;
wire [0:0] grid_io_top_9_bottom_width_0_height_0__pin_1_lower;
wire [0:0] grid_io_top_9_bottom_width_0_height_0__pin_1_upper;
wire [0:0] grid_io_top_9_ccff_tail;
wire [0:19] sb_0__0__0_chanx_right_out;
wire [0:19] sb_0__0__0_chany_top_out;
wire [0:0] sb_0__12__0_ccff_tail;
wire [0:19] sb_0__12__0_chanx_right_out;
wire [0:19] sb_0__12__0_chany_bottom_out;
wire [0:0] sb_0__1__0_ccff_tail;
wire [0:19] sb_0__1__0_chanx_right_out;
wire [0:19] sb_0__1__0_chany_bottom_out;
wire [0:19] sb_0__1__0_chany_top_out;
wire [0:0] sb_0__1__10_ccff_tail;
wire [0:19] sb_0__1__10_chanx_right_out;
wire [0:19] sb_0__1__10_chany_bottom_out;
wire [0:19] sb_0__1__10_chany_top_out;
wire [0:0] sb_0__1__1_ccff_tail;
wire [0:19] sb_0__1__1_chanx_right_out;
wire [0:19] sb_0__1__1_chany_bottom_out;
wire [0:19] sb_0__1__1_chany_top_out;
wire [0:0] sb_0__1__2_ccff_tail;
wire [0:19] sb_0__1__2_chanx_right_out;
wire [0:19] sb_0__1__2_chany_bottom_out;
wire [0:19] sb_0__1__2_chany_top_out;
wire [0:0] sb_0__1__3_ccff_tail;
wire [0:19] sb_0__1__3_chanx_right_out;
wire [0:19] sb_0__1__3_chany_bottom_out;
wire [0:19] sb_0__1__3_chany_top_out;
wire [0:0] sb_0__1__4_ccff_tail;
wire [0:19] sb_0__1__4_chanx_right_out;
wire [0:19] sb_0__1__4_chany_bottom_out;
wire [0:19] sb_0__1__4_chany_top_out;
wire [0:0] sb_0__1__5_ccff_tail;
wire [0:19] sb_0__1__5_chanx_right_out;
wire [0:19] sb_0__1__5_chany_bottom_out;
wire [0:19] sb_0__1__5_chany_top_out;
wire [0:0] sb_0__1__6_ccff_tail;
wire [0:19] sb_0__1__6_chanx_right_out;
wire [0:19] sb_0__1__6_chany_bottom_out;
wire [0:19] sb_0__1__6_chany_top_out;
wire [0:0] sb_0__1__7_ccff_tail;
wire [0:19] sb_0__1__7_chanx_right_out;
wire [0:19] sb_0__1__7_chany_bottom_out;
wire [0:19] sb_0__1__7_chany_top_out;
wire [0:0] sb_0__1__8_ccff_tail;
wire [0:19] sb_0__1__8_chanx_right_out;
wire [0:19] sb_0__1__8_chany_bottom_out;
wire [0:19] sb_0__1__8_chany_top_out;
wire [0:0] sb_0__1__9_ccff_tail;
wire [0:19] sb_0__1__9_chanx_right_out;
wire [0:19] sb_0__1__9_chany_bottom_out;
wire [0:19] sb_0__1__9_chany_top_out;
wire [0:0] sb_12__0__0_ccff_tail;
wire [0:19] sb_12__0__0_chanx_left_out;
wire [0:19] sb_12__0__0_chany_top_out;
wire [0:0] sb_12__12__0_ccff_tail;
wire [0:19] sb_12__12__0_chanx_left_out;
wire [0:19] sb_12__12__0_chany_bottom_out;
wire [0:0] sb_12__1__0_ccff_tail;
wire [0:19] sb_12__1__0_chanx_left_out;
wire [0:19] sb_12__1__0_chany_bottom_out;
wire [0:19] sb_12__1__0_chany_top_out;
wire [0:0] sb_12__1__10_ccff_tail;
wire [0:19] sb_12__1__10_chanx_left_out;
wire [0:19] sb_12__1__10_chany_bottom_out;
wire [0:19] sb_12__1__10_chany_top_out;
wire [0:0] sb_12__1__1_ccff_tail;
wire [0:19] sb_12__1__1_chanx_left_out;
wire [0:19] sb_12__1__1_chany_bottom_out;
wire [0:19] sb_12__1__1_chany_top_out;
wire [0:0] sb_12__1__2_ccff_tail;
wire [0:19] sb_12__1__2_chanx_left_out;
wire [0:19] sb_12__1__2_chany_bottom_out;
wire [0:19] sb_12__1__2_chany_top_out;
wire [0:0] sb_12__1__3_ccff_tail;
wire [0:19] sb_12__1__3_chanx_left_out;
wire [0:19] sb_12__1__3_chany_bottom_out;
wire [0:19] sb_12__1__3_chany_top_out;
wire [0:0] sb_12__1__4_ccff_tail;
wire [0:19] sb_12__1__4_chanx_left_out;
wire [0:19] sb_12__1__4_chany_bottom_out;
wire [0:19] sb_12__1__4_chany_top_out;
wire [0:0] sb_12__1__5_ccff_tail;
wire [0:19] sb_12__1__5_chanx_left_out;
wire [0:19] sb_12__1__5_chany_bottom_out;
wire [0:19] sb_12__1__5_chany_top_out;
wire [0:0] sb_12__1__6_ccff_tail;
wire [0:19] sb_12__1__6_chanx_left_out;
wire [0:19] sb_12__1__6_chany_bottom_out;
wire [0:19] sb_12__1__6_chany_top_out;
wire [0:0] sb_12__1__7_ccff_tail;
wire [0:19] sb_12__1__7_chanx_left_out;
wire [0:19] sb_12__1__7_chany_bottom_out;
wire [0:19] sb_12__1__7_chany_top_out;
wire [0:0] sb_12__1__8_ccff_tail;
wire [0:19] sb_12__1__8_chanx_left_out;
wire [0:19] sb_12__1__8_chany_bottom_out;
wire [0:19] sb_12__1__8_chany_top_out;
wire [0:0] sb_12__1__9_ccff_tail;
wire [0:19] sb_12__1__9_chanx_left_out;
wire [0:19] sb_12__1__9_chany_bottom_out;
wire [0:19] sb_12__1__9_chany_top_out;
wire [0:0] sb_1__0__0_ccff_tail;
wire [0:19] sb_1__0__0_chanx_left_out;
wire [0:19] sb_1__0__0_chanx_right_out;
wire [0:19] sb_1__0__0_chany_top_out;
wire [0:0] sb_1__0__10_ccff_tail;
wire [0:19] sb_1__0__10_chanx_left_out;
wire [0:19] sb_1__0__10_chanx_right_out;
wire [0:19] sb_1__0__10_chany_top_out;
wire [0:0] sb_1__0__1_ccff_tail;
wire [0:19] sb_1__0__1_chanx_left_out;
wire [0:19] sb_1__0__1_chanx_right_out;
wire [0:19] sb_1__0__1_chany_top_out;
wire [0:0] sb_1__0__2_ccff_tail;
wire [0:19] sb_1__0__2_chanx_left_out;
wire [0:19] sb_1__0__2_chanx_right_out;
wire [0:19] sb_1__0__2_chany_top_out;
wire [0:0] sb_1__0__3_ccff_tail;
wire [0:19] sb_1__0__3_chanx_left_out;
wire [0:19] sb_1__0__3_chanx_right_out;
wire [0:19] sb_1__0__3_chany_top_out;
wire [0:0] sb_1__0__4_ccff_tail;
wire [0:19] sb_1__0__4_chanx_left_out;
wire [0:19] sb_1__0__4_chanx_right_out;
wire [0:19] sb_1__0__4_chany_top_out;
wire [0:0] sb_1__0__5_ccff_tail;
wire [0:19] sb_1__0__5_chanx_left_out;
wire [0:19] sb_1__0__5_chanx_right_out;
wire [0:19] sb_1__0__5_chany_top_out;
wire [0:0] sb_1__0__6_ccff_tail;
wire [0:19] sb_1__0__6_chanx_left_out;
wire [0:19] sb_1__0__6_chanx_right_out;
wire [0:19] sb_1__0__6_chany_top_out;
wire [0:0] sb_1__0__7_ccff_tail;
wire [0:19] sb_1__0__7_chanx_left_out;
wire [0:19] sb_1__0__7_chanx_right_out;
wire [0:19] sb_1__0__7_chany_top_out;
wire [0:0] sb_1__0__8_ccff_tail;
wire [0:19] sb_1__0__8_chanx_left_out;
wire [0:19] sb_1__0__8_chanx_right_out;
wire [0:19] sb_1__0__8_chany_top_out;
wire [0:0] sb_1__0__9_ccff_tail;
wire [0:19] sb_1__0__9_chanx_left_out;
wire [0:19] sb_1__0__9_chanx_right_out;
wire [0:19] sb_1__0__9_chany_top_out;
wire [0:0] sb_1__12__0_ccff_tail;
wire [0:19] sb_1__12__0_chanx_left_out;
wire [0:19] sb_1__12__0_chanx_right_out;
wire [0:19] sb_1__12__0_chany_bottom_out;
wire [0:0] sb_1__12__10_ccff_tail;
wire [0:19] sb_1__12__10_chanx_left_out;
wire [0:19] sb_1__12__10_chanx_right_out;
wire [0:19] sb_1__12__10_chany_bottom_out;
wire [0:0] sb_1__12__1_ccff_tail;
wire [0:19] sb_1__12__1_chanx_left_out;
wire [0:19] sb_1__12__1_chanx_right_out;
wire [0:19] sb_1__12__1_chany_bottom_out;
wire [0:0] sb_1__12__2_ccff_tail;
wire [0:19] sb_1__12__2_chanx_left_out;
wire [0:19] sb_1__12__2_chanx_right_out;
wire [0:19] sb_1__12__2_chany_bottom_out;
wire [0:0] sb_1__12__3_ccff_tail;
wire [0:19] sb_1__12__3_chanx_left_out;
wire [0:19] sb_1__12__3_chanx_right_out;
wire [0:19] sb_1__12__3_chany_bottom_out;
wire [0:0] sb_1__12__4_ccff_tail;
wire [0:19] sb_1__12__4_chanx_left_out;
wire [0:19] sb_1__12__4_chanx_right_out;
wire [0:19] sb_1__12__4_chany_bottom_out;
wire [0:0] sb_1__12__5_ccff_tail;
wire [0:19] sb_1__12__5_chanx_left_out;
wire [0:19] sb_1__12__5_chanx_right_out;
wire [0:19] sb_1__12__5_chany_bottom_out;
wire [0:0] sb_1__12__6_ccff_tail;
wire [0:19] sb_1__12__6_chanx_left_out;
wire [0:19] sb_1__12__6_chanx_right_out;
wire [0:19] sb_1__12__6_chany_bottom_out;
wire [0:0] sb_1__12__7_ccff_tail;
wire [0:19] sb_1__12__7_chanx_left_out;
wire [0:19] sb_1__12__7_chanx_right_out;
wire [0:19] sb_1__12__7_chany_bottom_out;
wire [0:0] sb_1__12__8_ccff_tail;
wire [0:19] sb_1__12__8_chanx_left_out;
wire [0:19] sb_1__12__8_chanx_right_out;
wire [0:19] sb_1__12__8_chany_bottom_out;
wire [0:0] sb_1__12__9_ccff_tail;
wire [0:19] sb_1__12__9_chanx_left_out;
wire [0:19] sb_1__12__9_chanx_right_out;
wire [0:19] sb_1__12__9_chany_bottom_out;
wire [0:0] sb_1__1__0_ccff_tail;
wire [0:19] sb_1__1__0_chanx_left_out;
wire [0:19] sb_1__1__0_chanx_right_out;
wire [0:19] sb_1__1__0_chany_bottom_out;
wire [0:19] sb_1__1__0_chany_top_out;
wire [0:0] sb_1__1__100_ccff_tail;
wire [0:19] sb_1__1__100_chanx_left_out;
wire [0:19] sb_1__1__100_chanx_right_out;
wire [0:19] sb_1__1__100_chany_bottom_out;
wire [0:19] sb_1__1__100_chany_top_out;
wire [0:0] sb_1__1__101_ccff_tail;
wire [0:19] sb_1__1__101_chanx_left_out;
wire [0:19] sb_1__1__101_chanx_right_out;
wire [0:19] sb_1__1__101_chany_bottom_out;
wire [0:19] sb_1__1__101_chany_top_out;
wire [0:0] sb_1__1__102_ccff_tail;
wire [0:19] sb_1__1__102_chanx_left_out;
wire [0:19] sb_1__1__102_chanx_right_out;
wire [0:19] sb_1__1__102_chany_bottom_out;
wire [0:19] sb_1__1__102_chany_top_out;
wire [0:0] sb_1__1__103_ccff_tail;
wire [0:19] sb_1__1__103_chanx_left_out;
wire [0:19] sb_1__1__103_chanx_right_out;
wire [0:19] sb_1__1__103_chany_bottom_out;
wire [0:19] sb_1__1__103_chany_top_out;
wire [0:0] sb_1__1__104_ccff_tail;
wire [0:19] sb_1__1__104_chanx_left_out;
wire [0:19] sb_1__1__104_chanx_right_out;
wire [0:19] sb_1__1__104_chany_bottom_out;
wire [0:19] sb_1__1__104_chany_top_out;
wire [0:0] sb_1__1__105_ccff_tail;
wire [0:19] sb_1__1__105_chanx_left_out;
wire [0:19] sb_1__1__105_chanx_right_out;
wire [0:19] sb_1__1__105_chany_bottom_out;
wire [0:19] sb_1__1__105_chany_top_out;
wire [0:0] sb_1__1__106_ccff_tail;
wire [0:19] sb_1__1__106_chanx_left_out;
wire [0:19] sb_1__1__106_chanx_right_out;
wire [0:19] sb_1__1__106_chany_bottom_out;
wire [0:19] sb_1__1__106_chany_top_out;
wire [0:0] sb_1__1__107_ccff_tail;
wire [0:19] sb_1__1__107_chanx_left_out;
wire [0:19] sb_1__1__107_chanx_right_out;
wire [0:19] sb_1__1__107_chany_bottom_out;
wire [0:19] sb_1__1__107_chany_top_out;
wire [0:0] sb_1__1__108_ccff_tail;
wire [0:19] sb_1__1__108_chanx_left_out;
wire [0:19] sb_1__1__108_chanx_right_out;
wire [0:19] sb_1__1__108_chany_bottom_out;
wire [0:19] sb_1__1__108_chany_top_out;
wire [0:0] sb_1__1__109_ccff_tail;
wire [0:19] sb_1__1__109_chanx_left_out;
wire [0:19] sb_1__1__109_chanx_right_out;
wire [0:19] sb_1__1__109_chany_bottom_out;
wire [0:19] sb_1__1__109_chany_top_out;
wire [0:0] sb_1__1__10_ccff_tail;
wire [0:19] sb_1__1__10_chanx_left_out;
wire [0:19] sb_1__1__10_chanx_right_out;
wire [0:19] sb_1__1__10_chany_bottom_out;
wire [0:19] sb_1__1__10_chany_top_out;
wire [0:0] sb_1__1__110_ccff_tail;
wire [0:19] sb_1__1__110_chanx_left_out;
wire [0:19] sb_1__1__110_chanx_right_out;
wire [0:19] sb_1__1__110_chany_bottom_out;
wire [0:19] sb_1__1__110_chany_top_out;
wire [0:0] sb_1__1__111_ccff_tail;
wire [0:19] sb_1__1__111_chanx_left_out;
wire [0:19] sb_1__1__111_chanx_right_out;
wire [0:19] sb_1__1__111_chany_bottom_out;
wire [0:19] sb_1__1__111_chany_top_out;
wire [0:0] sb_1__1__112_ccff_tail;
wire [0:19] sb_1__1__112_chanx_left_out;
wire [0:19] sb_1__1__112_chanx_right_out;
wire [0:19] sb_1__1__112_chany_bottom_out;
wire [0:19] sb_1__1__112_chany_top_out;
wire [0:0] sb_1__1__113_ccff_tail;
wire [0:19] sb_1__1__113_chanx_left_out;
wire [0:19] sb_1__1__113_chanx_right_out;
wire [0:19] sb_1__1__113_chany_bottom_out;
wire [0:19] sb_1__1__113_chany_top_out;
wire [0:0] sb_1__1__114_ccff_tail;
wire [0:19] sb_1__1__114_chanx_left_out;
wire [0:19] sb_1__1__114_chanx_right_out;
wire [0:19] sb_1__1__114_chany_bottom_out;
wire [0:19] sb_1__1__114_chany_top_out;
wire [0:0] sb_1__1__115_ccff_tail;
wire [0:19] sb_1__1__115_chanx_left_out;
wire [0:19] sb_1__1__115_chanx_right_out;
wire [0:19] sb_1__1__115_chany_bottom_out;
wire [0:19] sb_1__1__115_chany_top_out;
wire [0:0] sb_1__1__116_ccff_tail;
wire [0:19] sb_1__1__116_chanx_left_out;
wire [0:19] sb_1__1__116_chanx_right_out;
wire [0:19] sb_1__1__116_chany_bottom_out;
wire [0:19] sb_1__1__116_chany_top_out;
wire [0:0] sb_1__1__117_ccff_tail;
wire [0:19] sb_1__1__117_chanx_left_out;
wire [0:19] sb_1__1__117_chanx_right_out;
wire [0:19] sb_1__1__117_chany_bottom_out;
wire [0:19] sb_1__1__117_chany_top_out;
wire [0:0] sb_1__1__118_ccff_tail;
wire [0:19] sb_1__1__118_chanx_left_out;
wire [0:19] sb_1__1__118_chanx_right_out;
wire [0:19] sb_1__1__118_chany_bottom_out;
wire [0:19] sb_1__1__118_chany_top_out;
wire [0:0] sb_1__1__119_ccff_tail;
wire [0:19] sb_1__1__119_chanx_left_out;
wire [0:19] sb_1__1__119_chanx_right_out;
wire [0:19] sb_1__1__119_chany_bottom_out;
wire [0:19] sb_1__1__119_chany_top_out;
wire [0:0] sb_1__1__11_ccff_tail;
wire [0:19] sb_1__1__11_chanx_left_out;
wire [0:19] sb_1__1__11_chanx_right_out;
wire [0:19] sb_1__1__11_chany_bottom_out;
wire [0:19] sb_1__1__11_chany_top_out;
wire [0:0] sb_1__1__120_ccff_tail;
wire [0:19] sb_1__1__120_chanx_left_out;
wire [0:19] sb_1__1__120_chanx_right_out;
wire [0:19] sb_1__1__120_chany_bottom_out;
wire [0:19] sb_1__1__120_chany_top_out;
wire [0:0] sb_1__1__12_ccff_tail;
wire [0:19] sb_1__1__12_chanx_left_out;
wire [0:19] sb_1__1__12_chanx_right_out;
wire [0:19] sb_1__1__12_chany_bottom_out;
wire [0:19] sb_1__1__12_chany_top_out;
wire [0:0] sb_1__1__13_ccff_tail;
wire [0:19] sb_1__1__13_chanx_left_out;
wire [0:19] sb_1__1__13_chanx_right_out;
wire [0:19] sb_1__1__13_chany_bottom_out;
wire [0:19] sb_1__1__13_chany_top_out;
wire [0:0] sb_1__1__14_ccff_tail;
wire [0:19] sb_1__1__14_chanx_left_out;
wire [0:19] sb_1__1__14_chanx_right_out;
wire [0:19] sb_1__1__14_chany_bottom_out;
wire [0:19] sb_1__1__14_chany_top_out;
wire [0:0] sb_1__1__15_ccff_tail;
wire [0:19] sb_1__1__15_chanx_left_out;
wire [0:19] sb_1__1__15_chanx_right_out;
wire [0:19] sb_1__1__15_chany_bottom_out;
wire [0:19] sb_1__1__15_chany_top_out;
wire [0:0] sb_1__1__16_ccff_tail;
wire [0:19] sb_1__1__16_chanx_left_out;
wire [0:19] sb_1__1__16_chanx_right_out;
wire [0:19] sb_1__1__16_chany_bottom_out;
wire [0:19] sb_1__1__16_chany_top_out;
wire [0:0] sb_1__1__17_ccff_tail;
wire [0:19] sb_1__1__17_chanx_left_out;
wire [0:19] sb_1__1__17_chanx_right_out;
wire [0:19] sb_1__1__17_chany_bottom_out;
wire [0:19] sb_1__1__17_chany_top_out;
wire [0:0] sb_1__1__18_ccff_tail;
wire [0:19] sb_1__1__18_chanx_left_out;
wire [0:19] sb_1__1__18_chanx_right_out;
wire [0:19] sb_1__1__18_chany_bottom_out;
wire [0:19] sb_1__1__18_chany_top_out;
wire [0:0] sb_1__1__19_ccff_tail;
wire [0:19] sb_1__1__19_chanx_left_out;
wire [0:19] sb_1__1__19_chanx_right_out;
wire [0:19] sb_1__1__19_chany_bottom_out;
wire [0:19] sb_1__1__19_chany_top_out;
wire [0:0] sb_1__1__1_ccff_tail;
wire [0:19] sb_1__1__1_chanx_left_out;
wire [0:19] sb_1__1__1_chanx_right_out;
wire [0:19] sb_1__1__1_chany_bottom_out;
wire [0:19] sb_1__1__1_chany_top_out;
wire [0:0] sb_1__1__20_ccff_tail;
wire [0:19] sb_1__1__20_chanx_left_out;
wire [0:19] sb_1__1__20_chanx_right_out;
wire [0:19] sb_1__1__20_chany_bottom_out;
wire [0:19] sb_1__1__20_chany_top_out;
wire [0:0] sb_1__1__21_ccff_tail;
wire [0:19] sb_1__1__21_chanx_left_out;
wire [0:19] sb_1__1__21_chanx_right_out;
wire [0:19] sb_1__1__21_chany_bottom_out;
wire [0:19] sb_1__1__21_chany_top_out;
wire [0:0] sb_1__1__22_ccff_tail;
wire [0:19] sb_1__1__22_chanx_left_out;
wire [0:19] sb_1__1__22_chanx_right_out;
wire [0:19] sb_1__1__22_chany_bottom_out;
wire [0:19] sb_1__1__22_chany_top_out;
wire [0:0] sb_1__1__23_ccff_tail;
wire [0:19] sb_1__1__23_chanx_left_out;
wire [0:19] sb_1__1__23_chanx_right_out;
wire [0:19] sb_1__1__23_chany_bottom_out;
wire [0:19] sb_1__1__23_chany_top_out;
wire [0:0] sb_1__1__24_ccff_tail;
wire [0:19] sb_1__1__24_chanx_left_out;
wire [0:19] sb_1__1__24_chanx_right_out;
wire [0:19] sb_1__1__24_chany_bottom_out;
wire [0:19] sb_1__1__24_chany_top_out;
wire [0:0] sb_1__1__25_ccff_tail;
wire [0:19] sb_1__1__25_chanx_left_out;
wire [0:19] sb_1__1__25_chanx_right_out;
wire [0:19] sb_1__1__25_chany_bottom_out;
wire [0:19] sb_1__1__25_chany_top_out;
wire [0:0] sb_1__1__26_ccff_tail;
wire [0:19] sb_1__1__26_chanx_left_out;
wire [0:19] sb_1__1__26_chanx_right_out;
wire [0:19] sb_1__1__26_chany_bottom_out;
wire [0:19] sb_1__1__26_chany_top_out;
wire [0:0] sb_1__1__27_ccff_tail;
wire [0:19] sb_1__1__27_chanx_left_out;
wire [0:19] sb_1__1__27_chanx_right_out;
wire [0:19] sb_1__1__27_chany_bottom_out;
wire [0:19] sb_1__1__27_chany_top_out;
wire [0:0] sb_1__1__28_ccff_tail;
wire [0:19] sb_1__1__28_chanx_left_out;
wire [0:19] sb_1__1__28_chanx_right_out;
wire [0:19] sb_1__1__28_chany_bottom_out;
wire [0:19] sb_1__1__28_chany_top_out;
wire [0:0] sb_1__1__29_ccff_tail;
wire [0:19] sb_1__1__29_chanx_left_out;
wire [0:19] sb_1__1__29_chanx_right_out;
wire [0:19] sb_1__1__29_chany_bottom_out;
wire [0:19] sb_1__1__29_chany_top_out;
wire [0:0] sb_1__1__2_ccff_tail;
wire [0:19] sb_1__1__2_chanx_left_out;
wire [0:19] sb_1__1__2_chanx_right_out;
wire [0:19] sb_1__1__2_chany_bottom_out;
wire [0:19] sb_1__1__2_chany_top_out;
wire [0:0] sb_1__1__30_ccff_tail;
wire [0:19] sb_1__1__30_chanx_left_out;
wire [0:19] sb_1__1__30_chanx_right_out;
wire [0:19] sb_1__1__30_chany_bottom_out;
wire [0:19] sb_1__1__30_chany_top_out;
wire [0:0] sb_1__1__31_ccff_tail;
wire [0:19] sb_1__1__31_chanx_left_out;
wire [0:19] sb_1__1__31_chanx_right_out;
wire [0:19] sb_1__1__31_chany_bottom_out;
wire [0:19] sb_1__1__31_chany_top_out;
wire [0:0] sb_1__1__32_ccff_tail;
wire [0:19] sb_1__1__32_chanx_left_out;
wire [0:19] sb_1__1__32_chanx_right_out;
wire [0:19] sb_1__1__32_chany_bottom_out;
wire [0:19] sb_1__1__32_chany_top_out;
wire [0:0] sb_1__1__33_ccff_tail;
wire [0:19] sb_1__1__33_chanx_left_out;
wire [0:19] sb_1__1__33_chanx_right_out;
wire [0:19] sb_1__1__33_chany_bottom_out;
wire [0:19] sb_1__1__33_chany_top_out;
wire [0:0] sb_1__1__34_ccff_tail;
wire [0:19] sb_1__1__34_chanx_left_out;
wire [0:19] sb_1__1__34_chanx_right_out;
wire [0:19] sb_1__1__34_chany_bottom_out;
wire [0:19] sb_1__1__34_chany_top_out;
wire [0:0] sb_1__1__35_ccff_tail;
wire [0:19] sb_1__1__35_chanx_left_out;
wire [0:19] sb_1__1__35_chanx_right_out;
wire [0:19] sb_1__1__35_chany_bottom_out;
wire [0:19] sb_1__1__35_chany_top_out;
wire [0:0] sb_1__1__36_ccff_tail;
wire [0:19] sb_1__1__36_chanx_left_out;
wire [0:19] sb_1__1__36_chanx_right_out;
wire [0:19] sb_1__1__36_chany_bottom_out;
wire [0:19] sb_1__1__36_chany_top_out;
wire [0:0] sb_1__1__37_ccff_tail;
wire [0:19] sb_1__1__37_chanx_left_out;
wire [0:19] sb_1__1__37_chanx_right_out;
wire [0:19] sb_1__1__37_chany_bottom_out;
wire [0:19] sb_1__1__37_chany_top_out;
wire [0:0] sb_1__1__38_ccff_tail;
wire [0:19] sb_1__1__38_chanx_left_out;
wire [0:19] sb_1__1__38_chanx_right_out;
wire [0:19] sb_1__1__38_chany_bottom_out;
wire [0:19] sb_1__1__38_chany_top_out;
wire [0:0] sb_1__1__39_ccff_tail;
wire [0:19] sb_1__1__39_chanx_left_out;
wire [0:19] sb_1__1__39_chanx_right_out;
wire [0:19] sb_1__1__39_chany_bottom_out;
wire [0:19] sb_1__1__39_chany_top_out;
wire [0:0] sb_1__1__3_ccff_tail;
wire [0:19] sb_1__1__3_chanx_left_out;
wire [0:19] sb_1__1__3_chanx_right_out;
wire [0:19] sb_1__1__3_chany_bottom_out;
wire [0:19] sb_1__1__3_chany_top_out;
wire [0:0] sb_1__1__40_ccff_tail;
wire [0:19] sb_1__1__40_chanx_left_out;
wire [0:19] sb_1__1__40_chanx_right_out;
wire [0:19] sb_1__1__40_chany_bottom_out;
wire [0:19] sb_1__1__40_chany_top_out;
wire [0:0] sb_1__1__41_ccff_tail;
wire [0:19] sb_1__1__41_chanx_left_out;
wire [0:19] sb_1__1__41_chanx_right_out;
wire [0:19] sb_1__1__41_chany_bottom_out;
wire [0:19] sb_1__1__41_chany_top_out;
wire [0:0] sb_1__1__42_ccff_tail;
wire [0:19] sb_1__1__42_chanx_left_out;
wire [0:19] sb_1__1__42_chanx_right_out;
wire [0:19] sb_1__1__42_chany_bottom_out;
wire [0:19] sb_1__1__42_chany_top_out;
wire [0:0] sb_1__1__43_ccff_tail;
wire [0:19] sb_1__1__43_chanx_left_out;
wire [0:19] sb_1__1__43_chanx_right_out;
wire [0:19] sb_1__1__43_chany_bottom_out;
wire [0:19] sb_1__1__43_chany_top_out;
wire [0:0] sb_1__1__44_ccff_tail;
wire [0:19] sb_1__1__44_chanx_left_out;
wire [0:19] sb_1__1__44_chanx_right_out;
wire [0:19] sb_1__1__44_chany_bottom_out;
wire [0:19] sb_1__1__44_chany_top_out;
wire [0:0] sb_1__1__45_ccff_tail;
wire [0:19] sb_1__1__45_chanx_left_out;
wire [0:19] sb_1__1__45_chanx_right_out;
wire [0:19] sb_1__1__45_chany_bottom_out;
wire [0:19] sb_1__1__45_chany_top_out;
wire [0:0] sb_1__1__46_ccff_tail;
wire [0:19] sb_1__1__46_chanx_left_out;
wire [0:19] sb_1__1__46_chanx_right_out;
wire [0:19] sb_1__1__46_chany_bottom_out;
wire [0:19] sb_1__1__46_chany_top_out;
wire [0:0] sb_1__1__47_ccff_tail;
wire [0:19] sb_1__1__47_chanx_left_out;
wire [0:19] sb_1__1__47_chanx_right_out;
wire [0:19] sb_1__1__47_chany_bottom_out;
wire [0:19] sb_1__1__47_chany_top_out;
wire [0:0] sb_1__1__48_ccff_tail;
wire [0:19] sb_1__1__48_chanx_left_out;
wire [0:19] sb_1__1__48_chanx_right_out;
wire [0:19] sb_1__1__48_chany_bottom_out;
wire [0:19] sb_1__1__48_chany_top_out;
wire [0:0] sb_1__1__49_ccff_tail;
wire [0:19] sb_1__1__49_chanx_left_out;
wire [0:19] sb_1__1__49_chanx_right_out;
wire [0:19] sb_1__1__49_chany_bottom_out;
wire [0:19] sb_1__1__49_chany_top_out;
wire [0:0] sb_1__1__4_ccff_tail;
wire [0:19] sb_1__1__4_chanx_left_out;
wire [0:19] sb_1__1__4_chanx_right_out;
wire [0:19] sb_1__1__4_chany_bottom_out;
wire [0:19] sb_1__1__4_chany_top_out;
wire [0:0] sb_1__1__50_ccff_tail;
wire [0:19] sb_1__1__50_chanx_left_out;
wire [0:19] sb_1__1__50_chanx_right_out;
wire [0:19] sb_1__1__50_chany_bottom_out;
wire [0:19] sb_1__1__50_chany_top_out;
wire [0:0] sb_1__1__51_ccff_tail;
wire [0:19] sb_1__1__51_chanx_left_out;
wire [0:19] sb_1__1__51_chanx_right_out;
wire [0:19] sb_1__1__51_chany_bottom_out;
wire [0:19] sb_1__1__51_chany_top_out;
wire [0:0] sb_1__1__52_ccff_tail;
wire [0:19] sb_1__1__52_chanx_left_out;
wire [0:19] sb_1__1__52_chanx_right_out;
wire [0:19] sb_1__1__52_chany_bottom_out;
wire [0:19] sb_1__1__52_chany_top_out;
wire [0:0] sb_1__1__53_ccff_tail;
wire [0:19] sb_1__1__53_chanx_left_out;
wire [0:19] sb_1__1__53_chanx_right_out;
wire [0:19] sb_1__1__53_chany_bottom_out;
wire [0:19] sb_1__1__53_chany_top_out;
wire [0:0] sb_1__1__54_ccff_tail;
wire [0:19] sb_1__1__54_chanx_left_out;
wire [0:19] sb_1__1__54_chanx_right_out;
wire [0:19] sb_1__1__54_chany_bottom_out;
wire [0:19] sb_1__1__54_chany_top_out;
wire [0:0] sb_1__1__55_ccff_tail;
wire [0:19] sb_1__1__55_chanx_left_out;
wire [0:19] sb_1__1__55_chanx_right_out;
wire [0:19] sb_1__1__55_chany_bottom_out;
wire [0:19] sb_1__1__55_chany_top_out;
wire [0:0] sb_1__1__56_ccff_tail;
wire [0:19] sb_1__1__56_chanx_left_out;
wire [0:19] sb_1__1__56_chanx_right_out;
wire [0:19] sb_1__1__56_chany_bottom_out;
wire [0:19] sb_1__1__56_chany_top_out;
wire [0:0] sb_1__1__57_ccff_tail;
wire [0:19] sb_1__1__57_chanx_left_out;
wire [0:19] sb_1__1__57_chanx_right_out;
wire [0:19] sb_1__1__57_chany_bottom_out;
wire [0:19] sb_1__1__57_chany_top_out;
wire [0:0] sb_1__1__58_ccff_tail;
wire [0:19] sb_1__1__58_chanx_left_out;
wire [0:19] sb_1__1__58_chanx_right_out;
wire [0:19] sb_1__1__58_chany_bottom_out;
wire [0:19] sb_1__1__58_chany_top_out;
wire [0:0] sb_1__1__59_ccff_tail;
wire [0:19] sb_1__1__59_chanx_left_out;
wire [0:19] sb_1__1__59_chanx_right_out;
wire [0:19] sb_1__1__59_chany_bottom_out;
wire [0:19] sb_1__1__59_chany_top_out;
wire [0:0] sb_1__1__5_ccff_tail;
wire [0:19] sb_1__1__5_chanx_left_out;
wire [0:19] sb_1__1__5_chanx_right_out;
wire [0:19] sb_1__1__5_chany_bottom_out;
wire [0:19] sb_1__1__5_chany_top_out;
wire [0:0] sb_1__1__60_ccff_tail;
wire [0:19] sb_1__1__60_chanx_left_out;
wire [0:19] sb_1__1__60_chanx_right_out;
wire [0:19] sb_1__1__60_chany_bottom_out;
wire [0:19] sb_1__1__60_chany_top_out;
wire [0:0] sb_1__1__61_ccff_tail;
wire [0:19] sb_1__1__61_chanx_left_out;
wire [0:19] sb_1__1__61_chanx_right_out;
wire [0:19] sb_1__1__61_chany_bottom_out;
wire [0:19] sb_1__1__61_chany_top_out;
wire [0:0] sb_1__1__62_ccff_tail;
wire [0:19] sb_1__1__62_chanx_left_out;
wire [0:19] sb_1__1__62_chanx_right_out;
wire [0:19] sb_1__1__62_chany_bottom_out;
wire [0:19] sb_1__1__62_chany_top_out;
wire [0:0] sb_1__1__63_ccff_tail;
wire [0:19] sb_1__1__63_chanx_left_out;
wire [0:19] sb_1__1__63_chanx_right_out;
wire [0:19] sb_1__1__63_chany_bottom_out;
wire [0:19] sb_1__1__63_chany_top_out;
wire [0:0] sb_1__1__64_ccff_tail;
wire [0:19] sb_1__1__64_chanx_left_out;
wire [0:19] sb_1__1__64_chanx_right_out;
wire [0:19] sb_1__1__64_chany_bottom_out;
wire [0:19] sb_1__1__64_chany_top_out;
wire [0:0] sb_1__1__65_ccff_tail;
wire [0:19] sb_1__1__65_chanx_left_out;
wire [0:19] sb_1__1__65_chanx_right_out;
wire [0:19] sb_1__1__65_chany_bottom_out;
wire [0:19] sb_1__1__65_chany_top_out;
wire [0:0] sb_1__1__66_ccff_tail;
wire [0:19] sb_1__1__66_chanx_left_out;
wire [0:19] sb_1__1__66_chanx_right_out;
wire [0:19] sb_1__1__66_chany_bottom_out;
wire [0:19] sb_1__1__66_chany_top_out;
wire [0:0] sb_1__1__67_ccff_tail;
wire [0:19] sb_1__1__67_chanx_left_out;
wire [0:19] sb_1__1__67_chanx_right_out;
wire [0:19] sb_1__1__67_chany_bottom_out;
wire [0:19] sb_1__1__67_chany_top_out;
wire [0:0] sb_1__1__68_ccff_tail;
wire [0:19] sb_1__1__68_chanx_left_out;
wire [0:19] sb_1__1__68_chanx_right_out;
wire [0:19] sb_1__1__68_chany_bottom_out;
wire [0:19] sb_1__1__68_chany_top_out;
wire [0:0] sb_1__1__69_ccff_tail;
wire [0:19] sb_1__1__69_chanx_left_out;
wire [0:19] sb_1__1__69_chanx_right_out;
wire [0:19] sb_1__1__69_chany_bottom_out;
wire [0:19] sb_1__1__69_chany_top_out;
wire [0:0] sb_1__1__6_ccff_tail;
wire [0:19] sb_1__1__6_chanx_left_out;
wire [0:19] sb_1__1__6_chanx_right_out;
wire [0:19] sb_1__1__6_chany_bottom_out;
wire [0:19] sb_1__1__6_chany_top_out;
wire [0:0] sb_1__1__70_ccff_tail;
wire [0:19] sb_1__1__70_chanx_left_out;
wire [0:19] sb_1__1__70_chanx_right_out;
wire [0:19] sb_1__1__70_chany_bottom_out;
wire [0:19] sb_1__1__70_chany_top_out;
wire [0:0] sb_1__1__71_ccff_tail;
wire [0:19] sb_1__1__71_chanx_left_out;
wire [0:19] sb_1__1__71_chanx_right_out;
wire [0:19] sb_1__1__71_chany_bottom_out;
wire [0:19] sb_1__1__71_chany_top_out;
wire [0:0] sb_1__1__72_ccff_tail;
wire [0:19] sb_1__1__72_chanx_left_out;
wire [0:19] sb_1__1__72_chanx_right_out;
wire [0:19] sb_1__1__72_chany_bottom_out;
wire [0:19] sb_1__1__72_chany_top_out;
wire [0:0] sb_1__1__73_ccff_tail;
wire [0:19] sb_1__1__73_chanx_left_out;
wire [0:19] sb_1__1__73_chanx_right_out;
wire [0:19] sb_1__1__73_chany_bottom_out;
wire [0:19] sb_1__1__73_chany_top_out;
wire [0:0] sb_1__1__74_ccff_tail;
wire [0:19] sb_1__1__74_chanx_left_out;
wire [0:19] sb_1__1__74_chanx_right_out;
wire [0:19] sb_1__1__74_chany_bottom_out;
wire [0:19] sb_1__1__74_chany_top_out;
wire [0:0] sb_1__1__75_ccff_tail;
wire [0:19] sb_1__1__75_chanx_left_out;
wire [0:19] sb_1__1__75_chanx_right_out;
wire [0:19] sb_1__1__75_chany_bottom_out;
wire [0:19] sb_1__1__75_chany_top_out;
wire [0:0] sb_1__1__76_ccff_tail;
wire [0:19] sb_1__1__76_chanx_left_out;
wire [0:19] sb_1__1__76_chanx_right_out;
wire [0:19] sb_1__1__76_chany_bottom_out;
wire [0:19] sb_1__1__76_chany_top_out;
wire [0:0] sb_1__1__77_ccff_tail;
wire [0:19] sb_1__1__77_chanx_left_out;
wire [0:19] sb_1__1__77_chanx_right_out;
wire [0:19] sb_1__1__77_chany_bottom_out;
wire [0:19] sb_1__1__77_chany_top_out;
wire [0:0] sb_1__1__78_ccff_tail;
wire [0:19] sb_1__1__78_chanx_left_out;
wire [0:19] sb_1__1__78_chanx_right_out;
wire [0:19] sb_1__1__78_chany_bottom_out;
wire [0:19] sb_1__1__78_chany_top_out;
wire [0:0] sb_1__1__79_ccff_tail;
wire [0:19] sb_1__1__79_chanx_left_out;
wire [0:19] sb_1__1__79_chanx_right_out;
wire [0:19] sb_1__1__79_chany_bottom_out;
wire [0:19] sb_1__1__79_chany_top_out;
wire [0:0] sb_1__1__7_ccff_tail;
wire [0:19] sb_1__1__7_chanx_left_out;
wire [0:19] sb_1__1__7_chanx_right_out;
wire [0:19] sb_1__1__7_chany_bottom_out;
wire [0:19] sb_1__1__7_chany_top_out;
wire [0:0] sb_1__1__80_ccff_tail;
wire [0:19] sb_1__1__80_chanx_left_out;
wire [0:19] sb_1__1__80_chanx_right_out;
wire [0:19] sb_1__1__80_chany_bottom_out;
wire [0:19] sb_1__1__80_chany_top_out;
wire [0:0] sb_1__1__81_ccff_tail;
wire [0:19] sb_1__1__81_chanx_left_out;
wire [0:19] sb_1__1__81_chanx_right_out;
wire [0:19] sb_1__1__81_chany_bottom_out;
wire [0:19] sb_1__1__81_chany_top_out;
wire [0:0] sb_1__1__82_ccff_tail;
wire [0:19] sb_1__1__82_chanx_left_out;
wire [0:19] sb_1__1__82_chanx_right_out;
wire [0:19] sb_1__1__82_chany_bottom_out;
wire [0:19] sb_1__1__82_chany_top_out;
wire [0:0] sb_1__1__83_ccff_tail;
wire [0:19] sb_1__1__83_chanx_left_out;
wire [0:19] sb_1__1__83_chanx_right_out;
wire [0:19] sb_1__1__83_chany_bottom_out;
wire [0:19] sb_1__1__83_chany_top_out;
wire [0:0] sb_1__1__84_ccff_tail;
wire [0:19] sb_1__1__84_chanx_left_out;
wire [0:19] sb_1__1__84_chanx_right_out;
wire [0:19] sb_1__1__84_chany_bottom_out;
wire [0:19] sb_1__1__84_chany_top_out;
wire [0:0] sb_1__1__85_ccff_tail;
wire [0:19] sb_1__1__85_chanx_left_out;
wire [0:19] sb_1__1__85_chanx_right_out;
wire [0:19] sb_1__1__85_chany_bottom_out;
wire [0:19] sb_1__1__85_chany_top_out;
wire [0:0] sb_1__1__86_ccff_tail;
wire [0:19] sb_1__1__86_chanx_left_out;
wire [0:19] sb_1__1__86_chanx_right_out;
wire [0:19] sb_1__1__86_chany_bottom_out;
wire [0:19] sb_1__1__86_chany_top_out;
wire [0:0] sb_1__1__87_ccff_tail;
wire [0:19] sb_1__1__87_chanx_left_out;
wire [0:19] sb_1__1__87_chanx_right_out;
wire [0:19] sb_1__1__87_chany_bottom_out;
wire [0:19] sb_1__1__87_chany_top_out;
wire [0:0] sb_1__1__88_ccff_tail;
wire [0:19] sb_1__1__88_chanx_left_out;
wire [0:19] sb_1__1__88_chanx_right_out;
wire [0:19] sb_1__1__88_chany_bottom_out;
wire [0:19] sb_1__1__88_chany_top_out;
wire [0:0] sb_1__1__89_ccff_tail;
wire [0:19] sb_1__1__89_chanx_left_out;
wire [0:19] sb_1__1__89_chanx_right_out;
wire [0:19] sb_1__1__89_chany_bottom_out;
wire [0:19] sb_1__1__89_chany_top_out;
wire [0:0] sb_1__1__8_ccff_tail;
wire [0:19] sb_1__1__8_chanx_left_out;
wire [0:19] sb_1__1__8_chanx_right_out;
wire [0:19] sb_1__1__8_chany_bottom_out;
wire [0:19] sb_1__1__8_chany_top_out;
wire [0:0] sb_1__1__90_ccff_tail;
wire [0:19] sb_1__1__90_chanx_left_out;
wire [0:19] sb_1__1__90_chanx_right_out;
wire [0:19] sb_1__1__90_chany_bottom_out;
wire [0:19] sb_1__1__90_chany_top_out;
wire [0:0] sb_1__1__91_ccff_tail;
wire [0:19] sb_1__1__91_chanx_left_out;
wire [0:19] sb_1__1__91_chanx_right_out;
wire [0:19] sb_1__1__91_chany_bottom_out;
wire [0:19] sb_1__1__91_chany_top_out;
wire [0:0] sb_1__1__92_ccff_tail;
wire [0:19] sb_1__1__92_chanx_left_out;
wire [0:19] sb_1__1__92_chanx_right_out;
wire [0:19] sb_1__1__92_chany_bottom_out;
wire [0:19] sb_1__1__92_chany_top_out;
wire [0:0] sb_1__1__93_ccff_tail;
wire [0:19] sb_1__1__93_chanx_left_out;
wire [0:19] sb_1__1__93_chanx_right_out;
wire [0:19] sb_1__1__93_chany_bottom_out;
wire [0:19] sb_1__1__93_chany_top_out;
wire [0:0] sb_1__1__94_ccff_tail;
wire [0:19] sb_1__1__94_chanx_left_out;
wire [0:19] sb_1__1__94_chanx_right_out;
wire [0:19] sb_1__1__94_chany_bottom_out;
wire [0:19] sb_1__1__94_chany_top_out;
wire [0:0] sb_1__1__95_ccff_tail;
wire [0:19] sb_1__1__95_chanx_left_out;
wire [0:19] sb_1__1__95_chanx_right_out;
wire [0:19] sb_1__1__95_chany_bottom_out;
wire [0:19] sb_1__1__95_chany_top_out;
wire [0:0] sb_1__1__96_ccff_tail;
wire [0:19] sb_1__1__96_chanx_left_out;
wire [0:19] sb_1__1__96_chanx_right_out;
wire [0:19] sb_1__1__96_chany_bottom_out;
wire [0:19] sb_1__1__96_chany_top_out;
wire [0:0] sb_1__1__97_ccff_tail;
wire [0:19] sb_1__1__97_chanx_left_out;
wire [0:19] sb_1__1__97_chanx_right_out;
wire [0:19] sb_1__1__97_chany_bottom_out;
wire [0:19] sb_1__1__97_chany_top_out;
wire [0:0] sb_1__1__98_ccff_tail;
wire [0:19] sb_1__1__98_chanx_left_out;
wire [0:19] sb_1__1__98_chanx_right_out;
wire [0:19] sb_1__1__98_chany_bottom_out;
wire [0:19] sb_1__1__98_chany_top_out;
wire [0:0] sb_1__1__99_ccff_tail;
wire [0:19] sb_1__1__99_chanx_left_out;
wire [0:19] sb_1__1__99_chanx_right_out;
wire [0:19] sb_1__1__99_chany_bottom_out;
wire [0:19] sb_1__1__99_chany_top_out;
wire [0:0] sb_1__1__9_ccff_tail;
wire [0:19] sb_1__1__9_chanx_left_out;
wire [0:19] sb_1__1__9_chanx_right_out;
wire [0:19] sb_1__1__9_chany_bottom_out;
wire [0:19] sb_1__1__9_chany_top_out;

//
//
//
//

	grid_clb grid_clb_1__1_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_0_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_143_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__0_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__0_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__0_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__0_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__0_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__0_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__0_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__0_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__0_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__0_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__0_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__0_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__0_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__0_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__0_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__0_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__0__0_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__0__0_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__0__0_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__0__0_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__0__0_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__0__0_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__0__0_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__0__0_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__0__0_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__0__0_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__0__0_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__0__0_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__0__0_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__0__0_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__0__0_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__0__0_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_0__1__0_right_grid_pin_52_[0]),
		.ccff_head(grid_io_left_0_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_0_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_0_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_0_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_0_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_0_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_0_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_0_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_0_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_0_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_0_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_0_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_0_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_0_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_0_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_0_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_0_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_0_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_0_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_0_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_0_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_0_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_0_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_0_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_0_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_0_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_0_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_0_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_0_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_0_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_0_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_0_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_0_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_0_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_0_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_0_ccff_tail[0]));

	grid_clb grid_clb_1__2_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_1_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_144_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__1_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__1_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__1_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__1_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__1_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__1_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__1_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__1_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__1_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__1_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__1_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__1_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__1_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__1_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__1_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__1_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__0_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__0_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__0_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__0_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__0_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__0_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__0_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__0_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__0_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__0_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__0_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__0_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__0_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__0_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__0_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__0_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_0__1__1_right_grid_pin_52_[0]),
		.ccff_head(grid_io_left_1_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_1_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_1_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_1_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_1_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_1_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_1_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_1_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_1_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_1_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_1_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_1_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_1_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_1_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_1_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_1_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_1_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_1_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_1_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_1_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_1_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_1_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_1_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_1_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_1_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_1_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_1_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_1_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_1_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_1_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_1_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_1_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_1_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_1_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_1_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_1_ccff_tail[0]));

	grid_clb grid_clb_1__3_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_2_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_145_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__2_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__2_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__2_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__2_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__2_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__2_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__2_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__2_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__2_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__2_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__2_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__2_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__2_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__2_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__2_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__2_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__1_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__1_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__1_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__1_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__1_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__1_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__1_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__1_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__1_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__1_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__1_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__1_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__1_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__1_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__1_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__1_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_0__1__2_right_grid_pin_52_[0]),
		.ccff_head(grid_io_left_2_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_2_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_2_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_2_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_2_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_2_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_2_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_2_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_2_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_2_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_2_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_2_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_2_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_2_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_2_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_2_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_2_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_2_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_2_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_2_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_2_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_2_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_2_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_2_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_2_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_2_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_2_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_2_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_2_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_2_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_2_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_2_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_2_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_2_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_2_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_2_ccff_tail[0]));

	grid_clb grid_clb_1__4_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_3_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_146_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__3_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__3_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__3_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__3_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__3_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__3_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__3_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__3_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__3_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__3_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__3_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__3_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__3_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__3_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__3_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__3_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__2_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__2_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__2_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__2_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__2_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__2_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__2_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__2_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__2_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__2_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__2_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__2_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__2_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__2_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__2_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__2_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_0__1__3_right_grid_pin_52_[0]),
		.ccff_head(grid_io_left_3_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_3_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_3_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_3_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_3_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_3_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_3_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_3_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_3_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_3_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_3_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_3_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_3_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_3_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_3_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_3_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_3_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_3_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_3_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_3_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_3_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_3_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_3_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_3_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_3_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_3_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_3_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_3_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_3_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_3_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_3_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_3_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_3_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_3_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_3_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_3_ccff_tail[0]));

	grid_clb grid_clb_1__5_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_4_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_147_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__4_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__4_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__4_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__4_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__4_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__4_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__4_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__4_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__4_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__4_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__4_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__4_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__4_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__4_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__4_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__4_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__3_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__3_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__3_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__3_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__3_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__3_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__3_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__3_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__3_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__3_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__3_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__3_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__3_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__3_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__3_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__3_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_0__1__4_right_grid_pin_52_[0]),
		.ccff_head(grid_io_left_4_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_4_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_4_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_4_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_4_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_4_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_4_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_4_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_4_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_4_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_4_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_4_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_4_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_4_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_4_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_4_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_4_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_4_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_4_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_4_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_4_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_4_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_4_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_4_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_4_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_4_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_4_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_4_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_4_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_4_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_4_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_4_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_4_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_4_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_4_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_4_ccff_tail[0]));

	grid_clb grid_clb_1__6_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_5_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_148_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__5_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__5_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__5_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__5_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__5_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__5_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__5_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__5_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__5_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__5_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__5_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__5_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__5_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__5_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__5_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__5_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__4_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__4_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__4_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__4_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__4_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__4_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__4_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__4_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__4_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__4_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__4_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__4_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__4_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__4_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__4_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__4_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_0__1__5_right_grid_pin_52_[0]),
		.ccff_head(grid_io_left_5_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_5_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_5_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_5_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_5_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_5_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_5_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_5_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_5_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_5_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_5_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_5_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_5_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_5_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_5_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_5_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_5_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_5_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_5_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_5_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_5_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_5_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_5_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_5_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_5_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_5_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_5_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_5_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_5_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_5_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_5_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_5_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_5_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_5_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_5_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_5_ccff_tail[0]));

	grid_clb grid_clb_1__7_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_6_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_149_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__6_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__6_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__6_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__6_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__6_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__6_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__6_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__6_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__6_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__6_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__6_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__6_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__6_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__6_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__6_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__6_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__5_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__5_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__5_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__5_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__5_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__5_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__5_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__5_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__5_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__5_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__5_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__5_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__5_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__5_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__5_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__5_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_0__1__6_right_grid_pin_52_[0]),
		.ccff_head(grid_io_left_6_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_6_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_6_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_6_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_6_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_6_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_6_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_6_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_6_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_6_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_6_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_6_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_6_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_6_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_6_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_6_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_6_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_6_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_6_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_6_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_6_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_6_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_6_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_6_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_6_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_6_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_6_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_6_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_6_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_6_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_6_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_6_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_6_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_6_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_6_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_6_ccff_tail[0]));

	grid_clb grid_clb_1__8_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_7_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_150_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__7_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__7_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__7_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__7_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__7_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__7_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__7_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__7_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__7_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__7_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__7_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__7_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__7_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__7_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__7_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__7_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__6_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__6_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__6_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__6_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__6_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__6_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__6_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__6_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__6_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__6_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__6_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__6_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__6_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__6_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__6_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__6_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_0__1__7_right_grid_pin_52_[0]),
		.ccff_head(grid_io_left_7_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_7_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_7_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_7_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_7_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_7_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_7_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_7_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_7_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_7_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_7_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_7_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_7_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_7_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_7_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_7_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_7_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_7_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_7_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_7_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_7_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_7_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_7_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_7_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_7_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_7_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_7_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_7_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_7_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_7_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_7_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_7_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_7_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_7_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_7_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_7_ccff_tail[0]));

	grid_clb grid_clb_1__9_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_8_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_151_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__8_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__8_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__8_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__8_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__8_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__8_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__8_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__8_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__8_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__8_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__8_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__8_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__8_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__8_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__8_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__8_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__7_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__7_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__7_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__7_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__7_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__7_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__7_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__7_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__7_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__7_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__7_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__7_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__7_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__7_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__7_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__7_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_0__1__8_right_grid_pin_52_[0]),
		.ccff_head(grid_io_left_8_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_8_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_8_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_8_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_8_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_8_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_8_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_8_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_8_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_8_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_8_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_8_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_8_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_8_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_8_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_8_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_8_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_8_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_8_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_8_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_8_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_8_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_8_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_8_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_8_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_8_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_8_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_8_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_8_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_8_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_8_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_8_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_8_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_8_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_8_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_8_ccff_tail[0]));

	grid_clb grid_clb_1__10_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_9_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_152_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__9_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__9_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__9_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__9_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__9_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__9_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__9_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__9_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__9_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__9_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__9_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__9_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__9_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__9_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__9_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__9_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__8_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__8_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__8_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__8_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__8_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__8_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__8_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__8_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__8_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__8_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__8_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__8_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__8_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__8_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__8_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__8_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_0__1__9_right_grid_pin_52_[0]),
		.ccff_head(grid_io_left_9_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_9_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_9_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_9_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_9_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_9_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_9_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_9_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_9_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_9_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_9_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_9_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_9_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_9_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_9_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_9_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_9_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_9_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_9_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_9_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_9_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_9_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_9_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_9_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_9_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_9_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_9_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_9_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_9_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_9_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_9_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_9_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_9_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_9_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_9_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_9_ccff_tail[0]));

	grid_clb grid_clb_1__11_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_10_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_153_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__10_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__10_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__10_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__10_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__10_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__10_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__10_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__10_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__10_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__10_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__10_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__10_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__10_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__10_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__10_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__10_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__9_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__9_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__9_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__9_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__9_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__9_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__9_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__9_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__9_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__9_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__9_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__9_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__9_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__9_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__9_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__9_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_0__1__10_right_grid_pin_52_[0]),
		.ccff_head(grid_io_left_10_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_10_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_10_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_10_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_10_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_10_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_10_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_10_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_10_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_10_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_10_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_10_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_10_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_10_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_10_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_10_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_10_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_10_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_10_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_10_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_10_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_10_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_10_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_10_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_10_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_10_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_10_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_10_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_10_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_10_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_10_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_10_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_10_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_10_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_10_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_10_ccff_tail[0]));

	grid_clb grid_clb_1__12_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(grid_clb_1__12__undriven_top_width_0_height_0__pin_32_[0]),
		.top_width_0_height_0__pin_33_(grid_clb_1__12__undriven_top_width_0_height_0__pin_33_[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__11_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__11_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__11_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__11_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__11_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__11_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__11_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__11_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__11_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__11_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__11_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__11_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__11_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__11_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__11_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__11_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__10_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__10_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__10_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__10_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__10_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__10_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__10_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__10_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__10_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__10_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__10_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__10_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__10_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__10_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__10_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__10_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_0__1__11_right_grid_pin_52_[0]),
		.ccff_head(grid_io_left_11_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_11_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_11_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_11_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_11_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_11_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_11_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_11_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_11_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_11_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_11_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_11_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_11_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_11_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_11_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_11_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_11_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_11_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_11_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_11_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_11_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_11_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_11_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_11_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_11_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_11_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_11_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_11_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_11_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_11_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_11_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_11_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_11_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_11_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_11_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_11_ccff_tail[0]));

	grid_clb grid_clb_2__1_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_11_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_154_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__12_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__12_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__12_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__12_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__12_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__12_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__12_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__12_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__12_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__12_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__12_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__12_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__12_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__12_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__12_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__12_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__0__1_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__0__1_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__0__1_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__0__1_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__0__1_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__0__1_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__0__1_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__0__1_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__0__1_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__0__1_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__0__1_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__0__1_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__0__1_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__0__1_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__0__1_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__0__1_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__0_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__0_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_12_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_12_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_12_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_12_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_12_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_12_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_12_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_12_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_12_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_12_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_12_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_12_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_12_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_12_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_12_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_12_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_12_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_12_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_12_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_12_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_12_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_12_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_12_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_12_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_12_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_12_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_12_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_12_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_12_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_12_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_12_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_12_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_12_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_12_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_12_ccff_tail[0]));

	grid_clb grid_clb_2__2_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_12_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_155_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__13_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__13_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__13_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__13_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__13_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__13_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__13_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__13_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__13_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__13_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__13_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__13_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__13_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__13_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__13_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__13_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__11_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__11_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__11_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__11_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__11_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__11_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__11_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__11_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__11_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__11_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__11_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__11_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__11_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__11_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__11_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__11_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__1_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__1_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_13_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_13_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_13_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_13_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_13_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_13_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_13_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_13_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_13_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_13_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_13_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_13_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_13_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_13_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_13_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_13_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_13_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_13_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_13_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_13_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_13_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_13_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_13_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_13_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_13_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_13_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_13_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_13_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_13_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_13_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_13_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_13_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_13_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_13_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_13_ccff_tail[0]));

	grid_clb grid_clb_2__3_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_13_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_156_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__14_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__14_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__14_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__14_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__14_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__14_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__14_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__14_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__14_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__14_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__14_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__14_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__14_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__14_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__14_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__14_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__12_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__12_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__12_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__12_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__12_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__12_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__12_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__12_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__12_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__12_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__12_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__12_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__12_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__12_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__12_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__12_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__2_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__2_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_14_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_14_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_14_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_14_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_14_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_14_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_14_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_14_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_14_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_14_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_14_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_14_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_14_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_14_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_14_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_14_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_14_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_14_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_14_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_14_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_14_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_14_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_14_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_14_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_14_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_14_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_14_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_14_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_14_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_14_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_14_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_14_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_14_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_14_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_14_ccff_tail[0]));

	grid_clb grid_clb_2__4_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_14_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_157_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__15_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__15_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__15_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__15_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__15_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__15_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__15_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__15_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__15_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__15_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__15_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__15_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__15_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__15_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__15_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__15_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__13_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__13_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__13_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__13_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__13_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__13_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__13_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__13_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__13_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__13_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__13_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__13_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__13_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__13_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__13_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__13_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__3_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__3_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_15_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_15_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_15_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_15_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_15_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_15_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_15_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_15_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_15_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_15_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_15_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_15_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_15_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_15_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_15_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_15_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_15_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_15_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_15_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_15_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_15_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_15_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_15_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_15_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_15_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_15_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_15_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_15_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_15_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_15_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_15_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_15_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_15_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_15_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_15_ccff_tail[0]));

	grid_clb grid_clb_2__5_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_15_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_158_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__16_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__16_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__16_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__16_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__16_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__16_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__16_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__16_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__16_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__16_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__16_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__16_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__16_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__16_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__16_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__16_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__14_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__14_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__14_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__14_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__14_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__14_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__14_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__14_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__14_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__14_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__14_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__14_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__14_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__14_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__14_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__14_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__4_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__4_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_16_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_16_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_16_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_16_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_16_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_16_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_16_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_16_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_16_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_16_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_16_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_16_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_16_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_16_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_16_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_16_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_16_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_16_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_16_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_16_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_16_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_16_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_16_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_16_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_16_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_16_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_16_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_16_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_16_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_16_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_16_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_16_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_16_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_16_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_16_ccff_tail[0]));

	grid_clb grid_clb_2__6_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_16_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_159_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__17_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__17_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__17_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__17_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__17_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__17_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__17_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__17_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__17_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__17_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__17_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__17_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__17_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__17_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__17_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__17_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__15_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__15_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__15_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__15_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__15_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__15_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__15_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__15_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__15_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__15_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__15_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__15_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__15_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__15_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__15_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__15_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__5_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__5_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_17_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_17_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_17_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_17_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_17_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_17_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_17_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_17_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_17_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_17_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_17_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_17_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_17_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_17_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_17_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_17_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_17_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_17_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_17_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_17_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_17_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_17_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_17_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_17_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_17_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_17_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_17_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_17_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_17_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_17_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_17_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_17_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_17_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_17_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_17_ccff_tail[0]));

	grid_clb grid_clb_2__7_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_17_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_160_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__18_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__18_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__18_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__18_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__18_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__18_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__18_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__18_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__18_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__18_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__18_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__18_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__18_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__18_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__18_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__18_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__16_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__16_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__16_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__16_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__16_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__16_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__16_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__16_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__16_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__16_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__16_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__16_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__16_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__16_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__16_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__16_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__6_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__6_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_18_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_18_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_18_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_18_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_18_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_18_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_18_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_18_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_18_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_18_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_18_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_18_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_18_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_18_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_18_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_18_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_18_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_18_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_18_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_18_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_18_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_18_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_18_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_18_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_18_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_18_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_18_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_18_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_18_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_18_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_18_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_18_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_18_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_18_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_18_ccff_tail[0]));

	grid_clb grid_clb_2__8_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_18_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_161_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__19_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__19_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__19_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__19_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__19_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__19_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__19_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__19_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__19_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__19_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__19_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__19_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__19_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__19_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__19_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__19_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__17_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__17_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__17_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__17_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__17_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__17_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__17_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__17_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__17_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__17_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__17_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__17_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__17_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__17_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__17_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__17_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__7_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__7_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_19_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_19_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_19_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_19_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_19_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_19_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_19_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_19_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_19_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_19_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_19_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_19_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_19_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_19_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_19_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_19_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_19_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_19_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_19_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_19_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_19_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_19_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_19_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_19_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_19_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_19_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_19_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_19_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_19_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_19_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_19_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_19_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_19_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_19_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_19_ccff_tail[0]));

	grid_clb grid_clb_2__9_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_19_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_162_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__20_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__20_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__20_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__20_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__20_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__20_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__20_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__20_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__20_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__20_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__20_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__20_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__20_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__20_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__20_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__20_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__18_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__18_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__18_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__18_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__18_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__18_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__18_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__18_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__18_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__18_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__18_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__18_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__18_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__18_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__18_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__18_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__8_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__8_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_20_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_20_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_20_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_20_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_20_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_20_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_20_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_20_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_20_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_20_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_20_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_20_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_20_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_20_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_20_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_20_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_20_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_20_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_20_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_20_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_20_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_20_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_20_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_20_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_20_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_20_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_20_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_20_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_20_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_20_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_20_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_20_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_20_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_20_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_20_ccff_tail[0]));

	grid_clb grid_clb_2__10_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_20_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_163_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__21_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__21_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__21_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__21_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__21_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__21_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__21_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__21_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__21_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__21_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__21_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__21_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__21_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__21_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__21_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__21_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__19_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__19_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__19_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__19_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__19_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__19_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__19_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__19_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__19_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__19_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__19_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__19_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__19_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__19_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__19_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__19_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__9_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__9_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_21_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_21_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_21_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_21_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_21_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_21_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_21_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_21_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_21_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_21_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_21_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_21_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_21_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_21_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_21_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_21_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_21_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_21_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_21_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_21_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_21_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_21_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_21_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_21_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_21_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_21_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_21_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_21_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_21_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_21_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_21_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_21_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_21_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_21_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_21_ccff_tail[0]));

	grid_clb grid_clb_2__11_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_21_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_164_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__22_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__22_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__22_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__22_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__22_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__22_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__22_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__22_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__22_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__22_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__22_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__22_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__22_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__22_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__22_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__22_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__20_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__20_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__20_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__20_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__20_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__20_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__20_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__20_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__20_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__20_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__20_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__20_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__20_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__20_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__20_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__20_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__10_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__10_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_22_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_22_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_22_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_22_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_22_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_22_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_22_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_22_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_22_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_22_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_22_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_22_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_22_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_22_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_22_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_22_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_22_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_22_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_22_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_22_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_22_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_22_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_22_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_22_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_22_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_22_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_22_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_22_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_22_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_22_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_22_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_22_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_22_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_22_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_22_ccff_tail[0]));

	grid_clb grid_clb_2__12_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_132_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_275_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__23_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__23_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__23_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__23_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__23_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__23_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__23_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__23_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__23_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__23_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__23_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__23_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__23_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__23_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__23_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__23_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__21_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__21_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__21_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__21_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__21_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__21_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__21_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__21_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__21_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__21_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__21_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__21_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__21_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__21_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__21_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__21_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__11_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__11_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_23_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_23_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_23_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_23_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_23_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_23_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_23_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_23_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_23_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_23_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_23_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_23_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_23_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_23_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_23_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_23_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_23_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_23_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_23_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_23_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_23_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_23_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_23_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_23_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_23_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_23_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_23_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_23_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_23_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_23_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_23_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_23_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_23_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_23_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_23_ccff_tail[0]));

	grid_clb grid_clb_3__1_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_22_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_165_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__24_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__24_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__24_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__24_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__24_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__24_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__24_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__24_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__24_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__24_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__24_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__24_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__24_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__24_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__24_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__24_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__0__2_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__0__2_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__0__2_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__0__2_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__0__2_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__0__2_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__0__2_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__0__2_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__0__2_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__0__2_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__0__2_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__0__2_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__0__2_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__0__2_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__0__2_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__0__2_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__12_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__12_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_24_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_24_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_24_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_24_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_24_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_24_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_24_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_24_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_24_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_24_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_24_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_24_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_24_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_24_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_24_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_24_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_24_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_24_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_24_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_24_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_24_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_24_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_24_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_24_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_24_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_24_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_24_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_24_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_24_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_24_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_24_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_24_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_24_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_24_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_24_ccff_tail[0]));

	grid_clb grid_clb_3__2_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_23_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_166_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__25_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__25_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__25_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__25_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__25_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__25_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__25_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__25_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__25_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__25_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__25_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__25_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__25_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__25_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__25_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__25_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__22_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__22_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__22_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__22_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__22_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__22_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__22_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__22_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__22_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__22_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__22_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__22_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__22_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__22_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__22_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__22_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__13_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__13_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_25_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_25_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_25_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_25_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_25_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_25_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_25_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_25_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_25_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_25_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_25_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_25_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_25_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_25_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_25_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_25_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_25_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_25_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_25_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_25_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_25_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_25_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_25_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_25_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_25_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_25_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_25_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_25_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_25_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_25_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_25_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_25_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_25_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_25_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_25_ccff_tail[0]));

	grid_clb grid_clb_3__3_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_24_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_167_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__26_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__26_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__26_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__26_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__26_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__26_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__26_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__26_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__26_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__26_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__26_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__26_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__26_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__26_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__26_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__26_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__23_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__23_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__23_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__23_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__23_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__23_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__23_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__23_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__23_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__23_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__23_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__23_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__23_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__23_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__23_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__23_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__14_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__14_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_26_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_26_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_26_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_26_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_26_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_26_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_26_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_26_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_26_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_26_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_26_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_26_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_26_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_26_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_26_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_26_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_26_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_26_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_26_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_26_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_26_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_26_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_26_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_26_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_26_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_26_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_26_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_26_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_26_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_26_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_26_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_26_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_26_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_26_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_26_ccff_tail[0]));

	grid_clb grid_clb_3__4_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_25_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_168_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__27_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__27_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__27_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__27_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__27_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__27_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__27_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__27_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__27_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__27_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__27_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__27_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__27_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__27_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__27_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__27_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__24_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__24_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__24_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__24_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__24_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__24_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__24_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__24_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__24_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__24_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__24_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__24_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__24_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__24_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__24_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__24_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__15_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__15_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_27_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_27_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_27_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_27_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_27_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_27_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_27_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_27_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_27_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_27_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_27_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_27_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_27_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_27_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_27_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_27_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_27_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_27_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_27_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_27_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_27_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_27_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_27_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_27_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_27_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_27_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_27_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_27_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_27_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_27_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_27_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_27_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_27_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_27_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_27_ccff_tail[0]));

	grid_clb grid_clb_3__5_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_26_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_169_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__28_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__28_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__28_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__28_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__28_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__28_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__28_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__28_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__28_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__28_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__28_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__28_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__28_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__28_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__28_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__28_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__25_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__25_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__25_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__25_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__25_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__25_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__25_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__25_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__25_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__25_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__25_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__25_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__25_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__25_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__25_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__25_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__16_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__16_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_28_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_28_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_28_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_28_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_28_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_28_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_28_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_28_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_28_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_28_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_28_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_28_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_28_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_28_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_28_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_28_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_28_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_28_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_28_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_28_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_28_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_28_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_28_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_28_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_28_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_28_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_28_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_28_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_28_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_28_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_28_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_28_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_28_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_28_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_28_ccff_tail[0]));

	grid_clb grid_clb_3__6_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_27_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_170_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__29_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__29_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__29_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__29_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__29_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__29_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__29_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__29_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__29_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__29_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__29_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__29_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__29_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__29_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__29_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__29_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__26_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__26_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__26_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__26_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__26_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__26_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__26_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__26_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__26_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__26_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__26_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__26_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__26_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__26_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__26_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__26_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__17_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__17_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_29_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_29_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_29_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_29_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_29_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_29_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_29_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_29_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_29_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_29_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_29_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_29_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_29_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_29_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_29_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_29_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_29_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_29_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_29_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_29_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_29_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_29_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_29_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_29_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_29_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_29_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_29_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_29_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_29_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_29_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_29_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_29_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_29_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_29_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_29_ccff_tail[0]));

	grid_clb grid_clb_3__7_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_28_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_171_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__30_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__30_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__30_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__30_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__30_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__30_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__30_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__30_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__30_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__30_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__30_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__30_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__30_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__30_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__30_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__30_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__27_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__27_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__27_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__27_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__27_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__27_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__27_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__27_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__27_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__27_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__27_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__27_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__27_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__27_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__27_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__27_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__18_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__18_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_30_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_30_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_30_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_30_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_30_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_30_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_30_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_30_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_30_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_30_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_30_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_30_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_30_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_30_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_30_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_30_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_30_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_30_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_30_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_30_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_30_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_30_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_30_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_30_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_30_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_30_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_30_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_30_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_30_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_30_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_30_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_30_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_30_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_30_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_30_ccff_tail[0]));

	grid_clb grid_clb_3__8_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_29_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_172_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__31_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__31_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__31_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__31_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__31_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__31_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__31_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__31_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__31_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__31_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__31_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__31_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__31_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__31_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__31_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__31_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__28_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__28_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__28_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__28_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__28_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__28_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__28_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__28_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__28_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__28_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__28_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__28_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__28_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__28_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__28_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__28_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__19_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__19_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_31_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_31_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_31_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_31_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_31_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_31_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_31_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_31_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_31_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_31_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_31_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_31_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_31_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_31_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_31_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_31_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_31_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_31_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_31_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_31_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_31_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_31_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_31_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_31_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_31_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_31_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_31_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_31_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_31_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_31_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_31_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_31_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_31_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_31_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_31_ccff_tail[0]));

	grid_clb grid_clb_3__9_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_30_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_173_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__32_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__32_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__32_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__32_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__32_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__32_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__32_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__32_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__32_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__32_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__32_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__32_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__32_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__32_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__32_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__32_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__29_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__29_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__29_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__29_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__29_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__29_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__29_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__29_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__29_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__29_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__29_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__29_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__29_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__29_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__29_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__29_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__20_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__20_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_32_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_32_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_32_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_32_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_32_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_32_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_32_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_32_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_32_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_32_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_32_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_32_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_32_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_32_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_32_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_32_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_32_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_32_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_32_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_32_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_32_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_32_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_32_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_32_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_32_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_32_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_32_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_32_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_32_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_32_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_32_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_32_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_32_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_32_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_32_ccff_tail[0]));

	grid_clb grid_clb_3__10_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_31_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_174_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__33_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__33_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__33_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__33_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__33_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__33_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__33_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__33_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__33_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__33_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__33_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__33_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__33_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__33_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__33_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__33_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__30_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__30_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__30_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__30_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__30_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__30_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__30_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__30_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__30_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__30_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__30_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__30_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__30_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__30_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__30_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__30_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__21_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__21_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_33_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_33_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_33_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_33_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_33_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_33_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_33_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_33_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_33_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_33_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_33_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_33_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_33_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_33_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_33_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_33_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_33_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_33_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_33_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_33_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_33_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_33_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_33_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_33_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_33_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_33_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_33_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_33_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_33_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_33_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_33_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_33_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_33_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_33_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_33_ccff_tail[0]));

	grid_clb grid_clb_3__11_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_32_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_175_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__34_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__34_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__34_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__34_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__34_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__34_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__34_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__34_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__34_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__34_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__34_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__34_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__34_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__34_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__34_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__34_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__31_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__31_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__31_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__31_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__31_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__31_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__31_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__31_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__31_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__31_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__31_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__31_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__31_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__31_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__31_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__31_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__22_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__22_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_34_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_34_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_34_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_34_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_34_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_34_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_34_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_34_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_34_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_34_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_34_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_34_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_34_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_34_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_34_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_34_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_34_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_34_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_34_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_34_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_34_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_34_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_34_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_34_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_34_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_34_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_34_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_34_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_34_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_34_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_34_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_34_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_34_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_34_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_34_ccff_tail[0]));

	grid_clb grid_clb_3__12_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_133_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_276_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__35_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__35_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__35_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__35_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__35_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__35_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__35_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__35_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__35_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__35_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__35_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__35_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__35_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__35_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__35_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__35_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__32_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__32_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__32_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__32_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__32_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__32_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__32_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__32_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__32_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__32_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__32_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__32_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__32_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__32_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__32_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__32_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__23_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__23_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_35_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_35_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_35_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_35_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_35_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_35_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_35_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_35_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_35_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_35_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_35_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_35_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_35_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_35_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_35_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_35_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_35_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_35_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_35_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_35_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_35_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_35_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_35_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_35_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_35_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_35_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_35_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_35_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_35_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_35_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_35_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_35_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_35_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_35_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_35_ccff_tail[0]));

	grid_clb grid_clb_4__1_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_33_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_176_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__36_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__36_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__36_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__36_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__36_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__36_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__36_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__36_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__36_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__36_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__36_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__36_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__36_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__36_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__36_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__36_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__0__3_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__0__3_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__0__3_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__0__3_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__0__3_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__0__3_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__0__3_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__0__3_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__0__3_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__0__3_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__0__3_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__0__3_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__0__3_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__0__3_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__0__3_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__0__3_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__24_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__24_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_36_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_36_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_36_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_36_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_36_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_36_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_36_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_36_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_36_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_36_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_36_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_36_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_36_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_36_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_36_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_36_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_36_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_36_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_36_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_36_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_36_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_36_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_36_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_36_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_36_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_36_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_36_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_36_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_36_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_36_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_36_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_36_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_36_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_36_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_36_ccff_tail[0]));

	grid_clb grid_clb_4__2_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_34_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_177_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__37_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__37_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__37_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__37_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__37_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__37_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__37_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__37_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__37_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__37_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__37_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__37_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__37_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__37_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__37_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__37_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__33_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__33_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__33_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__33_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__33_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__33_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__33_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__33_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__33_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__33_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__33_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__33_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__33_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__33_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__33_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__33_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__25_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__25_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_37_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_37_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_37_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_37_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_37_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_37_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_37_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_37_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_37_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_37_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_37_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_37_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_37_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_37_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_37_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_37_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_37_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_37_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_37_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_37_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_37_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_37_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_37_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_37_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_37_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_37_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_37_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_37_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_37_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_37_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_37_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_37_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_37_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_37_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_37_ccff_tail[0]));

	grid_clb grid_clb_4__3_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_35_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_178_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__38_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__38_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__38_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__38_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__38_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__38_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__38_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__38_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__38_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__38_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__38_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__38_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__38_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__38_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__38_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__38_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__34_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__34_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__34_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__34_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__34_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__34_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__34_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__34_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__34_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__34_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__34_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__34_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__34_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__34_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__34_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__34_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__26_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__26_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_38_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_38_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_38_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_38_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_38_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_38_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_38_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_38_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_38_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_38_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_38_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_38_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_38_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_38_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_38_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_38_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_38_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_38_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_38_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_38_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_38_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_38_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_38_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_38_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_38_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_38_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_38_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_38_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_38_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_38_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_38_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_38_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_38_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_38_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_38_ccff_tail[0]));

	grid_clb grid_clb_4__4_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_36_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_179_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__39_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__39_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__39_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__39_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__39_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__39_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__39_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__39_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__39_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__39_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__39_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__39_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__39_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__39_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__39_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__39_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__35_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__35_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__35_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__35_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__35_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__35_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__35_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__35_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__35_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__35_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__35_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__35_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__35_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__35_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__35_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__35_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__27_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__27_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_39_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_39_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_39_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_39_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_39_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_39_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_39_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_39_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_39_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_39_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_39_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_39_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_39_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_39_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_39_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_39_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_39_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_39_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_39_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_39_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_39_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_39_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_39_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_39_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_39_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_39_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_39_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_39_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_39_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_39_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_39_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_39_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_39_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_39_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_39_ccff_tail[0]));

	grid_clb grid_clb_4__5_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_37_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_180_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__40_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__40_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__40_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__40_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__40_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__40_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__40_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__40_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__40_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__40_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__40_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__40_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__40_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__40_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__40_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__40_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__36_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__36_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__36_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__36_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__36_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__36_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__36_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__36_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__36_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__36_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__36_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__36_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__36_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__36_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__36_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__36_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__28_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__28_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_40_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_40_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_40_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_40_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_40_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_40_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_40_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_40_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_40_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_40_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_40_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_40_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_40_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_40_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_40_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_40_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_40_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_40_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_40_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_40_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_40_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_40_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_40_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_40_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_40_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_40_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_40_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_40_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_40_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_40_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_40_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_40_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_40_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_40_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_40_ccff_tail[0]));

	grid_clb grid_clb_4__6_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_38_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_181_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__41_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__41_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__41_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__41_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__41_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__41_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__41_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__41_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__41_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__41_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__41_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__41_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__41_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__41_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__41_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__41_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__37_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__37_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__37_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__37_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__37_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__37_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__37_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__37_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__37_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__37_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__37_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__37_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__37_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__37_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__37_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__37_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__29_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__29_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_41_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_41_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_41_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_41_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_41_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_41_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_41_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_41_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_41_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_41_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_41_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_41_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_41_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_41_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_41_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_41_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_41_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_41_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_41_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_41_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_41_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_41_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_41_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_41_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_41_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_41_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_41_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_41_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_41_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_41_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_41_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_41_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_41_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_41_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_41_ccff_tail[0]));

	grid_clb grid_clb_4__7_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_39_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_182_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__42_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__42_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__42_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__42_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__42_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__42_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__42_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__42_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__42_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__42_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__42_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__42_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__42_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__42_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__42_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__42_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__38_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__38_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__38_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__38_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__38_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__38_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__38_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__38_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__38_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__38_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__38_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__38_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__38_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__38_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__38_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__38_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__30_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__30_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_42_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_42_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_42_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_42_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_42_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_42_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_42_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_42_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_42_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_42_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_42_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_42_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_42_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_42_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_42_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_42_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_42_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_42_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_42_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_42_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_42_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_42_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_42_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_42_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_42_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_42_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_42_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_42_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_42_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_42_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_42_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_42_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_42_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_42_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_42_ccff_tail[0]));

	grid_clb grid_clb_4__8_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_40_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_183_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__43_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__43_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__43_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__43_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__43_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__43_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__43_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__43_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__43_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__43_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__43_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__43_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__43_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__43_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__43_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__43_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__39_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__39_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__39_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__39_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__39_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__39_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__39_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__39_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__39_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__39_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__39_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__39_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__39_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__39_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__39_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__39_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__31_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__31_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_43_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_43_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_43_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_43_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_43_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_43_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_43_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_43_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_43_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_43_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_43_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_43_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_43_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_43_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_43_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_43_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_43_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_43_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_43_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_43_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_43_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_43_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_43_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_43_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_43_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_43_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_43_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_43_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_43_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_43_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_43_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_43_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_43_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_43_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_43_ccff_tail[0]));

	grid_clb grid_clb_4__9_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_41_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_184_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__44_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__44_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__44_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__44_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__44_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__44_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__44_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__44_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__44_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__44_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__44_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__44_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__44_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__44_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__44_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__44_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__40_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__40_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__40_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__40_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__40_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__40_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__40_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__40_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__40_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__40_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__40_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__40_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__40_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__40_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__40_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__40_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__32_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__32_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_44_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_44_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_44_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_44_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_44_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_44_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_44_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_44_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_44_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_44_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_44_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_44_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_44_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_44_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_44_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_44_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_44_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_44_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_44_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_44_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_44_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_44_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_44_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_44_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_44_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_44_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_44_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_44_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_44_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_44_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_44_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_44_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_44_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_44_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_44_ccff_tail[0]));

	grid_clb grid_clb_4__10_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_42_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_185_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__45_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__45_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__45_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__45_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__45_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__45_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__45_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__45_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__45_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__45_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__45_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__45_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__45_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__45_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__45_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__45_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__41_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__41_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__41_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__41_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__41_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__41_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__41_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__41_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__41_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__41_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__41_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__41_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__41_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__41_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__41_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__41_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__33_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__33_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_45_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_45_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_45_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_45_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_45_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_45_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_45_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_45_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_45_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_45_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_45_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_45_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_45_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_45_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_45_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_45_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_45_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_45_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_45_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_45_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_45_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_45_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_45_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_45_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_45_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_45_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_45_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_45_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_45_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_45_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_45_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_45_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_45_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_45_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_45_ccff_tail[0]));

	grid_clb grid_clb_4__11_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_43_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_186_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__46_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__46_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__46_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__46_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__46_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__46_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__46_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__46_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__46_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__46_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__46_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__46_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__46_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__46_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__46_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__46_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__42_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__42_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__42_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__42_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__42_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__42_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__42_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__42_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__42_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__42_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__42_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__42_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__42_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__42_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__42_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__42_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__34_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__34_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_46_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_46_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_46_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_46_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_46_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_46_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_46_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_46_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_46_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_46_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_46_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_46_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_46_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_46_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_46_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_46_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_46_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_46_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_46_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_46_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_46_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_46_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_46_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_46_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_46_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_46_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_46_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_46_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_46_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_46_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_46_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_46_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_46_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_46_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_46_ccff_tail[0]));

	grid_clb grid_clb_4__12_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_134_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_277_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__47_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__47_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__47_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__47_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__47_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__47_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__47_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__47_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__47_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__47_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__47_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__47_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__47_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__47_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__47_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__47_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__43_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__43_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__43_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__43_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__43_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__43_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__43_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__43_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__43_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__43_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__43_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__43_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__43_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__43_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__43_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__43_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__35_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__35_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_47_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_47_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_47_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_47_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_47_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_47_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_47_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_47_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_47_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_47_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_47_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_47_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_47_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_47_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_47_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_47_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_47_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_47_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_47_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_47_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_47_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_47_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_47_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_47_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_47_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_47_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_47_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_47_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_47_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_47_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_47_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_47_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_47_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_47_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_47_ccff_tail[0]));

	grid_clb grid_clb_5__1_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_44_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_187_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__48_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__48_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__48_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__48_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__48_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__48_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__48_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__48_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__48_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__48_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__48_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__48_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__48_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__48_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__48_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__48_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__0__4_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__0__4_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__0__4_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__0__4_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__0__4_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__0__4_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__0__4_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__0__4_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__0__4_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__0__4_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__0__4_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__0__4_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__0__4_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__0__4_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__0__4_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__0__4_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__36_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__36_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_48_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_48_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_48_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_48_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_48_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_48_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_48_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_48_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_48_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_48_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_48_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_48_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_48_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_48_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_48_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_48_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_48_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_48_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_48_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_48_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_48_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_48_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_48_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_48_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_48_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_48_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_48_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_48_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_48_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_48_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_48_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_48_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_48_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_48_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_48_ccff_tail[0]));

	grid_clb grid_clb_5__2_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_45_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_188_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__49_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__49_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__49_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__49_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__49_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__49_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__49_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__49_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__49_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__49_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__49_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__49_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__49_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__49_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__49_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__49_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__44_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__44_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__44_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__44_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__44_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__44_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__44_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__44_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__44_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__44_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__44_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__44_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__44_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__44_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__44_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__44_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__37_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__37_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_49_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_49_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_49_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_49_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_49_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_49_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_49_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_49_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_49_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_49_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_49_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_49_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_49_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_49_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_49_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_49_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_49_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_49_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_49_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_49_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_49_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_49_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_49_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_49_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_49_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_49_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_49_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_49_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_49_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_49_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_49_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_49_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_49_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_49_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_49_ccff_tail[0]));

	grid_clb grid_clb_5__3_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_46_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_189_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__50_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__50_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__50_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__50_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__50_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__50_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__50_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__50_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__50_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__50_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__50_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__50_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__50_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__50_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__50_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__50_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__45_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__45_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__45_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__45_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__45_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__45_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__45_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__45_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__45_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__45_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__45_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__45_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__45_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__45_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__45_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__45_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__38_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__38_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_50_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_50_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_50_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_50_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_50_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_50_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_50_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_50_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_50_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_50_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_50_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_50_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_50_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_50_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_50_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_50_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_50_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_50_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_50_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_50_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_50_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_50_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_50_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_50_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_50_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_50_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_50_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_50_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_50_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_50_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_50_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_50_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_50_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_50_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_50_ccff_tail[0]));

	grid_clb grid_clb_5__4_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_47_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_190_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__51_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__51_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__51_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__51_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__51_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__51_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__51_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__51_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__51_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__51_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__51_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__51_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__51_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__51_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__51_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__51_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__46_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__46_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__46_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__46_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__46_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__46_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__46_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__46_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__46_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__46_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__46_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__46_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__46_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__46_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__46_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__46_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__39_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__39_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_51_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_51_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_51_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_51_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_51_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_51_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_51_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_51_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_51_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_51_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_51_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_51_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_51_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_51_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_51_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_51_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_51_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_51_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_51_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_51_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_51_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_51_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_51_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_51_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_51_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_51_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_51_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_51_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_51_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_51_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_51_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_51_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_51_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_51_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_51_ccff_tail[0]));

	grid_clb grid_clb_5__5_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_48_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_191_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__52_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__52_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__52_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__52_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__52_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__52_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__52_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__52_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__52_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__52_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__52_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__52_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__52_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__52_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__52_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__52_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__47_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__47_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__47_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__47_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__47_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__47_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__47_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__47_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__47_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__47_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__47_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__47_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__47_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__47_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__47_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__47_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__40_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__40_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_52_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_52_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_52_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_52_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_52_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_52_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_52_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_52_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_52_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_52_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_52_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_52_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_52_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_52_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_52_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_52_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_52_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_52_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_52_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_52_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_52_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_52_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_52_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_52_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_52_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_52_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_52_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_52_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_52_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_52_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_52_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_52_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_52_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_52_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_52_ccff_tail[0]));

	grid_clb grid_clb_5__6_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_49_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_192_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__53_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__53_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__53_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__53_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__53_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__53_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__53_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__53_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__53_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__53_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__53_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__53_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__53_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__53_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__53_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__53_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__48_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__48_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__48_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__48_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__48_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__48_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__48_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__48_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__48_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__48_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__48_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__48_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__48_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__48_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__48_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__48_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__41_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__41_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_53_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_53_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_53_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_53_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_53_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_53_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_53_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_53_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_53_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_53_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_53_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_53_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_53_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_53_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_53_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_53_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_53_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_53_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_53_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_53_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_53_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_53_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_53_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_53_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_53_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_53_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_53_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_53_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_53_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_53_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_53_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_53_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_53_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_53_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_53_ccff_tail[0]));

	grid_clb grid_clb_5__7_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_50_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_193_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__54_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__54_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__54_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__54_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__54_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__54_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__54_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__54_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__54_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__54_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__54_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__54_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__54_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__54_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__54_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__54_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__49_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__49_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__49_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__49_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__49_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__49_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__49_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__49_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__49_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__49_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__49_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__49_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__49_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__49_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__49_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__49_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__42_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__42_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_54_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_54_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_54_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_54_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_54_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_54_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_54_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_54_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_54_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_54_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_54_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_54_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_54_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_54_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_54_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_54_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_54_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_54_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_54_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_54_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_54_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_54_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_54_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_54_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_54_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_54_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_54_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_54_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_54_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_54_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_54_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_54_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_54_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_54_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_54_ccff_tail[0]));

	grid_clb grid_clb_5__8_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_51_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_194_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__55_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__55_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__55_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__55_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__55_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__55_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__55_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__55_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__55_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__55_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__55_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__55_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__55_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__55_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__55_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__55_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__50_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__50_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__50_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__50_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__50_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__50_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__50_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__50_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__50_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__50_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__50_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__50_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__50_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__50_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__50_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__50_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__43_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__43_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_55_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_55_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_55_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_55_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_55_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_55_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_55_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_55_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_55_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_55_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_55_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_55_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_55_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_55_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_55_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_55_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_55_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_55_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_55_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_55_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_55_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_55_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_55_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_55_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_55_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_55_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_55_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_55_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_55_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_55_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_55_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_55_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_55_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_55_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_55_ccff_tail[0]));

	grid_clb grid_clb_5__9_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_52_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_195_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__56_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__56_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__56_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__56_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__56_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__56_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__56_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__56_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__56_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__56_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__56_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__56_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__56_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__56_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__56_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__56_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__51_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__51_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__51_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__51_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__51_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__51_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__51_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__51_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__51_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__51_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__51_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__51_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__51_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__51_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__51_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__51_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__44_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__44_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_56_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_56_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_56_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_56_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_56_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_56_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_56_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_56_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_56_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_56_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_56_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_56_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_56_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_56_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_56_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_56_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_56_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_56_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_56_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_56_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_56_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_56_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_56_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_56_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_56_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_56_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_56_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_56_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_56_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_56_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_56_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_56_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_56_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_56_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_56_ccff_tail[0]));

	grid_clb grid_clb_5__10_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_53_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_196_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__57_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__57_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__57_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__57_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__57_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__57_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__57_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__57_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__57_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__57_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__57_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__57_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__57_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__57_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__57_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__57_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__52_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__52_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__52_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__52_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__52_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__52_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__52_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__52_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__52_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__52_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__52_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__52_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__52_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__52_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__52_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__52_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__45_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__45_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_57_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_57_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_57_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_57_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_57_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_57_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_57_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_57_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_57_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_57_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_57_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_57_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_57_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_57_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_57_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_57_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_57_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_57_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_57_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_57_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_57_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_57_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_57_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_57_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_57_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_57_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_57_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_57_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_57_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_57_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_57_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_57_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_57_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_57_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_57_ccff_tail[0]));

	grid_clb grid_clb_5__11_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_54_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_197_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__58_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__58_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__58_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__58_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__58_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__58_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__58_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__58_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__58_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__58_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__58_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__58_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__58_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__58_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__58_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__58_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__53_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__53_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__53_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__53_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__53_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__53_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__53_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__53_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__53_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__53_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__53_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__53_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__53_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__53_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__53_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__53_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__46_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__46_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_58_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_58_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_58_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_58_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_58_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_58_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_58_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_58_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_58_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_58_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_58_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_58_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_58_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_58_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_58_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_58_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_58_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_58_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_58_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_58_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_58_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_58_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_58_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_58_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_58_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_58_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_58_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_58_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_58_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_58_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_58_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_58_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_58_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_58_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_58_ccff_tail[0]));

	grid_clb grid_clb_5__12_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_135_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_278_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__59_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__59_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__59_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__59_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__59_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__59_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__59_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__59_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__59_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__59_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__59_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__59_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__59_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__59_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__59_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__59_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__54_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__54_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__54_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__54_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__54_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__54_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__54_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__54_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__54_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__54_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__54_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__54_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__54_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__54_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__54_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__54_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__47_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__47_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_59_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_59_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_59_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_59_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_59_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_59_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_59_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_59_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_59_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_59_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_59_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_59_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_59_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_59_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_59_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_59_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_59_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_59_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_59_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_59_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_59_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_59_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_59_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_59_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_59_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_59_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_59_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_59_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_59_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_59_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_59_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_59_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_59_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_59_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_59_ccff_tail[0]));

	grid_clb grid_clb_6__1_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_55_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_198_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__60_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__60_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__60_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__60_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__60_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__60_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__60_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__60_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__60_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__60_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__60_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__60_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__60_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__60_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__60_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__60_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__0__5_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__0__5_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__0__5_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__0__5_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__0__5_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__0__5_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__0__5_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__0__5_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__0__5_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__0__5_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__0__5_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__0__5_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__0__5_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__0__5_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__0__5_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__0__5_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__48_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__48_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_60_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_60_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_60_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_60_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_60_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_60_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_60_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_60_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_60_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_60_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_60_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_60_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_60_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_60_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_60_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_60_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_60_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_60_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_60_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_60_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_60_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_60_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_60_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_60_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_60_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_60_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_60_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_60_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_60_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_60_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_60_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_60_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_60_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_60_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_60_ccff_tail[0]));

	grid_clb grid_clb_6__2_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_56_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_199_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__61_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__61_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__61_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__61_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__61_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__61_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__61_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__61_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__61_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__61_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__61_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__61_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__61_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__61_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__61_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__61_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__55_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__55_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__55_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__55_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__55_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__55_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__55_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__55_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__55_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__55_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__55_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__55_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__55_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__55_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__55_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__55_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__49_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__49_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_61_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_61_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_61_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_61_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_61_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_61_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_61_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_61_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_61_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_61_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_61_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_61_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_61_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_61_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_61_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_61_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_61_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_61_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_61_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_61_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_61_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_61_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_61_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_61_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_61_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_61_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_61_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_61_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_61_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_61_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_61_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_61_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_61_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_61_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_61_ccff_tail[0]));

	grid_clb grid_clb_6__3_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_57_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_200_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__62_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__62_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__62_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__62_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__62_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__62_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__62_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__62_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__62_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__62_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__62_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__62_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__62_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__62_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__62_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__62_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__56_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__56_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__56_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__56_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__56_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__56_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__56_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__56_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__56_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__56_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__56_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__56_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__56_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__56_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__56_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__56_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__50_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__50_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_62_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_62_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_62_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_62_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_62_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_62_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_62_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_62_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_62_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_62_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_62_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_62_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_62_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_62_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_62_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_62_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_62_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_62_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_62_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_62_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_62_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_62_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_62_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_62_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_62_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_62_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_62_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_62_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_62_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_62_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_62_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_62_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_62_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_62_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_62_ccff_tail[0]));

	grid_clb grid_clb_6__4_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_58_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_201_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__63_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__63_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__63_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__63_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__63_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__63_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__63_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__63_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__63_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__63_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__63_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__63_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__63_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__63_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__63_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__63_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__57_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__57_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__57_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__57_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__57_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__57_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__57_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__57_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__57_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__57_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__57_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__57_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__57_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__57_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__57_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__57_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__51_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__51_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_63_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_63_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_63_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_63_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_63_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_63_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_63_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_63_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_63_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_63_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_63_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_63_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_63_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_63_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_63_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_63_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_63_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_63_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_63_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_63_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_63_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_63_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_63_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_63_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_63_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_63_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_63_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_63_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_63_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_63_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_63_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_63_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_63_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_63_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_63_ccff_tail[0]));

	grid_clb grid_clb_6__5_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_59_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_202_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__64_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__64_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__64_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__64_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__64_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__64_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__64_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__64_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__64_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__64_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__64_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__64_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__64_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__64_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__64_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__64_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__58_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__58_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__58_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__58_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__58_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__58_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__58_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__58_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__58_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__58_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__58_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__58_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__58_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__58_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__58_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__58_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__52_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__52_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_64_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_64_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_64_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_64_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_64_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_64_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_64_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_64_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_64_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_64_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_64_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_64_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_64_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_64_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_64_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_64_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_64_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_64_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_64_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_64_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_64_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_64_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_64_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_64_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_64_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_64_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_64_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_64_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_64_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_64_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_64_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_64_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_64_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_64_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_64_ccff_tail[0]));

	grid_clb grid_clb_6__6_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_60_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_203_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__65_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__65_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__65_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__65_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__65_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__65_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__65_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__65_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__65_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__65_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__65_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__65_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__65_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__65_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__65_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__65_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__59_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__59_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__59_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__59_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__59_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__59_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__59_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__59_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__59_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__59_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__59_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__59_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__59_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__59_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__59_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__59_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__53_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__53_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_65_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_65_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_65_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_65_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_65_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_65_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_65_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_65_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_65_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_65_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_65_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_65_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_65_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_65_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_65_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_65_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_65_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_65_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_65_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_65_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_65_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_65_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_65_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_65_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_65_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_65_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_65_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_65_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_65_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_65_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_65_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_65_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_65_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_65_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_65_ccff_tail[0]));

	grid_clb grid_clb_6__7_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_61_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_204_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__66_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__66_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__66_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__66_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__66_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__66_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__66_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__66_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__66_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__66_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__66_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__66_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__66_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__66_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__66_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__66_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__60_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__60_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__60_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__60_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__60_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__60_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__60_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__60_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__60_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__60_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__60_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__60_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__60_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__60_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__60_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__60_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__54_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__54_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_66_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_66_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_66_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_66_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_66_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_66_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_66_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_66_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_66_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_66_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_66_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_66_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_66_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_66_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_66_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_66_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_66_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_66_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_66_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_66_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_66_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_66_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_66_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_66_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_66_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_66_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_66_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_66_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_66_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_66_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_66_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_66_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_66_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_66_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_66_ccff_tail[0]));

	grid_clb grid_clb_6__8_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_62_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_205_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__67_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__67_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__67_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__67_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__67_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__67_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__67_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__67_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__67_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__67_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__67_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__67_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__67_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__67_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__67_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__67_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__61_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__61_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__61_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__61_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__61_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__61_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__61_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__61_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__61_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__61_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__61_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__61_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__61_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__61_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__61_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__61_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__55_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__55_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_67_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_67_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_67_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_67_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_67_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_67_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_67_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_67_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_67_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_67_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_67_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_67_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_67_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_67_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_67_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_67_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_67_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_67_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_67_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_67_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_67_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_67_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_67_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_67_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_67_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_67_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_67_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_67_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_67_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_67_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_67_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_67_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_67_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_67_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_67_ccff_tail[0]));

	grid_clb grid_clb_6__9_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_63_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_206_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__68_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__68_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__68_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__68_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__68_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__68_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__68_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__68_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__68_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__68_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__68_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__68_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__68_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__68_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__68_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__68_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__62_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__62_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__62_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__62_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__62_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__62_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__62_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__62_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__62_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__62_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__62_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__62_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__62_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__62_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__62_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__62_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__56_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__56_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_68_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_68_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_68_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_68_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_68_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_68_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_68_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_68_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_68_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_68_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_68_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_68_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_68_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_68_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_68_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_68_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_68_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_68_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_68_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_68_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_68_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_68_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_68_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_68_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_68_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_68_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_68_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_68_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_68_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_68_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_68_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_68_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_68_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_68_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_68_ccff_tail[0]));

	grid_clb grid_clb_6__10_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_64_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_207_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__69_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__69_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__69_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__69_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__69_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__69_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__69_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__69_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__69_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__69_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__69_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__69_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__69_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__69_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__69_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__69_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__63_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__63_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__63_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__63_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__63_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__63_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__63_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__63_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__63_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__63_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__63_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__63_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__63_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__63_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__63_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__63_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__57_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__57_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_69_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_69_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_69_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_69_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_69_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_69_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_69_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_69_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_69_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_69_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_69_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_69_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_69_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_69_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_69_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_69_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_69_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_69_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_69_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_69_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_69_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_69_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_69_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_69_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_69_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_69_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_69_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_69_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_69_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_69_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_69_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_69_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_69_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_69_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_69_ccff_tail[0]));

	grid_clb grid_clb_6__11_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_65_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_208_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__70_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__70_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__70_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__70_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__70_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__70_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__70_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__70_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__70_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__70_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__70_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__70_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__70_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__70_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__70_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__70_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__64_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__64_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__64_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__64_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__64_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__64_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__64_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__64_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__64_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__64_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__64_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__64_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__64_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__64_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__64_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__64_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__58_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__58_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_70_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_70_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_70_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_70_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_70_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_70_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_70_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_70_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_70_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_70_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_70_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_70_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_70_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_70_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_70_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_70_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_70_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_70_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_70_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_70_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_70_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_70_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_70_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_70_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_70_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_70_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_70_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_70_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_70_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_70_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_70_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_70_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_70_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_70_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_70_ccff_tail[0]));

	grid_clb grid_clb_6__12_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_136_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_279_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__71_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__71_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__71_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__71_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__71_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__71_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__71_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__71_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__71_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__71_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__71_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__71_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__71_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__71_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__71_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__71_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__65_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__65_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__65_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__65_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__65_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__65_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__65_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__65_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__65_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__65_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__65_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__65_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__65_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__65_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__65_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__65_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__59_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__59_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_71_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_71_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_71_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_71_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_71_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_71_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_71_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_71_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_71_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_71_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_71_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_71_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_71_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_71_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_71_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_71_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_71_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_71_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_71_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_71_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_71_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_71_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_71_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_71_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_71_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_71_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_71_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_71_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_71_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_71_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_71_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_71_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_71_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_71_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_71_ccff_tail[0]));

	grid_clb grid_clb_7__1_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_66_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_209_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__72_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__72_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__72_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__72_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__72_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__72_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__72_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__72_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__72_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__72_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__72_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__72_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__72_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__72_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__72_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__72_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__0__6_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__0__6_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__0__6_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__0__6_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__0__6_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__0__6_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__0__6_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__0__6_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__0__6_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__0__6_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__0__6_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__0__6_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__0__6_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__0__6_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__0__6_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__0__6_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__60_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__60_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_72_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_72_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_72_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_72_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_72_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_72_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_72_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_72_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_72_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_72_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_72_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_72_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_72_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_72_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_72_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_72_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_72_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_72_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_72_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_72_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_72_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_72_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_72_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_72_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_72_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_72_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_72_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_72_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_72_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_72_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_72_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_72_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_72_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_72_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_72_ccff_tail[0]));

	grid_clb grid_clb_7__2_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_67_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_210_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__73_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__73_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__73_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__73_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__73_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__73_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__73_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__73_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__73_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__73_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__73_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__73_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__73_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__73_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__73_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__73_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__66_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__66_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__66_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__66_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__66_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__66_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__66_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__66_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__66_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__66_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__66_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__66_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__66_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__66_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__66_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__66_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__61_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__61_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_73_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_73_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_73_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_73_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_73_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_73_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_73_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_73_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_73_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_73_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_73_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_73_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_73_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_73_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_73_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_73_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_73_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_73_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_73_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_73_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_73_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_73_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_73_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_73_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_73_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_73_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_73_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_73_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_73_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_73_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_73_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_73_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_73_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_73_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_73_ccff_tail[0]));

	grid_clb grid_clb_7__3_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_68_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_211_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__74_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__74_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__74_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__74_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__74_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__74_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__74_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__74_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__74_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__74_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__74_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__74_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__74_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__74_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__74_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__74_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__67_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__67_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__67_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__67_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__67_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__67_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__67_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__67_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__67_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__67_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__67_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__67_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__67_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__67_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__67_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__67_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__62_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__62_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_74_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_74_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_74_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_74_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_74_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_74_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_74_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_74_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_74_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_74_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_74_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_74_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_74_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_74_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_74_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_74_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_74_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_74_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_74_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_74_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_74_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_74_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_74_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_74_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_74_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_74_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_74_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_74_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_74_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_74_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_74_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_74_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_74_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_74_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_74_ccff_tail[0]));

	grid_clb grid_clb_7__4_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_69_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_212_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__75_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__75_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__75_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__75_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__75_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__75_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__75_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__75_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__75_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__75_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__75_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__75_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__75_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__75_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__75_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__75_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__68_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__68_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__68_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__68_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__68_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__68_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__68_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__68_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__68_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__68_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__68_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__68_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__68_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__68_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__68_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__68_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__63_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__63_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_75_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_75_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_75_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_75_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_75_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_75_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_75_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_75_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_75_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_75_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_75_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_75_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_75_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_75_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_75_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_75_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_75_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_75_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_75_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_75_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_75_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_75_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_75_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_75_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_75_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_75_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_75_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_75_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_75_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_75_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_75_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_75_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_75_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_75_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_75_ccff_tail[0]));

	grid_clb grid_clb_7__5_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_70_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_213_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__76_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__76_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__76_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__76_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__76_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__76_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__76_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__76_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__76_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__76_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__76_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__76_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__76_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__76_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__76_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__76_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__69_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__69_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__69_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__69_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__69_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__69_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__69_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__69_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__69_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__69_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__69_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__69_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__69_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__69_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__69_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__69_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__64_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__64_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_76_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_76_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_76_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_76_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_76_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_76_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_76_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_76_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_76_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_76_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_76_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_76_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_76_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_76_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_76_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_76_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_76_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_76_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_76_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_76_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_76_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_76_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_76_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_76_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_76_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_76_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_76_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_76_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_76_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_76_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_76_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_76_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_76_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_76_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_76_ccff_tail[0]));

	grid_clb grid_clb_7__6_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_71_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_214_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__77_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__77_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__77_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__77_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__77_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__77_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__77_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__77_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__77_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__77_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__77_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__77_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__77_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__77_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__77_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__77_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__70_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__70_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__70_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__70_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__70_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__70_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__70_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__70_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__70_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__70_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__70_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__70_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__70_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__70_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__70_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__70_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__65_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__65_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_77_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_77_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_77_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_77_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_77_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_77_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_77_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_77_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_77_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_77_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_77_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_77_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_77_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_77_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_77_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_77_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_77_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_77_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_77_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_77_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_77_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_77_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_77_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_77_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_77_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_77_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_77_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_77_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_77_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_77_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_77_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_77_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_77_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_77_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_77_ccff_tail[0]));

	grid_clb grid_clb_7__7_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_72_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_215_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__78_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__78_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__78_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__78_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__78_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__78_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__78_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__78_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__78_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__78_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__78_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__78_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__78_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__78_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__78_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__78_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__71_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__71_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__71_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__71_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__71_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__71_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__71_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__71_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__71_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__71_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__71_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__71_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__71_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__71_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__71_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__71_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__66_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__66_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_78_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_78_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_78_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_78_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_78_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_78_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_78_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_78_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_78_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_78_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_78_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_78_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_78_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_78_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_78_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_78_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_78_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_78_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_78_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_78_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_78_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_78_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_78_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_78_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_78_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_78_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_78_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_78_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_78_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_78_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_78_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_78_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_78_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_78_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_78_ccff_tail[0]));

	grid_clb grid_clb_7__8_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_73_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_216_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__79_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__79_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__79_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__79_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__79_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__79_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__79_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__79_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__79_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__79_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__79_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__79_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__79_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__79_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__79_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__79_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__72_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__72_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__72_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__72_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__72_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__72_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__72_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__72_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__72_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__72_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__72_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__72_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__72_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__72_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__72_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__72_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__67_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__67_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_79_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_79_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_79_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_79_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_79_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_79_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_79_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_79_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_79_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_79_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_79_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_79_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_79_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_79_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_79_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_79_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_79_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_79_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_79_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_79_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_79_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_79_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_79_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_79_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_79_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_79_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_79_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_79_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_79_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_79_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_79_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_79_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_79_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_79_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_79_ccff_tail[0]));

	grid_clb grid_clb_7__9_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_74_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_217_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__80_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__80_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__80_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__80_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__80_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__80_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__80_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__80_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__80_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__80_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__80_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__80_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__80_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__80_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__80_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__80_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__73_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__73_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__73_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__73_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__73_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__73_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__73_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__73_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__73_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__73_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__73_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__73_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__73_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__73_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__73_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__73_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__68_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__68_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_80_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_80_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_80_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_80_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_80_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_80_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_80_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_80_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_80_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_80_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_80_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_80_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_80_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_80_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_80_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_80_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_80_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_80_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_80_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_80_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_80_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_80_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_80_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_80_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_80_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_80_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_80_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_80_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_80_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_80_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_80_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_80_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_80_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_80_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_80_ccff_tail[0]));

	grid_clb grid_clb_7__10_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_75_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_218_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__81_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__81_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__81_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__81_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__81_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__81_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__81_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__81_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__81_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__81_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__81_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__81_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__81_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__81_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__81_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__81_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__74_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__74_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__74_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__74_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__74_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__74_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__74_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__74_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__74_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__74_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__74_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__74_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__74_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__74_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__74_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__74_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__69_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__69_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_81_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_81_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_81_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_81_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_81_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_81_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_81_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_81_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_81_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_81_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_81_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_81_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_81_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_81_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_81_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_81_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_81_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_81_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_81_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_81_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_81_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_81_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_81_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_81_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_81_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_81_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_81_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_81_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_81_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_81_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_81_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_81_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_81_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_81_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_81_ccff_tail[0]));

	grid_clb grid_clb_7__11_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_76_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_219_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__82_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__82_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__82_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__82_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__82_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__82_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__82_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__82_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__82_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__82_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__82_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__82_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__82_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__82_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__82_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__82_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__75_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__75_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__75_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__75_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__75_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__75_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__75_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__75_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__75_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__75_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__75_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__75_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__75_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__75_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__75_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__75_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__70_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__70_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_82_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_82_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_82_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_82_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_82_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_82_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_82_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_82_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_82_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_82_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_82_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_82_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_82_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_82_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_82_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_82_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_82_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_82_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_82_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_82_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_82_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_82_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_82_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_82_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_82_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_82_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_82_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_82_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_82_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_82_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_82_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_82_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_82_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_82_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_82_ccff_tail[0]));

	grid_clb grid_clb_7__12_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_137_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_280_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__83_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__83_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__83_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__83_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__83_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__83_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__83_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__83_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__83_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__83_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__83_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__83_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__83_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__83_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__83_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__83_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__76_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__76_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__76_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__76_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__76_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__76_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__76_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__76_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__76_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__76_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__76_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__76_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__76_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__76_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__76_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__76_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__71_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__71_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_83_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_83_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_83_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_83_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_83_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_83_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_83_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_83_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_83_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_83_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_83_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_83_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_83_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_83_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_83_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_83_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_83_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_83_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_83_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_83_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_83_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_83_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_83_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_83_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_83_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_83_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_83_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_83_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_83_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_83_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_83_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_83_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_83_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_83_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_83_ccff_tail[0]));

	grid_clb grid_clb_8__1_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_77_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_220_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__84_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__84_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__84_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__84_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__84_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__84_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__84_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__84_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__84_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__84_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__84_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__84_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__84_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__84_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__84_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__84_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__0__7_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__0__7_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__0__7_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__0__7_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__0__7_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__0__7_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__0__7_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__0__7_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__0__7_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__0__7_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__0__7_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__0__7_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__0__7_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__0__7_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__0__7_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__0__7_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__72_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__72_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_84_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_84_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_84_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_84_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_84_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_84_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_84_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_84_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_84_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_84_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_84_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_84_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_84_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_84_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_84_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_84_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_84_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_84_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_84_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_84_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_84_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_84_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_84_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_84_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_84_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_84_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_84_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_84_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_84_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_84_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_84_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_84_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_84_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_84_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_84_ccff_tail[0]));

	grid_clb grid_clb_8__2_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_78_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_221_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__85_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__85_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__85_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__85_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__85_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__85_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__85_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__85_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__85_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__85_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__85_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__85_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__85_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__85_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__85_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__85_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__77_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__77_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__77_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__77_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__77_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__77_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__77_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__77_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__77_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__77_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__77_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__77_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__77_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__77_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__77_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__77_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__73_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__73_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_85_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_85_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_85_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_85_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_85_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_85_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_85_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_85_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_85_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_85_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_85_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_85_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_85_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_85_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_85_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_85_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_85_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_85_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_85_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_85_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_85_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_85_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_85_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_85_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_85_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_85_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_85_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_85_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_85_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_85_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_85_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_85_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_85_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_85_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_85_ccff_tail[0]));

	grid_clb grid_clb_8__3_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_79_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_222_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__86_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__86_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__86_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__86_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__86_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__86_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__86_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__86_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__86_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__86_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__86_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__86_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__86_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__86_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__86_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__86_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__78_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__78_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__78_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__78_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__78_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__78_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__78_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__78_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__78_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__78_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__78_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__78_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__78_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__78_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__78_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__78_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__74_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__74_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_86_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_86_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_86_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_86_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_86_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_86_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_86_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_86_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_86_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_86_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_86_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_86_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_86_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_86_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_86_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_86_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_86_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_86_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_86_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_86_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_86_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_86_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_86_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_86_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_86_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_86_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_86_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_86_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_86_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_86_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_86_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_86_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_86_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_86_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_86_ccff_tail[0]));

	grid_clb grid_clb_8__4_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_80_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_223_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__87_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__87_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__87_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__87_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__87_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__87_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__87_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__87_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__87_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__87_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__87_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__87_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__87_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__87_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__87_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__87_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__79_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__79_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__79_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__79_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__79_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__79_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__79_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__79_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__79_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__79_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__79_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__79_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__79_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__79_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__79_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__79_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__75_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__75_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_87_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_87_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_87_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_87_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_87_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_87_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_87_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_87_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_87_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_87_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_87_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_87_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_87_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_87_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_87_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_87_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_87_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_87_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_87_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_87_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_87_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_87_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_87_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_87_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_87_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_87_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_87_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_87_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_87_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_87_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_87_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_87_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_87_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_87_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_87_ccff_tail[0]));

	grid_clb grid_clb_8__5_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_81_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_224_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__88_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__88_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__88_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__88_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__88_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__88_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__88_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__88_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__88_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__88_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__88_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__88_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__88_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__88_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__88_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__88_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__80_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__80_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__80_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__80_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__80_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__80_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__80_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__80_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__80_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__80_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__80_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__80_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__80_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__80_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__80_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__80_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__76_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__76_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_88_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_88_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_88_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_88_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_88_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_88_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_88_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_88_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_88_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_88_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_88_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_88_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_88_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_88_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_88_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_88_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_88_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_88_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_88_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_88_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_88_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_88_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_88_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_88_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_88_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_88_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_88_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_88_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_88_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_88_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_88_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_88_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_88_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_88_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_88_ccff_tail[0]));

	grid_clb grid_clb_8__6_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_82_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_225_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__89_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__89_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__89_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__89_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__89_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__89_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__89_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__89_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__89_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__89_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__89_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__89_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__89_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__89_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__89_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__89_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__81_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__81_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__81_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__81_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__81_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__81_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__81_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__81_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__81_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__81_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__81_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__81_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__81_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__81_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__81_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__81_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__77_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__77_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_89_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_89_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_89_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_89_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_89_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_89_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_89_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_89_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_89_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_89_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_89_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_89_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_89_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_89_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_89_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_89_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_89_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_89_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_89_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_89_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_89_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_89_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_89_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_89_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_89_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_89_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_89_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_89_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_89_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_89_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_89_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_89_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_89_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_89_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_89_ccff_tail[0]));

	grid_clb grid_clb_8__7_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_83_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_226_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__90_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__90_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__90_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__90_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__90_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__90_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__90_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__90_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__90_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__90_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__90_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__90_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__90_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__90_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__90_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__90_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__82_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__82_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__82_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__82_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__82_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__82_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__82_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__82_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__82_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__82_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__82_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__82_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__82_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__82_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__82_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__82_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__78_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__78_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_90_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_90_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_90_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_90_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_90_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_90_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_90_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_90_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_90_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_90_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_90_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_90_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_90_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_90_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_90_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_90_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_90_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_90_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_90_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_90_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_90_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_90_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_90_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_90_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_90_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_90_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_90_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_90_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_90_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_90_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_90_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_90_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_90_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_90_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_90_ccff_tail[0]));

	grid_clb grid_clb_8__8_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_84_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_227_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__91_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__91_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__91_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__91_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__91_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__91_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__91_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__91_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__91_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__91_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__91_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__91_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__91_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__91_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__91_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__91_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__83_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__83_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__83_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__83_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__83_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__83_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__83_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__83_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__83_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__83_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__83_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__83_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__83_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__83_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__83_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__83_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__79_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__79_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_91_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_91_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_91_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_91_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_91_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_91_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_91_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_91_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_91_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_91_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_91_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_91_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_91_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_91_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_91_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_91_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_91_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_91_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_91_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_91_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_91_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_91_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_91_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_91_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_91_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_91_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_91_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_91_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_91_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_91_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_91_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_91_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_91_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_91_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_91_ccff_tail[0]));

	grid_clb grid_clb_8__9_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_85_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_228_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__92_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__92_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__92_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__92_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__92_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__92_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__92_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__92_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__92_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__92_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__92_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__92_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__92_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__92_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__92_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__92_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__84_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__84_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__84_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__84_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__84_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__84_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__84_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__84_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__84_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__84_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__84_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__84_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__84_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__84_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__84_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__84_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__80_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__80_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_92_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_92_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_92_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_92_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_92_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_92_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_92_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_92_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_92_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_92_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_92_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_92_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_92_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_92_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_92_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_92_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_92_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_92_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_92_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_92_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_92_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_92_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_92_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_92_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_92_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_92_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_92_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_92_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_92_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_92_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_92_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_92_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_92_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_92_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_92_ccff_tail[0]));

	grid_clb grid_clb_8__10_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_86_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_229_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__93_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__93_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__93_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__93_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__93_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__93_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__93_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__93_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__93_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__93_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__93_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__93_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__93_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__93_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__93_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__93_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__85_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__85_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__85_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__85_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__85_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__85_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__85_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__85_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__85_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__85_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__85_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__85_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__85_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__85_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__85_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__85_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__81_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__81_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_93_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_93_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_93_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_93_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_93_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_93_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_93_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_93_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_93_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_93_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_93_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_93_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_93_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_93_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_93_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_93_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_93_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_93_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_93_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_93_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_93_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_93_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_93_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_93_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_93_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_93_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_93_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_93_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_93_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_93_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_93_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_93_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_93_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_93_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_93_ccff_tail[0]));

	grid_clb grid_clb_8__11_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_87_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_230_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__94_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__94_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__94_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__94_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__94_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__94_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__94_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__94_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__94_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__94_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__94_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__94_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__94_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__94_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__94_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__94_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__86_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__86_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__86_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__86_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__86_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__86_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__86_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__86_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__86_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__86_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__86_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__86_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__86_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__86_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__86_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__86_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__82_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__82_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_94_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_94_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_94_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_94_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_94_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_94_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_94_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_94_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_94_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_94_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_94_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_94_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_94_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_94_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_94_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_94_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_94_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_94_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_94_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_94_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_94_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_94_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_94_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_94_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_94_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_94_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_94_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_94_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_94_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_94_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_94_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_94_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_94_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_94_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_94_ccff_tail[0]));

	grid_clb grid_clb_8__12_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_138_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_281_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__95_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__95_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__95_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__95_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__95_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__95_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__95_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__95_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__95_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__95_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__95_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__95_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__95_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__95_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__95_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__95_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__87_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__87_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__87_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__87_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__87_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__87_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__87_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__87_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__87_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__87_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__87_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__87_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__87_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__87_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__87_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__87_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__83_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__83_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_95_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_95_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_95_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_95_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_95_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_95_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_95_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_95_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_95_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_95_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_95_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_95_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_95_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_95_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_95_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_95_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_95_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_95_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_95_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_95_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_95_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_95_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_95_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_95_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_95_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_95_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_95_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_95_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_95_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_95_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_95_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_95_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_95_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_95_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_95_ccff_tail[0]));

	grid_clb grid_clb_9__1_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_88_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_231_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__96_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__96_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__96_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__96_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__96_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__96_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__96_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__96_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__96_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__96_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__96_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__96_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__96_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__96_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__96_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__96_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__0__8_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__0__8_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__0__8_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__0__8_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__0__8_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__0__8_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__0__8_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__0__8_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__0__8_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__0__8_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__0__8_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__0__8_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__0__8_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__0__8_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__0__8_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__0__8_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__84_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__84_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_96_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_96_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_96_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_96_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_96_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_96_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_96_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_96_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_96_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_96_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_96_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_96_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_96_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_96_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_96_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_96_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_96_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_96_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_96_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_96_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_96_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_96_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_96_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_96_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_96_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_96_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_96_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_96_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_96_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_96_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_96_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_96_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_96_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_96_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_96_ccff_tail[0]));

	grid_clb grid_clb_9__2_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_89_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_232_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__97_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__97_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__97_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__97_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__97_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__97_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__97_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__97_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__97_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__97_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__97_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__97_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__97_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__97_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__97_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__97_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__88_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__88_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__88_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__88_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__88_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__88_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__88_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__88_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__88_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__88_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__88_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__88_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__88_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__88_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__88_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__88_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__85_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__85_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_97_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_97_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_97_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_97_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_97_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_97_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_97_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_97_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_97_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_97_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_97_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_97_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_97_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_97_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_97_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_97_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_97_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_97_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_97_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_97_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_97_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_97_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_97_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_97_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_97_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_97_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_97_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_97_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_97_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_97_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_97_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_97_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_97_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_97_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_97_ccff_tail[0]));

	grid_clb grid_clb_9__3_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_90_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_233_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__98_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__98_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__98_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__98_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__98_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__98_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__98_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__98_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__98_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__98_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__98_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__98_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__98_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__98_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__98_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__98_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__89_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__89_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__89_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__89_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__89_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__89_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__89_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__89_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__89_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__89_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__89_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__89_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__89_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__89_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__89_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__89_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__86_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__86_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_98_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_98_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_98_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_98_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_98_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_98_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_98_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_98_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_98_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_98_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_98_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_98_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_98_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_98_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_98_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_98_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_98_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_98_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_98_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_98_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_98_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_98_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_98_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_98_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_98_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_98_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_98_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_98_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_98_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_98_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_98_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_98_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_98_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_98_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_98_ccff_tail[0]));

	grid_clb grid_clb_9__4_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_91_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_234_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__99_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__99_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__99_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__99_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__99_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__99_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__99_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__99_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__99_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__99_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__99_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__99_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__99_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__99_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__99_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__99_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__90_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__90_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__90_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__90_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__90_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__90_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__90_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__90_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__90_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__90_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__90_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__90_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__90_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__90_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__90_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__90_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__87_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__87_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_99_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_99_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_99_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_99_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_99_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_99_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_99_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_99_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_99_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_99_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_99_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_99_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_99_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_99_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_99_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_99_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_99_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_99_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_99_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_99_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_99_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_99_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_99_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_99_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_99_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_99_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_99_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_99_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_99_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_99_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_99_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_99_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_99_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_99_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_99_ccff_tail[0]));

	grid_clb grid_clb_9__5_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_92_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_235_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__100_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__100_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__100_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__100_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__100_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__100_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__100_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__100_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__100_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__100_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__100_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__100_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__100_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__100_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__100_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__100_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__91_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__91_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__91_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__91_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__91_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__91_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__91_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__91_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__91_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__91_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__91_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__91_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__91_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__91_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__91_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__91_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__88_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__88_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_100_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_100_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_100_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_100_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_100_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_100_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_100_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_100_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_100_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_100_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_100_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_100_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_100_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_100_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_100_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_100_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_100_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_100_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_100_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_100_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_100_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_100_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_100_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_100_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_100_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_100_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_100_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_100_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_100_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_100_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_100_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_100_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_100_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_100_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_100_ccff_tail[0]));

	grid_clb grid_clb_9__6_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_93_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_236_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__101_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__101_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__101_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__101_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__101_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__101_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__101_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__101_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__101_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__101_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__101_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__101_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__101_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__101_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__101_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__101_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__92_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__92_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__92_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__92_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__92_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__92_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__92_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__92_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__92_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__92_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__92_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__92_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__92_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__92_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__92_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__92_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__89_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__89_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_101_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_101_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_101_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_101_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_101_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_101_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_101_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_101_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_101_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_101_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_101_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_101_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_101_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_101_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_101_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_101_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_101_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_101_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_101_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_101_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_101_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_101_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_101_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_101_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_101_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_101_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_101_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_101_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_101_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_101_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_101_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_101_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_101_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_101_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_101_ccff_tail[0]));

	grid_clb grid_clb_9__7_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_94_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_237_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__102_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__102_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__102_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__102_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__102_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__102_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__102_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__102_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__102_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__102_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__102_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__102_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__102_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__102_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__102_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__102_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__93_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__93_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__93_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__93_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__93_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__93_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__93_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__93_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__93_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__93_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__93_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__93_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__93_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__93_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__93_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__93_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__90_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__90_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_102_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_102_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_102_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_102_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_102_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_102_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_102_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_102_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_102_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_102_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_102_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_102_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_102_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_102_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_102_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_102_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_102_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_102_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_102_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_102_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_102_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_102_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_102_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_102_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_102_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_102_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_102_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_102_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_102_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_102_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_102_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_102_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_102_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_102_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_102_ccff_tail[0]));

	grid_clb grid_clb_9__8_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_95_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_238_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__103_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__103_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__103_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__103_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__103_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__103_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__103_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__103_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__103_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__103_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__103_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__103_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__103_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__103_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__103_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__103_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__94_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__94_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__94_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__94_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__94_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__94_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__94_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__94_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__94_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__94_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__94_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__94_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__94_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__94_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__94_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__94_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__91_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__91_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_103_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_103_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_103_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_103_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_103_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_103_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_103_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_103_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_103_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_103_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_103_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_103_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_103_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_103_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_103_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_103_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_103_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_103_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_103_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_103_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_103_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_103_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_103_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_103_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_103_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_103_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_103_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_103_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_103_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_103_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_103_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_103_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_103_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_103_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_103_ccff_tail[0]));

	grid_clb grid_clb_9__9_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_96_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_239_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__104_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__104_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__104_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__104_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__104_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__104_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__104_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__104_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__104_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__104_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__104_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__104_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__104_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__104_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__104_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__104_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__95_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__95_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__95_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__95_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__95_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__95_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__95_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__95_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__95_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__95_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__95_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__95_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__95_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__95_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__95_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__95_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__92_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__92_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_104_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_104_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_104_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_104_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_104_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_104_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_104_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_104_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_104_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_104_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_104_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_104_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_104_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_104_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_104_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_104_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_104_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_104_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_104_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_104_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_104_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_104_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_104_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_104_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_104_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_104_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_104_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_104_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_104_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_104_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_104_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_104_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_104_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_104_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_104_ccff_tail[0]));

	grid_clb grid_clb_9__10_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_97_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_240_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__105_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__105_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__105_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__105_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__105_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__105_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__105_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__105_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__105_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__105_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__105_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__105_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__105_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__105_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__105_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__105_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__96_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__96_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__96_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__96_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__96_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__96_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__96_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__96_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__96_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__96_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__96_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__96_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__96_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__96_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__96_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__96_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__93_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__93_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_105_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_105_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_105_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_105_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_105_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_105_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_105_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_105_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_105_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_105_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_105_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_105_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_105_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_105_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_105_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_105_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_105_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_105_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_105_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_105_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_105_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_105_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_105_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_105_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_105_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_105_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_105_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_105_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_105_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_105_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_105_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_105_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_105_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_105_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_105_ccff_tail[0]));

	grid_clb grid_clb_9__11_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_98_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_241_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__106_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__106_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__106_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__106_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__106_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__106_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__106_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__106_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__106_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__106_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__106_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__106_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__106_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__106_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__106_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__106_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__97_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__97_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__97_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__97_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__97_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__97_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__97_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__97_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__97_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__97_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__97_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__97_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__97_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__97_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__97_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__97_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__94_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__94_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_106_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_106_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_106_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_106_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_106_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_106_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_106_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_106_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_106_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_106_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_106_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_106_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_106_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_106_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_106_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_106_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_106_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_106_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_106_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_106_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_106_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_106_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_106_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_106_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_106_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_106_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_106_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_106_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_106_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_106_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_106_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_106_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_106_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_106_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_106_ccff_tail[0]));

	grid_clb grid_clb_9__12_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_139_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_282_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__107_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__107_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__107_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__107_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__107_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__107_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__107_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__107_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__107_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__107_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__107_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__107_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__107_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__107_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__107_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__107_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__98_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__98_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__98_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__98_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__98_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__98_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__98_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__98_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__98_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__98_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__98_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__98_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__98_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__98_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__98_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__98_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__95_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__95_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_107_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_107_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_107_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_107_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_107_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_107_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_107_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_107_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_107_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_107_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_107_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_107_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_107_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_107_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_107_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_107_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_107_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_107_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_107_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_107_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_107_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_107_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_107_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_107_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_107_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_107_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_107_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_107_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_107_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_107_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_107_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_107_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_107_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_107_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_107_ccff_tail[0]));

	grid_clb grid_clb_10__1_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_99_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_242_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__108_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__108_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__108_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__108_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__108_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__108_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__108_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__108_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__108_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__108_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__108_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__108_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__108_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__108_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__108_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__108_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__0__9_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__0__9_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__0__9_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__0__9_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__0__9_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__0__9_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__0__9_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__0__9_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__0__9_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__0__9_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__0__9_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__0__9_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__0__9_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__0__9_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__0__9_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__0__9_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__96_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__96_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_108_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_108_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_108_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_108_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_108_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_108_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_108_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_108_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_108_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_108_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_108_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_108_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_108_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_108_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_108_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_108_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_108_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_108_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_108_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_108_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_108_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_108_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_108_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_108_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_108_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_108_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_108_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_108_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_108_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_108_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_108_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_108_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_108_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_108_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_108_ccff_tail[0]));

	grid_clb grid_clb_10__2_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_100_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_243_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__109_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__109_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__109_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__109_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__109_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__109_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__109_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__109_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__109_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__109_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__109_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__109_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__109_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__109_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__109_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__109_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__99_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__99_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__99_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__99_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__99_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__99_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__99_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__99_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__99_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__99_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__99_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__99_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__99_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__99_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__99_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__99_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__97_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__97_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_109_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_109_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_109_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_109_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_109_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_109_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_109_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_109_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_109_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_109_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_109_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_109_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_109_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_109_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_109_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_109_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_109_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_109_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_109_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_109_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_109_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_109_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_109_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_109_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_109_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_109_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_109_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_109_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_109_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_109_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_109_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_109_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_109_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_109_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_109_ccff_tail[0]));

	grid_clb grid_clb_10__3_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_101_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_244_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__110_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__110_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__110_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__110_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__110_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__110_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__110_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__110_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__110_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__110_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__110_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__110_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__110_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__110_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__110_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__110_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__100_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__100_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__100_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__100_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__100_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__100_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__100_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__100_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__100_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__100_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__100_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__100_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__100_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__100_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__100_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__100_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__98_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__98_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_110_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_110_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_110_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_110_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_110_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_110_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_110_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_110_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_110_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_110_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_110_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_110_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_110_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_110_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_110_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_110_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_110_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_110_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_110_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_110_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_110_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_110_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_110_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_110_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_110_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_110_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_110_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_110_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_110_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_110_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_110_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_110_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_110_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_110_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_110_ccff_tail[0]));

	grid_clb grid_clb_10__4_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_102_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_245_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__111_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__111_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__111_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__111_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__111_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__111_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__111_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__111_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__111_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__111_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__111_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__111_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__111_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__111_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__111_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__111_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__101_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__101_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__101_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__101_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__101_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__101_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__101_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__101_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__101_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__101_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__101_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__101_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__101_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__101_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__101_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__101_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__99_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__99_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_111_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_111_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_111_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_111_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_111_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_111_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_111_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_111_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_111_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_111_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_111_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_111_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_111_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_111_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_111_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_111_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_111_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_111_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_111_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_111_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_111_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_111_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_111_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_111_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_111_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_111_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_111_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_111_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_111_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_111_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_111_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_111_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_111_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_111_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_111_ccff_tail[0]));

	grid_clb grid_clb_10__5_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_103_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_246_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__112_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__112_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__112_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__112_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__112_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__112_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__112_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__112_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__112_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__112_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__112_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__112_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__112_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__112_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__112_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__112_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__102_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__102_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__102_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__102_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__102_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__102_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__102_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__102_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__102_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__102_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__102_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__102_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__102_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__102_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__102_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__102_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__100_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__100_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_112_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_112_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_112_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_112_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_112_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_112_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_112_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_112_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_112_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_112_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_112_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_112_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_112_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_112_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_112_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_112_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_112_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_112_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_112_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_112_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_112_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_112_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_112_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_112_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_112_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_112_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_112_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_112_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_112_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_112_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_112_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_112_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_112_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_112_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_112_ccff_tail[0]));

	grid_clb grid_clb_10__6_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_104_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_247_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__113_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__113_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__113_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__113_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__113_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__113_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__113_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__113_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__113_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__113_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__113_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__113_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__113_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__113_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__113_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__113_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__103_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__103_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__103_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__103_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__103_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__103_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__103_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__103_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__103_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__103_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__103_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__103_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__103_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__103_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__103_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__103_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__101_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__101_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_113_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_113_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_113_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_113_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_113_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_113_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_113_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_113_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_113_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_113_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_113_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_113_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_113_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_113_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_113_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_113_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_113_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_113_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_113_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_113_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_113_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_113_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_113_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_113_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_113_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_113_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_113_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_113_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_113_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_113_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_113_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_113_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_113_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_113_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_113_ccff_tail[0]));

	grid_clb grid_clb_10__7_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_105_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_248_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__114_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__114_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__114_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__114_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__114_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__114_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__114_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__114_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__114_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__114_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__114_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__114_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__114_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__114_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__114_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__114_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__104_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__104_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__104_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__104_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__104_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__104_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__104_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__104_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__104_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__104_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__104_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__104_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__104_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__104_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__104_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__104_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__102_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__102_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_114_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_114_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_114_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_114_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_114_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_114_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_114_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_114_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_114_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_114_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_114_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_114_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_114_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_114_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_114_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_114_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_114_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_114_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_114_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_114_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_114_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_114_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_114_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_114_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_114_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_114_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_114_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_114_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_114_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_114_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_114_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_114_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_114_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_114_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_114_ccff_tail[0]));

	grid_clb grid_clb_10__8_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_106_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_249_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__115_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__115_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__115_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__115_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__115_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__115_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__115_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__115_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__115_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__115_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__115_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__115_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__115_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__115_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__115_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__115_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__105_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__105_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__105_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__105_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__105_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__105_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__105_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__105_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__105_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__105_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__105_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__105_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__105_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__105_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__105_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__105_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__103_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__103_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_115_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_115_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_115_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_115_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_115_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_115_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_115_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_115_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_115_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_115_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_115_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_115_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_115_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_115_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_115_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_115_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_115_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_115_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_115_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_115_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_115_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_115_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_115_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_115_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_115_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_115_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_115_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_115_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_115_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_115_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_115_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_115_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_115_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_115_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_115_ccff_tail[0]));

	grid_clb grid_clb_10__9_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_107_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_250_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__116_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__116_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__116_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__116_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__116_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__116_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__116_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__116_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__116_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__116_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__116_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__116_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__116_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__116_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__116_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__116_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__106_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__106_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__106_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__106_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__106_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__106_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__106_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__106_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__106_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__106_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__106_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__106_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__106_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__106_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__106_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__106_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__104_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__104_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_116_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_116_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_116_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_116_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_116_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_116_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_116_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_116_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_116_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_116_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_116_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_116_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_116_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_116_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_116_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_116_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_116_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_116_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_116_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_116_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_116_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_116_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_116_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_116_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_116_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_116_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_116_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_116_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_116_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_116_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_116_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_116_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_116_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_116_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_116_ccff_tail[0]));

	grid_clb grid_clb_10__10_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_108_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_251_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__117_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__117_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__117_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__117_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__117_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__117_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__117_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__117_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__117_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__117_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__117_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__117_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__117_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__117_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__117_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__117_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__107_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__107_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__107_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__107_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__107_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__107_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__107_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__107_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__107_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__107_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__107_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__107_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__107_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__107_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__107_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__107_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__105_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__105_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_117_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_117_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_117_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_117_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_117_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_117_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_117_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_117_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_117_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_117_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_117_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_117_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_117_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_117_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_117_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_117_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_117_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_117_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_117_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_117_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_117_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_117_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_117_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_117_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_117_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_117_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_117_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_117_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_117_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_117_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_117_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_117_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_117_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_117_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_117_ccff_tail[0]));

	grid_clb grid_clb_10__11_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_109_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_252_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__118_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__118_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__118_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__118_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__118_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__118_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__118_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__118_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__118_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__118_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__118_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__118_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__118_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__118_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__118_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__118_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__108_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__108_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__108_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__108_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__108_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__108_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__108_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__108_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__108_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__108_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__108_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__108_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__108_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__108_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__108_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__108_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__106_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__106_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_118_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_118_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_118_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_118_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_118_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_118_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_118_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_118_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_118_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_118_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_118_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_118_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_118_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_118_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_118_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_118_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_118_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_118_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_118_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_118_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_118_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_118_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_118_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_118_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_118_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_118_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_118_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_118_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_118_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_118_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_118_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_118_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_118_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_118_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_118_ccff_tail[0]));

	grid_clb grid_clb_10__12_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_140_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_283_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__119_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__119_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__119_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__119_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__119_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__119_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__119_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__119_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__119_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__119_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__119_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__119_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__119_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__119_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__119_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__119_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__109_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__109_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__109_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__109_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__109_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__109_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__109_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__109_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__109_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__109_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__109_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__109_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__109_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__109_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__109_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__109_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__107_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__107_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_119_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_119_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_119_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_119_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_119_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_119_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_119_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_119_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_119_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_119_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_119_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_119_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_119_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_119_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_119_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_119_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_119_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_119_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_119_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_119_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_119_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_119_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_119_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_119_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_119_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_119_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_119_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_119_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_119_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_119_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_119_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_119_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_119_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_119_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_119_ccff_tail[0]));

	grid_clb grid_clb_11__1_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_110_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_253_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__120_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__120_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__120_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__120_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__120_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__120_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__120_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__120_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__120_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__120_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__120_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__120_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__120_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__120_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__120_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__120_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__0__10_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__0__10_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__0__10_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__0__10_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__0__10_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__0__10_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__0__10_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__0__10_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__0__10_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__0__10_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__0__10_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__0__10_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__0__10_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__0__10_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__0__10_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__0__10_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__108_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__108_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_120_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_120_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_120_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_120_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_120_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_120_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_120_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_120_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_120_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_120_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_120_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_120_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_120_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_120_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_120_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_120_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_120_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_120_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_120_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_120_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_120_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_120_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_120_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_120_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_120_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_120_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_120_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_120_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_120_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_120_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_120_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_120_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_120_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_120_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_120_ccff_tail[0]));

	grid_clb grid_clb_11__2_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_111_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_254_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__121_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__121_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__121_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__121_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__121_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__121_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__121_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__121_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__121_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__121_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__121_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__121_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__121_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__121_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__121_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__121_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__110_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__110_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__110_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__110_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__110_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__110_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__110_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__110_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__110_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__110_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__110_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__110_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__110_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__110_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__110_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__110_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__109_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__109_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_121_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_121_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_121_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_121_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_121_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_121_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_121_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_121_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_121_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_121_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_121_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_121_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_121_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_121_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_121_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_121_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_121_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_121_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_121_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_121_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_121_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_121_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_121_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_121_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_121_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_121_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_121_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_121_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_121_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_121_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_121_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_121_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_121_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_121_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_121_ccff_tail[0]));

	grid_clb grid_clb_11__3_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_112_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_255_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__122_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__122_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__122_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__122_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__122_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__122_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__122_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__122_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__122_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__122_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__122_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__122_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__122_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__122_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__122_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__122_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__111_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__111_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__111_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__111_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__111_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__111_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__111_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__111_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__111_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__111_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__111_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__111_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__111_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__111_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__111_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__111_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__110_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__110_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_122_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_122_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_122_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_122_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_122_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_122_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_122_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_122_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_122_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_122_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_122_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_122_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_122_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_122_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_122_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_122_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_122_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_122_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_122_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_122_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_122_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_122_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_122_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_122_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_122_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_122_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_122_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_122_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_122_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_122_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_122_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_122_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_122_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_122_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_122_ccff_tail[0]));

	grid_clb grid_clb_11__4_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_113_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_256_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__123_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__123_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__123_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__123_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__123_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__123_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__123_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__123_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__123_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__123_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__123_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__123_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__123_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__123_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__123_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__123_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__112_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__112_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__112_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__112_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__112_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__112_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__112_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__112_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__112_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__112_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__112_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__112_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__112_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__112_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__112_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__112_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__111_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__111_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_123_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_123_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_123_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_123_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_123_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_123_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_123_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_123_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_123_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_123_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_123_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_123_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_123_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_123_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_123_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_123_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_123_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_123_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_123_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_123_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_123_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_123_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_123_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_123_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_123_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_123_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_123_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_123_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_123_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_123_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_123_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_123_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_123_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_123_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_123_ccff_tail[0]));

	grid_clb grid_clb_11__5_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_114_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_257_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__124_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__124_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__124_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__124_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__124_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__124_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__124_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__124_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__124_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__124_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__124_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__124_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__124_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__124_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__124_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__124_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__113_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__113_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__113_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__113_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__113_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__113_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__113_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__113_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__113_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__113_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__113_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__113_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__113_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__113_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__113_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__113_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__112_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__112_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_124_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_124_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_124_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_124_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_124_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_124_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_124_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_124_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_124_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_124_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_124_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_124_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_124_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_124_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_124_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_124_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_124_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_124_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_124_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_124_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_124_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_124_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_124_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_124_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_124_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_124_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_124_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_124_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_124_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_124_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_124_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_124_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_124_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_124_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_124_ccff_tail[0]));

	grid_clb grid_clb_11__6_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_115_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_258_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__125_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__125_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__125_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__125_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__125_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__125_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__125_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__125_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__125_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__125_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__125_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__125_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__125_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__125_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__125_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__125_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__114_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__114_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__114_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__114_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__114_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__114_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__114_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__114_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__114_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__114_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__114_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__114_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__114_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__114_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__114_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__114_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__113_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__113_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_125_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_125_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_125_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_125_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_125_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_125_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_125_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_125_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_125_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_125_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_125_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_125_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_125_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_125_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_125_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_125_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_125_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_125_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_125_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_125_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_125_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_125_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_125_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_125_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_125_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_125_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_125_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_125_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_125_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_125_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_125_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_125_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_125_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_125_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_125_ccff_tail[0]));

	grid_clb grid_clb_11__7_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_116_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_259_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__126_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__126_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__126_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__126_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__126_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__126_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__126_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__126_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__126_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__126_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__126_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__126_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__126_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__126_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__126_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__126_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__115_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__115_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__115_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__115_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__115_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__115_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__115_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__115_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__115_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__115_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__115_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__115_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__115_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__115_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__115_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__115_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__114_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__114_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_126_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_126_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_126_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_126_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_126_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_126_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_126_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_126_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_126_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_126_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_126_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_126_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_126_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_126_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_126_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_126_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_126_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_126_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_126_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_126_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_126_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_126_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_126_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_126_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_126_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_126_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_126_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_126_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_126_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_126_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_126_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_126_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_126_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_126_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_126_ccff_tail[0]));

	grid_clb grid_clb_11__8_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_117_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_260_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__127_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__127_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__127_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__127_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__127_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__127_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__127_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__127_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__127_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__127_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__127_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__127_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__127_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__127_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__127_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__127_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__116_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__116_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__116_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__116_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__116_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__116_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__116_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__116_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__116_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__116_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__116_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__116_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__116_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__116_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__116_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__116_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__115_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__115_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_127_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_127_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_127_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_127_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_127_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_127_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_127_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_127_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_127_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_127_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_127_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_127_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_127_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_127_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_127_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_127_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_127_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_127_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_127_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_127_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_127_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_127_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_127_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_127_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_127_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_127_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_127_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_127_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_127_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_127_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_127_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_127_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_127_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_127_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_127_ccff_tail[0]));

	grid_clb grid_clb_11__9_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_118_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_261_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__128_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__128_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__128_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__128_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__128_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__128_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__128_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__128_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__128_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__128_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__128_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__128_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__128_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__128_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__128_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__128_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__117_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__117_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__117_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__117_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__117_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__117_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__117_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__117_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__117_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__117_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__117_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__117_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__117_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__117_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__117_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__117_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__116_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__116_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_128_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_128_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_128_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_128_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_128_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_128_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_128_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_128_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_128_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_128_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_128_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_128_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_128_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_128_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_128_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_128_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_128_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_128_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_128_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_128_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_128_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_128_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_128_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_128_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_128_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_128_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_128_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_128_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_128_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_128_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_128_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_128_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_128_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_128_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_128_ccff_tail[0]));

	grid_clb grid_clb_11__10_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_119_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_262_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__129_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__129_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__129_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__129_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__129_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__129_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__129_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__129_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__129_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__129_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__129_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__129_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__129_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__129_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__129_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__129_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__118_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__118_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__118_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__118_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__118_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__118_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__118_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__118_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__118_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__118_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__118_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__118_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__118_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__118_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__118_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__118_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__117_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__117_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_129_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_129_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_129_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_129_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_129_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_129_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_129_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_129_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_129_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_129_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_129_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_129_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_129_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_129_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_129_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_129_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_129_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_129_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_129_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_129_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_129_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_129_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_129_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_129_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_129_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_129_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_129_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_129_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_129_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_129_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_129_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_129_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_129_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_129_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_129_ccff_tail[0]));

	grid_clb grid_clb_11__11_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_120_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_263_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__130_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__130_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__130_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__130_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__130_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__130_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__130_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__130_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__130_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__130_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__130_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__130_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__130_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__130_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__130_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__130_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__119_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__119_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__119_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__119_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__119_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__119_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__119_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__119_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__119_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__119_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__119_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__119_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__119_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__119_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__119_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__119_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__118_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__118_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_130_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_130_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_130_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_130_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_130_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_130_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_130_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_130_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_130_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_130_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_130_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_130_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_130_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_130_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_130_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_130_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_130_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_130_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_130_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_130_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_130_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_130_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_130_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_130_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_130_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_130_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_130_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_130_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_130_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_130_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_130_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_130_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_130_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_130_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_130_ccff_tail[0]));

	grid_clb grid_clb_11__12_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_141_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_284_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__131_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__131_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__131_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__131_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__131_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__131_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__131_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__131_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__131_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__131_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__131_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__131_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__131_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__131_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__131_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__131_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__120_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__120_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__120_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__120_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__120_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__120_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__120_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__120_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__120_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__120_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__120_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__120_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__120_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__120_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__120_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__120_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__119_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__119_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_131_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_131_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_131_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_131_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_131_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_131_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_131_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_131_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_131_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_131_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_131_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_131_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_131_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_131_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_131_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_131_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_131_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_131_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_131_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_131_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_131_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_131_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_131_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_131_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_131_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_131_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_131_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_131_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_131_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_131_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_131_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_131_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_131_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_131_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_131_ccff_tail[0]));

	grid_clb grid_clb_12__1_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_121_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_264_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__132_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__132_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__132_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__132_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__132_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__132_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__132_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__132_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__132_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__132_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__132_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__132_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__132_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__132_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__132_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__132_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__0__11_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__0__11_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__0__11_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__0__11_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__0__11_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__0__11_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__0__11_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__0__11_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__0__11_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__0__11_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__0__11_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__0__11_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__0__11_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__0__11_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__0__11_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__0__11_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__120_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__120_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_132_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_132_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_132_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_132_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_132_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_132_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_132_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_132_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_132_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_132_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_132_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_132_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_132_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_132_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_132_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_132_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_132_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_132_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_132_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_132_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_132_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_132_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_132_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_132_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_132_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_132_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_132_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_132_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_132_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_132_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_132_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_132_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_12__1__undriven_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_12__1__undriven_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_132_ccff_tail[0]));

	grid_clb grid_clb_12__2_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_122_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_265_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__133_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__133_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__133_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__133_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__133_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__133_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__133_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__133_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__133_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__133_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__133_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__133_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__133_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__133_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__133_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__133_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__121_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__121_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__121_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__121_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__121_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__121_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__121_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__121_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__121_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__121_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__121_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__121_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__121_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__121_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__121_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__121_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__121_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__121_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_133_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_133_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_133_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_133_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_133_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_133_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_133_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_133_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_133_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_133_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_133_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_133_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_133_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_133_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_133_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_133_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_133_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_133_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_133_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_133_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_133_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_133_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_133_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_133_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_133_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_133_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_133_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_133_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_133_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_133_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_133_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_133_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_133_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_133_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_133_ccff_tail[0]));

	grid_clb grid_clb_12__3_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_123_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_266_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__134_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__134_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__134_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__134_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__134_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__134_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__134_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__134_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__134_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__134_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__134_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__134_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__134_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__134_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__134_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__134_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__122_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__122_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__122_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__122_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__122_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__122_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__122_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__122_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__122_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__122_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__122_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__122_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__122_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__122_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__122_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__122_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__122_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__122_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_134_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_134_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_134_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_134_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_134_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_134_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_134_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_134_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_134_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_134_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_134_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_134_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_134_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_134_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_134_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_134_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_134_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_134_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_134_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_134_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_134_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_134_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_134_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_134_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_134_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_134_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_134_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_134_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_134_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_134_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_134_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_134_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_134_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_134_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_134_ccff_tail[0]));

	grid_clb grid_clb_12__4_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_124_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_267_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__135_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__135_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__135_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__135_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__135_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__135_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__135_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__135_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__135_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__135_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__135_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__135_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__135_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__135_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__135_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__135_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__123_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__123_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__123_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__123_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__123_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__123_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__123_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__123_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__123_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__123_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__123_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__123_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__123_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__123_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__123_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__123_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__123_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__123_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_135_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_135_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_135_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_135_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_135_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_135_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_135_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_135_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_135_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_135_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_135_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_135_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_135_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_135_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_135_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_135_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_135_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_135_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_135_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_135_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_135_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_135_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_135_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_135_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_135_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_135_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_135_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_135_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_135_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_135_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_135_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_135_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_135_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_135_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_135_ccff_tail[0]));

	grid_clb grid_clb_12__5_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_125_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_268_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__136_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__136_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__136_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__136_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__136_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__136_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__136_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__136_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__136_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__136_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__136_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__136_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__136_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__136_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__136_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__136_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__124_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__124_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__124_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__124_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__124_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__124_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__124_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__124_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__124_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__124_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__124_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__124_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__124_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__124_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__124_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__124_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__124_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__124_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_136_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_136_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_136_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_136_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_136_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_136_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_136_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_136_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_136_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_136_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_136_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_136_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_136_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_136_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_136_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_136_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_136_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_136_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_136_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_136_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_136_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_136_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_136_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_136_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_136_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_136_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_136_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_136_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_136_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_136_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_136_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_136_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_136_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_136_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_136_ccff_tail[0]));

	grid_clb grid_clb_12__6_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_126_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_269_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__137_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__137_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__137_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__137_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__137_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__137_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__137_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__137_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__137_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__137_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__137_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__137_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__137_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__137_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__137_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__137_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__125_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__125_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__125_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__125_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__125_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__125_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__125_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__125_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__125_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__125_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__125_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__125_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__125_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__125_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__125_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__125_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__125_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__125_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_137_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_137_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_137_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_137_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_137_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_137_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_137_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_137_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_137_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_137_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_137_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_137_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_137_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_137_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_137_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_137_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_137_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_137_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_137_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_137_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_137_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_137_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_137_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_137_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_137_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_137_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_137_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_137_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_137_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_137_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_137_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_137_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_137_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_137_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_137_ccff_tail[0]));

	grid_clb grid_clb_12__7_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_127_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_270_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__138_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__138_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__138_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__138_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__138_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__138_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__138_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__138_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__138_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__138_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__138_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__138_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__138_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__138_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__138_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__138_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__126_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__126_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__126_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__126_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__126_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__126_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__126_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__126_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__126_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__126_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__126_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__126_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__126_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__126_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__126_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__126_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__126_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__126_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_138_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_138_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_138_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_138_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_138_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_138_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_138_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_138_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_138_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_138_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_138_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_138_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_138_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_138_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_138_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_138_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_138_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_138_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_138_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_138_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_138_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_138_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_138_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_138_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_138_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_138_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_138_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_138_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_138_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_138_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_138_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_138_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_138_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_138_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_138_ccff_tail[0]));

	grid_clb grid_clb_12__8_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_128_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_271_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__139_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__139_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__139_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__139_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__139_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__139_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__139_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__139_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__139_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__139_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__139_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__139_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__139_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__139_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__139_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__139_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__127_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__127_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__127_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__127_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__127_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__127_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__127_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__127_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__127_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__127_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__127_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__127_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__127_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__127_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__127_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__127_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__127_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__127_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_139_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_139_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_139_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_139_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_139_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_139_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_139_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_139_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_139_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_139_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_139_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_139_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_139_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_139_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_139_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_139_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_139_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_139_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_139_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_139_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_139_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_139_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_139_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_139_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_139_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_139_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_139_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_139_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_139_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_139_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_139_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_139_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_139_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_139_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_139_ccff_tail[0]));

	grid_clb grid_clb_12__9_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_129_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_272_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__140_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__140_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__140_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__140_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__140_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__140_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__140_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__140_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__140_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__140_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__140_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__140_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__140_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__140_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__140_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__140_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__128_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__128_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__128_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__128_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__128_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__128_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__128_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__128_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__128_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__128_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__128_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__128_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__128_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__128_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__128_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__128_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__128_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__128_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_140_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_140_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_140_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_140_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_140_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_140_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_140_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_140_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_140_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_140_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_140_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_140_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_140_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_140_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_140_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_140_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_140_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_140_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_140_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_140_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_140_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_140_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_140_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_140_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_140_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_140_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_140_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_140_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_140_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_140_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_140_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_140_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_140_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_140_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_140_ccff_tail[0]));

	grid_clb grid_clb_12__10_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_130_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_273_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__141_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__141_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__141_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__141_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__141_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__141_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__141_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__141_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__141_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__141_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__141_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__141_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__141_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__141_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__141_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__141_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__129_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__129_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__129_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__129_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__129_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__129_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__129_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__129_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__129_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__129_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__129_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__129_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__129_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__129_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__129_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__129_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__129_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__129_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_141_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_141_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_141_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_141_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_141_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_141_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_141_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_141_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_141_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_141_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_141_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_141_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_141_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_141_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_141_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_141_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_141_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_141_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_141_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_141_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_141_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_141_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_141_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_141_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_141_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_141_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_141_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_141_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_141_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_141_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_141_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_141_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_141_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_141_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_141_ccff_tail[0]));

	grid_clb grid_clb_12__11_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_131_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_274_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__142_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__142_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__142_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__142_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__142_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__142_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__142_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__142_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__142_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__142_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__142_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__142_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__142_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__142_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__142_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__142_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__130_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__130_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__130_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__130_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__130_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__130_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__130_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__130_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__130_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__130_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__130_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__130_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__130_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__130_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__130_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__130_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__130_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__130_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_142_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_142_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_142_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_142_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_142_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_142_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_142_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_142_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_142_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_142_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_142_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_142_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_142_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_142_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_142_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_142_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_142_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_142_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_142_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_142_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_142_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_142_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_142_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_142_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_142_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_142_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_142_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_142_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_142_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_142_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_142_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_142_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_142_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_142_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_142_ccff_tail[0]));

	grid_clb grid_clb_12__12_ (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.top_width_0_height_0__pin_32_(direct_interc_142_out[0]),
		.top_width_0_height_0__pin_33_(direct_interc_285_out[0]),
		.right_width_0_height_0__pin_0_(cby_1__1__143_left_grid_pin_0_[0]),
		.right_width_0_height_0__pin_1_(cby_1__1__143_left_grid_pin_1_[0]),
		.right_width_0_height_0__pin_2_(cby_1__1__143_left_grid_pin_2_[0]),
		.right_width_0_height_0__pin_3_(cby_1__1__143_left_grid_pin_3_[0]),
		.right_width_0_height_0__pin_4_(cby_1__1__143_left_grid_pin_4_[0]),
		.right_width_0_height_0__pin_5_(cby_1__1__143_left_grid_pin_5_[0]),
		.right_width_0_height_0__pin_6_(cby_1__1__143_left_grid_pin_6_[0]),
		.right_width_0_height_0__pin_7_(cby_1__1__143_left_grid_pin_7_[0]),
		.right_width_0_height_0__pin_8_(cby_1__1__143_left_grid_pin_8_[0]),
		.right_width_0_height_0__pin_9_(cby_1__1__143_left_grid_pin_9_[0]),
		.right_width_0_height_0__pin_10_(cby_1__1__143_left_grid_pin_10_[0]),
		.right_width_0_height_0__pin_11_(cby_1__1__143_left_grid_pin_11_[0]),
		.right_width_0_height_0__pin_12_(cby_1__1__143_left_grid_pin_12_[0]),
		.right_width_0_height_0__pin_13_(cby_1__1__143_left_grid_pin_13_[0]),
		.right_width_0_height_0__pin_14_(cby_1__1__143_left_grid_pin_14_[0]),
		.right_width_0_height_0__pin_15_(cby_1__1__143_left_grid_pin_15_[0]),
		.bottom_width_0_height_0__pin_16_(cbx_1__1__131_top_grid_pin_16_[0]),
		.bottom_width_0_height_0__pin_17_(cbx_1__1__131_top_grid_pin_17_[0]),
		.bottom_width_0_height_0__pin_18_(cbx_1__1__131_top_grid_pin_18_[0]),
		.bottom_width_0_height_0__pin_19_(cbx_1__1__131_top_grid_pin_19_[0]),
		.bottom_width_0_height_0__pin_20_(cbx_1__1__131_top_grid_pin_20_[0]),
		.bottom_width_0_height_0__pin_21_(cbx_1__1__131_top_grid_pin_21_[0]),
		.bottom_width_0_height_0__pin_22_(cbx_1__1__131_top_grid_pin_22_[0]),
		.bottom_width_0_height_0__pin_23_(cbx_1__1__131_top_grid_pin_23_[0]),
		.bottom_width_0_height_0__pin_24_(cbx_1__1__131_top_grid_pin_24_[0]),
		.bottom_width_0_height_0__pin_25_(cbx_1__1__131_top_grid_pin_25_[0]),
		.bottom_width_0_height_0__pin_26_(cbx_1__1__131_top_grid_pin_26_[0]),
		.bottom_width_0_height_0__pin_27_(cbx_1__1__131_top_grid_pin_27_[0]),
		.bottom_width_0_height_0__pin_28_(cbx_1__1__131_top_grid_pin_28_[0]),
		.bottom_width_0_height_0__pin_29_(cbx_1__1__131_top_grid_pin_29_[0]),
		.bottom_width_0_height_0__pin_30_(cbx_1__1__131_top_grid_pin_30_[0]),
		.bottom_width_0_height_0__pin_31_(cbx_1__1__131_top_grid_pin_31_[0]),
		.left_width_0_height_0__pin_52_(cby_1__1__131_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__131_ccff_tail[0]),
		.right_width_0_height_0__pin_34_upper(grid_clb_143_right_width_0_height_0__pin_34_upper[0]),
		.right_width_0_height_0__pin_34_lower(grid_clb_143_right_width_0_height_0__pin_34_lower[0]),
		.right_width_0_height_0__pin_35_upper(grid_clb_143_right_width_0_height_0__pin_35_upper[0]),
		.right_width_0_height_0__pin_35_lower(grid_clb_143_right_width_0_height_0__pin_35_lower[0]),
		.right_width_0_height_0__pin_36_upper(grid_clb_143_right_width_0_height_0__pin_36_upper[0]),
		.right_width_0_height_0__pin_36_lower(grid_clb_143_right_width_0_height_0__pin_36_lower[0]),
		.right_width_0_height_0__pin_37_upper(grid_clb_143_right_width_0_height_0__pin_37_upper[0]),
		.right_width_0_height_0__pin_37_lower(grid_clb_143_right_width_0_height_0__pin_37_lower[0]),
		.right_width_0_height_0__pin_38_upper(grid_clb_143_right_width_0_height_0__pin_38_upper[0]),
		.right_width_0_height_0__pin_38_lower(grid_clb_143_right_width_0_height_0__pin_38_lower[0]),
		.right_width_0_height_0__pin_39_upper(grid_clb_143_right_width_0_height_0__pin_39_upper[0]),
		.right_width_0_height_0__pin_39_lower(grid_clb_143_right_width_0_height_0__pin_39_lower[0]),
		.right_width_0_height_0__pin_40_upper(grid_clb_143_right_width_0_height_0__pin_40_upper[0]),
		.right_width_0_height_0__pin_40_lower(grid_clb_143_right_width_0_height_0__pin_40_lower[0]),
		.right_width_0_height_0__pin_41_upper(grid_clb_143_right_width_0_height_0__pin_41_upper[0]),
		.right_width_0_height_0__pin_41_lower(grid_clb_143_right_width_0_height_0__pin_41_lower[0]),
		.bottom_width_0_height_0__pin_42_upper(grid_clb_143_bottom_width_0_height_0__pin_42_upper[0]),
		.bottom_width_0_height_0__pin_42_lower(grid_clb_143_bottom_width_0_height_0__pin_42_lower[0]),
		.bottom_width_0_height_0__pin_43_upper(grid_clb_143_bottom_width_0_height_0__pin_43_upper[0]),
		.bottom_width_0_height_0__pin_43_lower(grid_clb_143_bottom_width_0_height_0__pin_43_lower[0]),
		.bottom_width_0_height_0__pin_44_upper(grid_clb_143_bottom_width_0_height_0__pin_44_upper[0]),
		.bottom_width_0_height_0__pin_44_lower(grid_clb_143_bottom_width_0_height_0__pin_44_lower[0]),
		.bottom_width_0_height_0__pin_45_upper(grid_clb_143_bottom_width_0_height_0__pin_45_upper[0]),
		.bottom_width_0_height_0__pin_45_lower(grid_clb_143_bottom_width_0_height_0__pin_45_lower[0]),
		.bottom_width_0_height_0__pin_46_upper(grid_clb_143_bottom_width_0_height_0__pin_46_upper[0]),
		.bottom_width_0_height_0__pin_46_lower(grid_clb_143_bottom_width_0_height_0__pin_46_lower[0]),
		.bottom_width_0_height_0__pin_47_upper(grid_clb_143_bottom_width_0_height_0__pin_47_upper[0]),
		.bottom_width_0_height_0__pin_47_lower(grid_clb_143_bottom_width_0_height_0__pin_47_lower[0]),
		.bottom_width_0_height_0__pin_48_upper(grid_clb_143_bottom_width_0_height_0__pin_48_upper[0]),
		.bottom_width_0_height_0__pin_48_lower(grid_clb_143_bottom_width_0_height_0__pin_48_lower[0]),
		.bottom_width_0_height_0__pin_49_upper(grid_clb_143_bottom_width_0_height_0__pin_49_upper[0]),
		.bottom_width_0_height_0__pin_49_lower(grid_clb_143_bottom_width_0_height_0__pin_49_lower[0]),
		.bottom_width_0_height_0__pin_50_(grid_clb_143_bottom_width_0_height_0__pin_50_[0]),
		.bottom_width_0_height_0__pin_51_(grid_clb_143_bottom_width_0_height_0__pin_51_[0]),
		.ccff_tail(grid_clb_143_ccff_tail[0]));

	grid_io_top grid_io_top_1__13_ (
		.prog_clk(prog_clk[0]),
		.gfpga_pad_GPIO_A(gfpga_pad_GPIO_A[0]),
		.gfpga_pad_GPIO_IE(gfpga_pad_GPIO_IE[0]),
		.gfpga_pad_GPIO_OE(gfpga_pad_GPIO_OE[0]),
		.gfpga_pad_GPIO_Y(gfpga_pad_GPIO_Y[0]),
		.bottom_width_0_height_0__pin_0_(cbx_1__12__0_top_grid_pin_0_[0]),
		.ccff_head(cbx_1__12__0_ccff_tail[0]),
		.bottom_width_0_height_0__pin_1_upper(grid_io_top_0_bottom_width_0_height_0__pin_1_upper[0]),
		.bottom_width_0_height_0__pin_1_lower(grid_io_top_0_bottom_width_0_height_0__pin_1_lower[0]),
		.ccff_tail(grid_io_top_0_ccff_tail[0]));

	grid_io_top grid_io_top_2__13_ (
		.prog_clk(prog_clk[0]),
		.gfpga_pad_GPIO_A(gfpga_pad_GPIO_A[1]),
		.gfpga_pad_GPIO_IE(gfpga_pad_GPIO_IE[1]),
		.gfpga_pad_GPIO_OE(gfpga_pad_GPIO_OE[1]),
		.gfpga_pad_GPIO_Y(gfpga_pad_GPIO_Y[1]),
		.bottom_width_0_height_0__pin_0_(cbx_1__12__1_top_grid_pin_0_[0]),
		.ccff_head(cbx_1__12__1_ccff_tail[0]),
		.bottom_width_0_height_0__pin_1_upper(grid_io_top_1_bottom_width_0_height_0__pin_1_upper[0]),
		.bottom_width_0_height_0__pin_1_lower(grid_io_top_1_bottom_width_0_height_0__pin_1_lower[0]),
		.ccff_tail(grid_io_top_1_ccff_tail[0]));

	grid_io_top grid_io_top_3__13_ (
		.prog_clk(prog_clk[0]),
		.gfpga_pad_GPIO_A(gfpga_pad_GPIO_A[2]),
		.gfpga_pad_GPIO_IE(gfpga_pad_GPIO_IE[2]),
		.gfpga_pad_GPIO_OE(gfpga_pad_GPIO_OE[2]),
		.gfpga_pad_GPIO_Y(gfpga_pad_GPIO_Y[2]),
		.bottom_width_0_height_0__pin_0_(cbx_1__12__2_top_grid_pin_0_[0]),
		.ccff_head(cbx_1__12__2_ccff_tail[0]),
		.bottom_width_0_height_0__pin_1_upper(grid_io_top_2_bottom_width_0_height_0__pin_1_upper[0]),
		.bottom_width_0_height_0__pin_1_lower(grid_io_top_2_bottom_width_0_height_0__pin_1_lower[0]),
		.ccff_tail(grid_io_top_2_ccff_tail[0]));

	grid_io_top grid_io_top_4__13_ (
		.prog_clk(prog_clk[0]),
		.gfpga_pad_GPIO_A(gfpga_pad_GPIO_A[3]),
		.gfpga_pad_GPIO_IE(gfpga_pad_GPIO_IE[3]),
		.gfpga_pad_GPIO_OE(gfpga_pad_GPIO_OE[3]),
		.gfpga_pad_GPIO_Y(gfpga_pad_GPIO_Y[3]),
		.bottom_width_0_height_0__pin_0_(cbx_1__12__3_top_grid_pin_0_[0]),
		.ccff_head(cbx_1__12__3_ccff_tail[0]),
		.bottom_width_0_height_0__pin_1_upper(grid_io_top_3_bottom_width_0_height_0__pin_1_upper[0]),
		.bottom_width_0_height_0__pin_1_lower(grid_io_top_3_bottom_width_0_height_0__pin_1_lower[0]),
		.ccff_tail(grid_io_top_3_ccff_tail[0]));

	grid_io_top grid_io_top_5__13_ (
		.prog_clk(prog_clk[0]),
		.gfpga_pad_GPIO_A(gfpga_pad_GPIO_A[4]),
		.gfpga_pad_GPIO_IE(gfpga_pad_GPIO_IE[4]),
		.gfpga_pad_GPIO_OE(gfpga_pad_GPIO_OE[4]),
		.gfpga_pad_GPIO_Y(gfpga_pad_GPIO_Y[4]),
		.bottom_width_0_height_0__pin_0_(cbx_1__12__4_top_grid_pin_0_[0]),
		.ccff_head(cbx_1__12__4_ccff_tail[0]),
		.bottom_width_0_height_0__pin_1_upper(grid_io_top_4_bottom_width_0_height_0__pin_1_upper[0]),
		.bottom_width_0_height_0__pin_1_lower(grid_io_top_4_bottom_width_0_height_0__pin_1_lower[0]),
		.ccff_tail(grid_io_top_4_ccff_tail[0]));

	grid_io_top grid_io_top_6__13_ (
		.prog_clk(prog_clk[0]),
		.gfpga_pad_GPIO_A(gfpga_pad_GPIO_A[5]),
		.gfpga_pad_GPIO_IE(gfpga_pad_GPIO_IE[5]),
		.gfpga_pad_GPIO_OE(gfpga_pad_GPIO_OE[5]),
		.gfpga_pad_GPIO_Y(gfpga_pad_GPIO_Y[5]),
		.bottom_width_0_height_0__pin_0_(cbx_1__12__5_top_grid_pin_0_[0]),
		.ccff_head(cbx_1__12__5_ccff_tail[0]),
		.bottom_width_0_height_0__pin_1_upper(grid_io_top_5_bottom_width_0_height_0__pin_1_upper[0]),
		.bottom_width_0_height_0__pin_1_lower(grid_io_top_5_bottom_width_0_height_0__pin_1_lower[0]),
		.ccff_tail(grid_io_top_5_ccff_tail[0]));

	grid_io_top grid_io_top_7__13_ (
		.prog_clk(prog_clk[0]),
		.gfpga_pad_GPIO_A(gfpga_pad_GPIO_A[6]),
		.gfpga_pad_GPIO_IE(gfpga_pad_GPIO_IE[6]),
		.gfpga_pad_GPIO_OE(gfpga_pad_GPIO_OE[6]),
		.gfpga_pad_GPIO_Y(gfpga_pad_GPIO_Y[6]),
		.bottom_width_0_height_0__pin_0_(cbx_1__12__6_top_grid_pin_0_[0]),
		.ccff_head(cbx_1__12__6_ccff_tail[0]),
		.bottom_width_0_height_0__pin_1_upper(grid_io_top_6_bottom_width_0_height_0__pin_1_upper[0]),
		.bottom_width_0_height_0__pin_1_lower(grid_io_top_6_bottom_width_0_height_0__pin_1_lower[0]),
		.ccff_tail(grid_io_top_6_ccff_tail[0]));

	grid_io_top grid_io_top_8__13_ (
		.prog_clk(prog_clk[0]),
		.gfpga_pad_GPIO_A(gfpga_pad_GPIO_A[7]),
		.gfpga_pad_GPIO_IE(gfpga_pad_GPIO_IE[7]),
		.gfpga_pad_GPIO_OE(gfpga_pad_GPIO_OE[7]),
		.gfpga_pad_GPIO_Y(gfpga_pad_GPIO_Y[7]),
		.bottom_width_0_height_0__pin_0_(cbx_1__12__7_top_grid_pin_0_[0]),
		.ccff_head(cbx_1__12__7_ccff_tail[0]),
		.bottom_width_0_height_0__pin_1_upper(grid_io_top_7_bottom_width_0_height_0__pin_1_upper[0]),
		.bottom_width_0_height_0__pin_1_lower(grid_io_top_7_bottom_width_0_height_0__pin_1_lower[0]),
		.ccff_tail(grid_io_top_7_ccff_tail[0]));

	grid_io_top grid_io_top_9__13_ (
		.prog_clk(prog_clk[0]),
		.gfpga_pad_GPIO_A(gfpga_pad_GPIO_A[8]),
		.gfpga_pad_GPIO_IE(gfpga_pad_GPIO_IE[8]),
		.gfpga_pad_GPIO_OE(gfpga_pad_GPIO_OE[8]),
		.gfpga_pad_GPIO_Y(gfpga_pad_GPIO_Y[8]),
		.bottom_width_0_height_0__pin_0_(cbx_1__12__8_top_grid_pin_0_[0]),
		.ccff_head(cbx_1__12__8_ccff_tail[0]),
		.bottom_width_0_height_0__pin_1_upper(grid_io_top_8_bottom_width_0_height_0__pin_1_upper[0]),
		.bottom_width_0_height_0__pin_1_lower(grid_io_top_8_bottom_width_0_height_0__pin_1_lower[0]),
		.ccff_tail(grid_io_top_8_ccff_tail[0]));

	grid_io_top grid_io_top_10__13_ (
		.prog_clk(prog_clk[0]),
		.gfpga_pad_GPIO_A(gfpga_pad_GPIO_A[9]),
		.gfpga_pad_GPIO_IE(gfpga_pad_GPIO_IE[9]),
		.gfpga_pad_GPIO_OE(gfpga_pad_GPIO_OE[9]),
		.gfpga_pad_GPIO_Y(gfpga_pad_GPIO_Y[9]),
		.bottom_width_0_height_0__pin_0_(cbx_1__12__9_top_grid_pin_0_[0]),
		.ccff_head(cbx_1__12__9_ccff_tail[0]),
		.bottom_width_0_height_0__pin_1_upper(grid_io_top_9_bottom_width_0_height_0__pin_1_upper[0]),
		.bottom_width_0_height_0__pin_1_lower(grid_io_top_9_bottom_width_0_height_0__pin_1_lower[0]),
		.ccff_tail(grid_io_top_9_ccff_tail[0]));

	grid_io_top grid_io_top_11__13_ (
		.prog_clk(prog_clk[0]),
		.gfpga_pad_GPIO_A(gfpga_pad_GPIO_A[10]),
		.gfpga_pad_GPIO_IE(gfpga_pad_GPIO_IE[10]),
		.gfpga_pad_GPIO_OE(gfpga_pad_GPIO_OE[10]),
		.gfpga_pad_GPIO_Y(gfpga_pad_GPIO_Y[10]),
		.bottom_width_0_height_0__pin_0_(cbx_1__12__10_top_grid_pin_0_[0]),
		.ccff_head(cbx_1__12__10_ccff_tail[0]),
		.bottom_width_0_height_0__pin_1_upper(grid_io_top_10_bottom_width_0_height_0__pin_1_upper[0]),
		.bottom_width_0_height_0__pin_1_lower(grid_io_top_10_bottom_width_0_height_0__pin_1_lower[0]),
		.ccff_tail(grid_io_top_10_ccff_tail[0]));

	grid_io_top grid_io_top_12__13_ (
		.prog_clk(prog_clk[0]),
		.gfpga_pad_GPIO_A(gfpga_pad_GPIO_A[11]),
		.gfpga_pad_GPIO_IE(gfpga_pad_GPIO_IE[11]),
		.gfpga_pad_GPIO_OE(gfpga_pad_GPIO_OE[11]),
		.gfpga_pad_GPIO_Y(gfpga_pad_GPIO_Y[11]),
		.bottom_width_0_height_0__pin_0_(cbx_1__12__11_top_grid_pin_0_[0]),
		.ccff_head(cbx_1__12__11_ccff_tail[0]),
		.bottom_width_0_height_0__pin_1_upper(grid_io_top_11_bottom_width_0_height_0__pin_1_upper[0]),
		.bottom_width_0_height_0__pin_1_lower(grid_io_top_11_bottom_width_0_height_0__pin_1_lower[0]),
		.ccff_tail(grid_io_top_11_ccff_tail[0]));

	grid_io_right grid_io_right_13__1_ (
		.prog_clk(prog_clk[0]),
		.gfpga_pad_GPIO_A(gfpga_pad_GPIO_A[12]),
		.gfpga_pad_GPIO_IE(gfpga_pad_GPIO_IE[12]),
		.gfpga_pad_GPIO_OE(gfpga_pad_GPIO_OE[12]),
		.gfpga_pad_GPIO_Y(gfpga_pad_GPIO_Y[12]),
		.left_width_0_height_0__pin_0_(cby_1__1__132_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__132_ccff_tail[0]),
		.left_width_0_height_0__pin_1_upper(grid_io_right_0_left_width_0_height_0__pin_1_upper[0]),
		.left_width_0_height_0__pin_1_lower(grid_io_right_0_left_width_0_height_0__pin_1_lower[0]),
		.ccff_tail(grid_io_right_0_ccff_tail[0]));

	grid_io_right grid_io_right_13__2_ (
		.prog_clk(prog_clk[0]),
		.gfpga_pad_GPIO_A(gfpga_pad_GPIO_A[13]),
		.gfpga_pad_GPIO_IE(gfpga_pad_GPIO_IE[13]),
		.gfpga_pad_GPIO_OE(gfpga_pad_GPIO_OE[13]),
		.gfpga_pad_GPIO_Y(gfpga_pad_GPIO_Y[13]),
		.left_width_0_height_0__pin_0_(cby_1__1__133_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__133_ccff_tail[0]),
		.left_width_0_height_0__pin_1_upper(grid_io_right_1_left_width_0_height_0__pin_1_upper[0]),
		.left_width_0_height_0__pin_1_lower(grid_io_right_1_left_width_0_height_0__pin_1_lower[0]),
		.ccff_tail(grid_io_right_1_ccff_tail[0]));

	grid_io_right grid_io_right_13__3_ (
		.prog_clk(prog_clk[0]),
		.gfpga_pad_GPIO_A(gfpga_pad_GPIO_A[14]),
		.gfpga_pad_GPIO_IE(gfpga_pad_GPIO_IE[14]),
		.gfpga_pad_GPIO_OE(gfpga_pad_GPIO_OE[14]),
		.gfpga_pad_GPIO_Y(gfpga_pad_GPIO_Y[14]),
		.left_width_0_height_0__pin_0_(cby_1__1__134_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__134_ccff_tail[0]),
		.left_width_0_height_0__pin_1_upper(grid_io_right_2_left_width_0_height_0__pin_1_upper[0]),
		.left_width_0_height_0__pin_1_lower(grid_io_right_2_left_width_0_height_0__pin_1_lower[0]),
		.ccff_tail(grid_io_right_2_ccff_tail[0]));

	grid_io_right grid_io_right_13__4_ (
		.prog_clk(prog_clk[0]),
		.gfpga_pad_GPIO_A(gfpga_pad_GPIO_A[15]),
		.gfpga_pad_GPIO_IE(gfpga_pad_GPIO_IE[15]),
		.gfpga_pad_GPIO_OE(gfpga_pad_GPIO_OE[15]),
		.gfpga_pad_GPIO_Y(gfpga_pad_GPIO_Y[15]),
		.left_width_0_height_0__pin_0_(cby_1__1__135_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__135_ccff_tail[0]),
		.left_width_0_height_0__pin_1_upper(grid_io_right_3_left_width_0_height_0__pin_1_upper[0]),
		.left_width_0_height_0__pin_1_lower(grid_io_right_3_left_width_0_height_0__pin_1_lower[0]),
		.ccff_tail(grid_io_right_3_ccff_tail[0]));

	grid_io_right grid_io_right_13__5_ (
		.prog_clk(prog_clk[0]),
		.gfpga_pad_GPIO_A(gfpga_pad_GPIO_A[16]),
		.gfpga_pad_GPIO_IE(gfpga_pad_GPIO_IE[16]),
		.gfpga_pad_GPIO_OE(gfpga_pad_GPIO_OE[16]),
		.gfpga_pad_GPIO_Y(gfpga_pad_GPIO_Y[16]),
		.left_width_0_height_0__pin_0_(cby_1__1__136_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__136_ccff_tail[0]),
		.left_width_0_height_0__pin_1_upper(grid_io_right_4_left_width_0_height_0__pin_1_upper[0]),
		.left_width_0_height_0__pin_1_lower(grid_io_right_4_left_width_0_height_0__pin_1_lower[0]),
		.ccff_tail(grid_io_right_4_ccff_tail[0]));

	grid_io_right grid_io_right_13__6_ (
		.prog_clk(prog_clk[0]),
		.gfpga_pad_GPIO_A(gfpga_pad_GPIO_A[17]),
		.gfpga_pad_GPIO_IE(gfpga_pad_GPIO_IE[17]),
		.gfpga_pad_GPIO_OE(gfpga_pad_GPIO_OE[17]),
		.gfpga_pad_GPIO_Y(gfpga_pad_GPIO_Y[17]),
		.left_width_0_height_0__pin_0_(cby_1__1__137_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__137_ccff_tail[0]),
		.left_width_0_height_0__pin_1_upper(grid_io_right_5_left_width_0_height_0__pin_1_upper[0]),
		.left_width_0_height_0__pin_1_lower(grid_io_right_5_left_width_0_height_0__pin_1_lower[0]),
		.ccff_tail(grid_io_right_5_ccff_tail[0]));

	grid_io_right grid_io_right_13__7_ (
		.prog_clk(prog_clk[0]),
		.gfpga_pad_GPIO_A(gfpga_pad_GPIO_A[18]),
		.gfpga_pad_GPIO_IE(gfpga_pad_GPIO_IE[18]),
		.gfpga_pad_GPIO_OE(gfpga_pad_GPIO_OE[18]),
		.gfpga_pad_GPIO_Y(gfpga_pad_GPIO_Y[18]),
		.left_width_0_height_0__pin_0_(cby_1__1__138_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__138_ccff_tail[0]),
		.left_width_0_height_0__pin_1_upper(grid_io_right_6_left_width_0_height_0__pin_1_upper[0]),
		.left_width_0_height_0__pin_1_lower(grid_io_right_6_left_width_0_height_0__pin_1_lower[0]),
		.ccff_tail(grid_io_right_6_ccff_tail[0]));

	grid_io_right grid_io_right_13__8_ (
		.prog_clk(prog_clk[0]),
		.gfpga_pad_GPIO_A(gfpga_pad_GPIO_A[19]),
		.gfpga_pad_GPIO_IE(gfpga_pad_GPIO_IE[19]),
		.gfpga_pad_GPIO_OE(gfpga_pad_GPIO_OE[19]),
		.gfpga_pad_GPIO_Y(gfpga_pad_GPIO_Y[19]),
		.left_width_0_height_0__pin_0_(cby_1__1__139_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__139_ccff_tail[0]),
		.left_width_0_height_0__pin_1_upper(grid_io_right_7_left_width_0_height_0__pin_1_upper[0]),
		.left_width_0_height_0__pin_1_lower(grid_io_right_7_left_width_0_height_0__pin_1_lower[0]),
		.ccff_tail(grid_io_right_7_ccff_tail[0]));

	grid_io_right grid_io_right_13__9_ (
		.prog_clk(prog_clk[0]),
		.gfpga_pad_GPIO_A(gfpga_pad_GPIO_A[20]),
		.gfpga_pad_GPIO_IE(gfpga_pad_GPIO_IE[20]),
		.gfpga_pad_GPIO_OE(gfpga_pad_GPIO_OE[20]),
		.gfpga_pad_GPIO_Y(gfpga_pad_GPIO_Y[20]),
		.left_width_0_height_0__pin_0_(cby_1__1__140_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__140_ccff_tail[0]),
		.left_width_0_height_0__pin_1_upper(grid_io_right_8_left_width_0_height_0__pin_1_upper[0]),
		.left_width_0_height_0__pin_1_lower(grid_io_right_8_left_width_0_height_0__pin_1_lower[0]),
		.ccff_tail(grid_io_right_8_ccff_tail[0]));

	grid_io_right grid_io_right_13__10_ (
		.prog_clk(prog_clk[0]),
		.gfpga_pad_GPIO_A(gfpga_pad_GPIO_A[21]),
		.gfpga_pad_GPIO_IE(gfpga_pad_GPIO_IE[21]),
		.gfpga_pad_GPIO_OE(gfpga_pad_GPIO_OE[21]),
		.gfpga_pad_GPIO_Y(gfpga_pad_GPIO_Y[21]),
		.left_width_0_height_0__pin_0_(cby_1__1__141_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__141_ccff_tail[0]),
		.left_width_0_height_0__pin_1_upper(grid_io_right_9_left_width_0_height_0__pin_1_upper[0]),
		.left_width_0_height_0__pin_1_lower(grid_io_right_9_left_width_0_height_0__pin_1_lower[0]),
		.ccff_tail(grid_io_right_9_ccff_tail[0]));

	grid_io_right grid_io_right_13__11_ (
		.prog_clk(prog_clk[0]),
		.gfpga_pad_GPIO_A(gfpga_pad_GPIO_A[22]),
		.gfpga_pad_GPIO_IE(gfpga_pad_GPIO_IE[22]),
		.gfpga_pad_GPIO_OE(gfpga_pad_GPIO_OE[22]),
		.gfpga_pad_GPIO_Y(gfpga_pad_GPIO_Y[22]),
		.left_width_0_height_0__pin_0_(cby_1__1__142_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__142_ccff_tail[0]),
		.left_width_0_height_0__pin_1_upper(grid_io_right_10_left_width_0_height_0__pin_1_upper[0]),
		.left_width_0_height_0__pin_1_lower(grid_io_right_10_left_width_0_height_0__pin_1_lower[0]),
		.ccff_tail(grid_io_right_10_ccff_tail[0]));

	grid_io_right grid_io_right_13__12_ (
		.prog_clk(prog_clk[0]),
		.gfpga_pad_GPIO_A(gfpga_pad_GPIO_A[23]),
		.gfpga_pad_GPIO_IE(gfpga_pad_GPIO_IE[23]),
		.gfpga_pad_GPIO_OE(gfpga_pad_GPIO_OE[23]),
		.gfpga_pad_GPIO_Y(gfpga_pad_GPIO_Y[23]),
		.left_width_0_height_0__pin_0_(cby_1__1__143_right_grid_pin_52_[0]),
		.ccff_head(cby_1__1__143_ccff_tail[0]),
		.left_width_0_height_0__pin_1_upper(grid_io_right_11_left_width_0_height_0__pin_1_upper[0]),
		.left_width_0_height_0__pin_1_lower(grid_io_right_11_left_width_0_height_0__pin_1_lower[0]),
		.ccff_tail(grid_io_right_11_ccff_tail[0]));

	grid_io_bottom grid_io_bottom_1__0_ (
		.prog_clk(prog_clk[0]),
		.gfpga_pad_GPIO_A(gfpga_pad_GPIO_A[24]),
		.gfpga_pad_GPIO_IE(gfpga_pad_GPIO_IE[24]),
		.gfpga_pad_GPIO_OE(gfpga_pad_GPIO_OE[24]),
		.gfpga_pad_GPIO_Y(gfpga_pad_GPIO_Y[24]),
		.top_width_0_height_0__pin_0_(cbx_1__0__0_bottom_grid_pin_0_[0]),
		.ccff_head(cbx_1__0__0_ccff_tail[0]),
		.top_width_0_height_0__pin_1_upper(grid_io_bottom_0_top_width_0_height_0__pin_1_upper[0]),
		.top_width_0_height_0__pin_1_lower(grid_io_bottom_0_top_width_0_height_0__pin_1_lower[0]),
		.ccff_tail(grid_io_bottom_0_ccff_tail[0]));

	grid_io_bottom grid_io_bottom_2__0_ (
		.prog_clk(prog_clk[0]),
		.gfpga_pad_GPIO_A(gfpga_pad_GPIO_A[25]),
		.gfpga_pad_GPIO_IE(gfpga_pad_GPIO_IE[25]),
		.gfpga_pad_GPIO_OE(gfpga_pad_GPIO_OE[25]),
		.gfpga_pad_GPIO_Y(gfpga_pad_GPIO_Y[25]),
		.top_width_0_height_0__pin_0_(cbx_1__0__1_bottom_grid_pin_0_[0]),
		.ccff_head(cbx_1__0__1_ccff_tail[0]),
		.top_width_0_height_0__pin_1_upper(grid_io_bottom_1_top_width_0_height_0__pin_1_upper[0]),
		.top_width_0_height_0__pin_1_lower(grid_io_bottom_1_top_width_0_height_0__pin_1_lower[0]),
		.ccff_tail(grid_io_bottom_1_ccff_tail[0]));

	grid_io_bottom grid_io_bottom_3__0_ (
		.prog_clk(prog_clk[0]),
		.gfpga_pad_GPIO_A(gfpga_pad_GPIO_A[26]),
		.gfpga_pad_GPIO_IE(gfpga_pad_GPIO_IE[26]),
		.gfpga_pad_GPIO_OE(gfpga_pad_GPIO_OE[26]),
		.gfpga_pad_GPIO_Y(gfpga_pad_GPIO_Y[26]),
		.top_width_0_height_0__pin_0_(cbx_1__0__2_bottom_grid_pin_0_[0]),
		.ccff_head(cbx_1__0__2_ccff_tail[0]),
		.top_width_0_height_0__pin_1_upper(grid_io_bottom_2_top_width_0_height_0__pin_1_upper[0]),
		.top_width_0_height_0__pin_1_lower(grid_io_bottom_2_top_width_0_height_0__pin_1_lower[0]),
		.ccff_tail(grid_io_bottom_2_ccff_tail[0]));

	grid_io_bottom grid_io_bottom_4__0_ (
		.prog_clk(prog_clk[0]),
		.gfpga_pad_GPIO_A(gfpga_pad_GPIO_A[27]),
		.gfpga_pad_GPIO_IE(gfpga_pad_GPIO_IE[27]),
		.gfpga_pad_GPIO_OE(gfpga_pad_GPIO_OE[27]),
		.gfpga_pad_GPIO_Y(gfpga_pad_GPIO_Y[27]),
		.top_width_0_height_0__pin_0_(cbx_1__0__3_bottom_grid_pin_0_[0]),
		.ccff_head(cbx_1__0__3_ccff_tail[0]),
		.top_width_0_height_0__pin_1_upper(grid_io_bottom_3_top_width_0_height_0__pin_1_upper[0]),
		.top_width_0_height_0__pin_1_lower(grid_io_bottom_3_top_width_0_height_0__pin_1_lower[0]),
		.ccff_tail(grid_io_bottom_3_ccff_tail[0]));

	grid_io_bottom grid_io_bottom_5__0_ (
		.prog_clk(prog_clk[0]),
		.gfpga_pad_GPIO_A(gfpga_pad_GPIO_A[28]),
		.gfpga_pad_GPIO_IE(gfpga_pad_GPIO_IE[28]),
		.gfpga_pad_GPIO_OE(gfpga_pad_GPIO_OE[28]),
		.gfpga_pad_GPIO_Y(gfpga_pad_GPIO_Y[28]),
		.top_width_0_height_0__pin_0_(cbx_1__0__4_bottom_grid_pin_0_[0]),
		.ccff_head(cbx_1__0__4_ccff_tail[0]),
		.top_width_0_height_0__pin_1_upper(grid_io_bottom_4_top_width_0_height_0__pin_1_upper[0]),
		.top_width_0_height_0__pin_1_lower(grid_io_bottom_4_top_width_0_height_0__pin_1_lower[0]),
		.ccff_tail(grid_io_bottom_4_ccff_tail[0]));

	grid_io_bottom grid_io_bottom_6__0_ (
		.prog_clk(prog_clk[0]),
		.gfpga_pad_GPIO_A(gfpga_pad_GPIO_A[29]),
		.gfpga_pad_GPIO_IE(gfpga_pad_GPIO_IE[29]),
		.gfpga_pad_GPIO_OE(gfpga_pad_GPIO_OE[29]),
		.gfpga_pad_GPIO_Y(gfpga_pad_GPIO_Y[29]),
		.top_width_0_height_0__pin_0_(cbx_1__0__5_bottom_grid_pin_0_[0]),
		.ccff_head(cbx_1__0__5_ccff_tail[0]),
		.top_width_0_height_0__pin_1_upper(grid_io_bottom_5_top_width_0_height_0__pin_1_upper[0]),
		.top_width_0_height_0__pin_1_lower(grid_io_bottom_5_top_width_0_height_0__pin_1_lower[0]),
		.ccff_tail(grid_io_bottom_5_ccff_tail[0]));

	grid_io_bottom grid_io_bottom_7__0_ (
		.prog_clk(prog_clk[0]),
		.gfpga_pad_GPIO_A(gfpga_pad_GPIO_A[30]),
		.gfpga_pad_GPIO_IE(gfpga_pad_GPIO_IE[30]),
		.gfpga_pad_GPIO_OE(gfpga_pad_GPIO_OE[30]),
		.gfpga_pad_GPIO_Y(gfpga_pad_GPIO_Y[30]),
		.top_width_0_height_0__pin_0_(cbx_1__0__6_bottom_grid_pin_0_[0]),
		.ccff_head(cbx_1__0__6_ccff_tail[0]),
		.top_width_0_height_0__pin_1_upper(grid_io_bottom_6_top_width_0_height_0__pin_1_upper[0]),
		.top_width_0_height_0__pin_1_lower(grid_io_bottom_6_top_width_0_height_0__pin_1_lower[0]),
		.ccff_tail(grid_io_bottom_6_ccff_tail[0]));

	grid_io_bottom grid_io_bottom_8__0_ (
		.prog_clk(prog_clk[0]),
		.gfpga_pad_GPIO_A(gfpga_pad_GPIO_A[31]),
		.gfpga_pad_GPIO_IE(gfpga_pad_GPIO_IE[31]),
		.gfpga_pad_GPIO_OE(gfpga_pad_GPIO_OE[31]),
		.gfpga_pad_GPIO_Y(gfpga_pad_GPIO_Y[31]),
		.top_width_0_height_0__pin_0_(cbx_1__0__7_bottom_grid_pin_0_[0]),
		.ccff_head(cbx_1__0__7_ccff_tail[0]),
		.top_width_0_height_0__pin_1_upper(grid_io_bottom_7_top_width_0_height_0__pin_1_upper[0]),
		.top_width_0_height_0__pin_1_lower(grid_io_bottom_7_top_width_0_height_0__pin_1_lower[0]),
		.ccff_tail(grid_io_bottom_7_ccff_tail[0]));

	grid_io_bottom grid_io_bottom_9__0_ (
		.prog_clk(prog_clk[0]),
		.gfpga_pad_GPIO_A(gfpga_pad_GPIO_A[32]),
		.gfpga_pad_GPIO_IE(gfpga_pad_GPIO_IE[32]),
		.gfpga_pad_GPIO_OE(gfpga_pad_GPIO_OE[32]),
		.gfpga_pad_GPIO_Y(gfpga_pad_GPIO_Y[32]),
		.top_width_0_height_0__pin_0_(cbx_1__0__8_bottom_grid_pin_0_[0]),
		.ccff_head(cbx_1__0__8_ccff_tail[0]),
		.top_width_0_height_0__pin_1_upper(grid_io_bottom_8_top_width_0_height_0__pin_1_upper[0]),
		.top_width_0_height_0__pin_1_lower(grid_io_bottom_8_top_width_0_height_0__pin_1_lower[0]),
		.ccff_tail(grid_io_bottom_8_ccff_tail[0]));

	grid_io_bottom grid_io_bottom_10__0_ (
		.prog_clk(prog_clk[0]),
		.gfpga_pad_GPIO_A(gfpga_pad_GPIO_A[33]),
		.gfpga_pad_GPIO_IE(gfpga_pad_GPIO_IE[33]),
		.gfpga_pad_GPIO_OE(gfpga_pad_GPIO_OE[33]),
		.gfpga_pad_GPIO_Y(gfpga_pad_GPIO_Y[33]),
		.top_width_0_height_0__pin_0_(cbx_1__0__9_bottom_grid_pin_0_[0]),
		.ccff_head(cbx_1__0__9_ccff_tail[0]),
		.top_width_0_height_0__pin_1_upper(grid_io_bottom_9_top_width_0_height_0__pin_1_upper[0]),
		.top_width_0_height_0__pin_1_lower(grid_io_bottom_9_top_width_0_height_0__pin_1_lower[0]),
		.ccff_tail(grid_io_bottom_9_ccff_tail[0]));

	grid_io_bottom grid_io_bottom_11__0_ (
		.prog_clk(prog_clk[0]),
		.gfpga_pad_GPIO_A(gfpga_pad_GPIO_A[34]),
		.gfpga_pad_GPIO_IE(gfpga_pad_GPIO_IE[34]),
		.gfpga_pad_GPIO_OE(gfpga_pad_GPIO_OE[34]),
		.gfpga_pad_GPIO_Y(gfpga_pad_GPIO_Y[34]),
		.top_width_0_height_0__pin_0_(cbx_1__0__10_bottom_grid_pin_0_[0]),
		.ccff_head(cbx_1__0__10_ccff_tail[0]),
		.top_width_0_height_0__pin_1_upper(grid_io_bottom_10_top_width_0_height_0__pin_1_upper[0]),
		.top_width_0_height_0__pin_1_lower(grid_io_bottom_10_top_width_0_height_0__pin_1_lower[0]),
		.ccff_tail(grid_io_bottom_10_ccff_tail[0]));

	grid_io_bottom grid_io_bottom_12__0_ (
		.prog_clk(prog_clk[0]),
		.gfpga_pad_GPIO_A(gfpga_pad_GPIO_A[35]),
		.gfpga_pad_GPIO_IE(gfpga_pad_GPIO_IE[35]),
		.gfpga_pad_GPIO_OE(gfpga_pad_GPIO_OE[35]),
		.gfpga_pad_GPIO_Y(gfpga_pad_GPIO_Y[35]),
		.top_width_0_height_0__pin_0_(cbx_1__0__11_bottom_grid_pin_0_[0]),
		.ccff_head(cbx_1__0__11_ccff_tail[0]),
		.top_width_0_height_0__pin_1_upper(grid_io_bottom_11_top_width_0_height_0__pin_1_upper[0]),
		.top_width_0_height_0__pin_1_lower(grid_io_bottom_11_top_width_0_height_0__pin_1_lower[0]),
		.ccff_tail(grid_io_bottom_11_ccff_tail[0]));

	grid_io_left grid_io_left_0__1_ (
		.prog_clk(prog_clk[0]),
		.gfpga_pad_GPIO_A(gfpga_pad_GPIO_A[36]),
		.gfpga_pad_GPIO_IE(gfpga_pad_GPIO_IE[36]),
		.gfpga_pad_GPIO_OE(gfpga_pad_GPIO_OE[36]),
		.gfpga_pad_GPIO_Y(gfpga_pad_GPIO_Y[36]),
		.right_width_0_height_0__pin_0_(cby_0__1__0_left_grid_pin_0_[0]),
		.ccff_head(cby_0__1__0_ccff_tail[0]),
		.right_width_0_height_0__pin_1_upper(grid_io_left_0_right_width_0_height_0__pin_1_upper[0]),
		.right_width_0_height_0__pin_1_lower(grid_io_left_0_right_width_0_height_0__pin_1_lower[0]),
		.ccff_tail(grid_io_left_0_ccff_tail[0]));

	grid_io_left grid_io_left_0__2_ (
		.prog_clk(prog_clk[0]),
		.gfpga_pad_GPIO_A(gfpga_pad_GPIO_A[37]),
		.gfpga_pad_GPIO_IE(gfpga_pad_GPIO_IE[37]),
		.gfpga_pad_GPIO_OE(gfpga_pad_GPIO_OE[37]),
		.gfpga_pad_GPIO_Y(gfpga_pad_GPIO_Y[37]),
		.right_width_0_height_0__pin_0_(cby_0__1__1_left_grid_pin_0_[0]),
		.ccff_head(cby_0__1__1_ccff_tail[0]),
		.right_width_0_height_0__pin_1_upper(grid_io_left_1_right_width_0_height_0__pin_1_upper[0]),
		.right_width_0_height_0__pin_1_lower(grid_io_left_1_right_width_0_height_0__pin_1_lower[0]),
		.ccff_tail(grid_io_left_1_ccff_tail[0]));

	grid_io_left grid_io_left_0__3_ (
		.prog_clk(prog_clk[0]),
		.gfpga_pad_GPIO_A(gfpga_pad_GPIO_A[38]),
		.gfpga_pad_GPIO_IE(gfpga_pad_GPIO_IE[38]),
		.gfpga_pad_GPIO_OE(gfpga_pad_GPIO_OE[38]),
		.gfpga_pad_GPIO_Y(gfpga_pad_GPIO_Y[38]),
		.right_width_0_height_0__pin_0_(cby_0__1__2_left_grid_pin_0_[0]),
		.ccff_head(cby_0__1__2_ccff_tail[0]),
		.right_width_0_height_0__pin_1_upper(grid_io_left_2_right_width_0_height_0__pin_1_upper[0]),
		.right_width_0_height_0__pin_1_lower(grid_io_left_2_right_width_0_height_0__pin_1_lower[0]),
		.ccff_tail(grid_io_left_2_ccff_tail[0]));

	grid_io_left grid_io_left_0__4_ (
		.prog_clk(prog_clk[0]),
		.gfpga_pad_GPIO_A(gfpga_pad_GPIO_A[39]),
		.gfpga_pad_GPIO_IE(gfpga_pad_GPIO_IE[39]),
		.gfpga_pad_GPIO_OE(gfpga_pad_GPIO_OE[39]),
		.gfpga_pad_GPIO_Y(gfpga_pad_GPIO_Y[39]),
		.right_width_0_height_0__pin_0_(cby_0__1__3_left_grid_pin_0_[0]),
		.ccff_head(cby_0__1__3_ccff_tail[0]),
		.right_width_0_height_0__pin_1_upper(grid_io_left_3_right_width_0_height_0__pin_1_upper[0]),
		.right_width_0_height_0__pin_1_lower(grid_io_left_3_right_width_0_height_0__pin_1_lower[0]),
		.ccff_tail(grid_io_left_3_ccff_tail[0]));

	grid_io_left grid_io_left_0__5_ (
		.prog_clk(prog_clk[0]),
		.gfpga_pad_GPIO_A(gfpga_pad_GPIO_A[40]),
		.gfpga_pad_GPIO_IE(gfpga_pad_GPIO_IE[40]),
		.gfpga_pad_GPIO_OE(gfpga_pad_GPIO_OE[40]),
		.gfpga_pad_GPIO_Y(gfpga_pad_GPIO_Y[40]),
		.right_width_0_height_0__pin_0_(cby_0__1__4_left_grid_pin_0_[0]),
		.ccff_head(cby_0__1__4_ccff_tail[0]),
		.right_width_0_height_0__pin_1_upper(grid_io_left_4_right_width_0_height_0__pin_1_upper[0]),
		.right_width_0_height_0__pin_1_lower(grid_io_left_4_right_width_0_height_0__pin_1_lower[0]),
		.ccff_tail(grid_io_left_4_ccff_tail[0]));

	grid_io_left grid_io_left_0__6_ (
		.prog_clk(prog_clk[0]),
		.gfpga_pad_GPIO_A(gfpga_pad_GPIO_A[41]),
		.gfpga_pad_GPIO_IE(gfpga_pad_GPIO_IE[41]),
		.gfpga_pad_GPIO_OE(gfpga_pad_GPIO_OE[41]),
		.gfpga_pad_GPIO_Y(gfpga_pad_GPIO_Y[41]),
		.right_width_0_height_0__pin_0_(cby_0__1__5_left_grid_pin_0_[0]),
		.ccff_head(cby_0__1__5_ccff_tail[0]),
		.right_width_0_height_0__pin_1_upper(grid_io_left_5_right_width_0_height_0__pin_1_upper[0]),
		.right_width_0_height_0__pin_1_lower(grid_io_left_5_right_width_0_height_0__pin_1_lower[0]),
		.ccff_tail(grid_io_left_5_ccff_tail[0]));

	grid_io_left grid_io_left_0__7_ (
		.prog_clk(prog_clk[0]),
		.gfpga_pad_GPIO_A(gfpga_pad_GPIO_A[42]),
		.gfpga_pad_GPIO_IE(gfpga_pad_GPIO_IE[42]),
		.gfpga_pad_GPIO_OE(gfpga_pad_GPIO_OE[42]),
		.gfpga_pad_GPIO_Y(gfpga_pad_GPIO_Y[42]),
		.right_width_0_height_0__pin_0_(cby_0__1__6_left_grid_pin_0_[0]),
		.ccff_head(cby_0__1__6_ccff_tail[0]),
		.right_width_0_height_0__pin_1_upper(grid_io_left_6_right_width_0_height_0__pin_1_upper[0]),
		.right_width_0_height_0__pin_1_lower(grid_io_left_6_right_width_0_height_0__pin_1_lower[0]),
		.ccff_tail(grid_io_left_6_ccff_tail[0]));

	grid_io_left grid_io_left_0__8_ (
		.prog_clk(prog_clk[0]),
		.gfpga_pad_GPIO_A(gfpga_pad_GPIO_A[43]),
		.gfpga_pad_GPIO_IE(gfpga_pad_GPIO_IE[43]),
		.gfpga_pad_GPIO_OE(gfpga_pad_GPIO_OE[43]),
		.gfpga_pad_GPIO_Y(gfpga_pad_GPIO_Y[43]),
		.right_width_0_height_0__pin_0_(cby_0__1__7_left_grid_pin_0_[0]),
		.ccff_head(cby_0__1__7_ccff_tail[0]),
		.right_width_0_height_0__pin_1_upper(grid_io_left_7_right_width_0_height_0__pin_1_upper[0]),
		.right_width_0_height_0__pin_1_lower(grid_io_left_7_right_width_0_height_0__pin_1_lower[0]),
		.ccff_tail(grid_io_left_7_ccff_tail[0]));

	grid_io_left grid_io_left_0__9_ (
		.prog_clk(prog_clk[0]),
		.gfpga_pad_GPIO_A(gfpga_pad_GPIO_A[44]),
		.gfpga_pad_GPIO_IE(gfpga_pad_GPIO_IE[44]),
		.gfpga_pad_GPIO_OE(gfpga_pad_GPIO_OE[44]),
		.gfpga_pad_GPIO_Y(gfpga_pad_GPIO_Y[44]),
		.right_width_0_height_0__pin_0_(cby_0__1__8_left_grid_pin_0_[0]),
		.ccff_head(cby_0__1__8_ccff_tail[0]),
		.right_width_0_height_0__pin_1_upper(grid_io_left_8_right_width_0_height_0__pin_1_upper[0]),
		.right_width_0_height_0__pin_1_lower(grid_io_left_8_right_width_0_height_0__pin_1_lower[0]),
		.ccff_tail(grid_io_left_8_ccff_tail[0]));

	grid_io_left grid_io_left_0__10_ (
		.prog_clk(prog_clk[0]),
		.gfpga_pad_GPIO_A(gfpga_pad_GPIO_A[45]),
		.gfpga_pad_GPIO_IE(gfpga_pad_GPIO_IE[45]),
		.gfpga_pad_GPIO_OE(gfpga_pad_GPIO_OE[45]),
		.gfpga_pad_GPIO_Y(gfpga_pad_GPIO_Y[45]),
		.right_width_0_height_0__pin_0_(cby_0__1__9_left_grid_pin_0_[0]),
		.ccff_head(cby_0__1__9_ccff_tail[0]),
		.right_width_0_height_0__pin_1_upper(grid_io_left_9_right_width_0_height_0__pin_1_upper[0]),
		.right_width_0_height_0__pin_1_lower(grid_io_left_9_right_width_0_height_0__pin_1_lower[0]),
		.ccff_tail(grid_io_left_9_ccff_tail[0]));

	grid_io_left grid_io_left_0__11_ (
		.prog_clk(prog_clk[0]),
		.gfpga_pad_GPIO_A(gfpga_pad_GPIO_A[46]),
		.gfpga_pad_GPIO_IE(gfpga_pad_GPIO_IE[46]),
		.gfpga_pad_GPIO_OE(gfpga_pad_GPIO_OE[46]),
		.gfpga_pad_GPIO_Y(gfpga_pad_GPIO_Y[46]),
		.right_width_0_height_0__pin_0_(cby_0__1__10_left_grid_pin_0_[0]),
		.ccff_head(cby_0__1__10_ccff_tail[0]),
		.right_width_0_height_0__pin_1_upper(grid_io_left_10_right_width_0_height_0__pin_1_upper[0]),
		.right_width_0_height_0__pin_1_lower(grid_io_left_10_right_width_0_height_0__pin_1_lower[0]),
		.ccff_tail(grid_io_left_10_ccff_tail[0]));

	grid_io_left grid_io_left_0__12_ (
		.prog_clk(prog_clk[0]),
		.gfpga_pad_GPIO_A(gfpga_pad_GPIO_A[47]),
		.gfpga_pad_GPIO_IE(gfpga_pad_GPIO_IE[47]),
		.gfpga_pad_GPIO_OE(gfpga_pad_GPIO_OE[47]),
		.gfpga_pad_GPIO_Y(gfpga_pad_GPIO_Y[47]),
		.right_width_0_height_0__pin_0_(cby_0__1__11_left_grid_pin_0_[0]),
		.ccff_head(cby_0__1__11_ccff_tail[0]),
		.right_width_0_height_0__pin_1_upper(grid_io_left_11_right_width_0_height_0__pin_1_upper[0]),
		.right_width_0_height_0__pin_1_lower(grid_io_left_11_right_width_0_height_0__pin_1_lower[0]),
		.ccff_tail(grid_io_left_11_ccff_tail[0]));

	sb_0__0_ sb_0__0_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_0__1__0_chany_bottom_out[0:19]),
		.top_left_grid_pin_1_(grid_io_left_0_right_width_0_height_0__pin_1_lower[0]),
		.chanx_right_in(cbx_1__0__0_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_0_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_0_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_0_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_0_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_0_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_0_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_0_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_0_bottom_width_0_height_0__pin_49_upper[0]),
		.right_bottom_grid_pin_1_(grid_io_bottom_0_top_width_0_height_0__pin_1_upper[0]),
		.ccff_head(grid_io_bottom_0_ccff_tail[0]),
		.chany_top_out(sb_0__0__0_chany_top_out[0:19]),
		.chanx_right_out(sb_0__0__0_chanx_right_out[0:19]),
		.ccff_tail(ccff_tail[0]));

	sb_0__1_ sb_0__1_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_0__1__1_chany_bottom_out[0:19]),
		.top_left_grid_pin_1_(grid_io_left_1_right_width_0_height_0__pin_1_lower[0]),
		.chanx_right_in(cbx_1__1__0_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_1_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_1_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_1_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_1_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_1_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_1_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_1_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_1_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_0__1__0_chany_top_out[0:19]),
		.bottom_left_grid_pin_1_(grid_io_left_0_right_width_0_height_0__pin_1_upper[0]),
		.ccff_head(cbx_1__1__0_ccff_tail[0]),
		.chany_top_out(sb_0__1__0_chany_top_out[0:19]),
		.chanx_right_out(sb_0__1__0_chanx_right_out[0:19]),
		.chany_bottom_out(sb_0__1__0_chany_bottom_out[0:19]),
		.ccff_tail(sb_0__1__0_ccff_tail[0]));

	sb_0__1_ sb_0__2_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_0__1__2_chany_bottom_out[0:19]),
		.top_left_grid_pin_1_(grid_io_left_2_right_width_0_height_0__pin_1_lower[0]),
		.chanx_right_in(cbx_1__1__1_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_2_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_2_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_2_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_2_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_2_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_2_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_2_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_2_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_0__1__1_chany_top_out[0:19]),
		.bottom_left_grid_pin_1_(grid_io_left_1_right_width_0_height_0__pin_1_upper[0]),
		.ccff_head(cbx_1__1__1_ccff_tail[0]),
		.chany_top_out(sb_0__1__1_chany_top_out[0:19]),
		.chanx_right_out(sb_0__1__1_chanx_right_out[0:19]),
		.chany_bottom_out(sb_0__1__1_chany_bottom_out[0:19]),
		.ccff_tail(sb_0__1__1_ccff_tail[0]));

	sb_0__1_ sb_0__3_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_0__1__3_chany_bottom_out[0:19]),
		.top_left_grid_pin_1_(grid_io_left_3_right_width_0_height_0__pin_1_lower[0]),
		.chanx_right_in(cbx_1__1__2_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_3_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_3_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_3_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_3_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_3_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_3_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_3_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_3_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_0__1__2_chany_top_out[0:19]),
		.bottom_left_grid_pin_1_(grid_io_left_2_right_width_0_height_0__pin_1_upper[0]),
		.ccff_head(cbx_1__1__2_ccff_tail[0]),
		.chany_top_out(sb_0__1__2_chany_top_out[0:19]),
		.chanx_right_out(sb_0__1__2_chanx_right_out[0:19]),
		.chany_bottom_out(sb_0__1__2_chany_bottom_out[0:19]),
		.ccff_tail(sb_0__1__2_ccff_tail[0]));

	sb_0__1_ sb_0__4_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_0__1__4_chany_bottom_out[0:19]),
		.top_left_grid_pin_1_(grid_io_left_4_right_width_0_height_0__pin_1_lower[0]),
		.chanx_right_in(cbx_1__1__3_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_4_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_4_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_4_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_4_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_4_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_4_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_4_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_4_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_0__1__3_chany_top_out[0:19]),
		.bottom_left_grid_pin_1_(grid_io_left_3_right_width_0_height_0__pin_1_upper[0]),
		.ccff_head(cbx_1__1__3_ccff_tail[0]),
		.chany_top_out(sb_0__1__3_chany_top_out[0:19]),
		.chanx_right_out(sb_0__1__3_chanx_right_out[0:19]),
		.chany_bottom_out(sb_0__1__3_chany_bottom_out[0:19]),
		.ccff_tail(sb_0__1__3_ccff_tail[0]));

	sb_0__1_ sb_0__5_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_0__1__5_chany_bottom_out[0:19]),
		.top_left_grid_pin_1_(grid_io_left_5_right_width_0_height_0__pin_1_lower[0]),
		.chanx_right_in(cbx_1__1__4_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_5_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_5_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_5_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_5_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_5_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_5_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_5_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_5_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_0__1__4_chany_top_out[0:19]),
		.bottom_left_grid_pin_1_(grid_io_left_4_right_width_0_height_0__pin_1_upper[0]),
		.ccff_head(cbx_1__1__4_ccff_tail[0]),
		.chany_top_out(sb_0__1__4_chany_top_out[0:19]),
		.chanx_right_out(sb_0__1__4_chanx_right_out[0:19]),
		.chany_bottom_out(sb_0__1__4_chany_bottom_out[0:19]),
		.ccff_tail(sb_0__1__4_ccff_tail[0]));

	sb_0__1_ sb_0__6_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_0__1__6_chany_bottom_out[0:19]),
		.top_left_grid_pin_1_(grid_io_left_6_right_width_0_height_0__pin_1_lower[0]),
		.chanx_right_in(cbx_1__1__5_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_6_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_6_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_6_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_6_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_6_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_6_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_6_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_6_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_0__1__5_chany_top_out[0:19]),
		.bottom_left_grid_pin_1_(grid_io_left_5_right_width_0_height_0__pin_1_upper[0]),
		.ccff_head(cbx_1__1__5_ccff_tail[0]),
		.chany_top_out(sb_0__1__5_chany_top_out[0:19]),
		.chanx_right_out(sb_0__1__5_chanx_right_out[0:19]),
		.chany_bottom_out(sb_0__1__5_chany_bottom_out[0:19]),
		.ccff_tail(sb_0__1__5_ccff_tail[0]));

	sb_0__1_ sb_0__7_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_0__1__7_chany_bottom_out[0:19]),
		.top_left_grid_pin_1_(grid_io_left_7_right_width_0_height_0__pin_1_lower[0]),
		.chanx_right_in(cbx_1__1__6_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_7_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_7_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_7_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_7_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_7_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_7_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_7_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_7_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_0__1__6_chany_top_out[0:19]),
		.bottom_left_grid_pin_1_(grid_io_left_6_right_width_0_height_0__pin_1_upper[0]),
		.ccff_head(cbx_1__1__6_ccff_tail[0]),
		.chany_top_out(sb_0__1__6_chany_top_out[0:19]),
		.chanx_right_out(sb_0__1__6_chanx_right_out[0:19]),
		.chany_bottom_out(sb_0__1__6_chany_bottom_out[0:19]),
		.ccff_tail(sb_0__1__6_ccff_tail[0]));

	sb_0__1_ sb_0__8_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_0__1__8_chany_bottom_out[0:19]),
		.top_left_grid_pin_1_(grid_io_left_8_right_width_0_height_0__pin_1_lower[0]),
		.chanx_right_in(cbx_1__1__7_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_8_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_8_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_8_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_8_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_8_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_8_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_8_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_8_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_0__1__7_chany_top_out[0:19]),
		.bottom_left_grid_pin_1_(grid_io_left_7_right_width_0_height_0__pin_1_upper[0]),
		.ccff_head(cbx_1__1__7_ccff_tail[0]),
		.chany_top_out(sb_0__1__7_chany_top_out[0:19]),
		.chanx_right_out(sb_0__1__7_chanx_right_out[0:19]),
		.chany_bottom_out(sb_0__1__7_chany_bottom_out[0:19]),
		.ccff_tail(sb_0__1__7_ccff_tail[0]));

	sb_0__1_ sb_0__9_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_0__1__9_chany_bottom_out[0:19]),
		.top_left_grid_pin_1_(grid_io_left_9_right_width_0_height_0__pin_1_lower[0]),
		.chanx_right_in(cbx_1__1__8_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_9_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_9_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_9_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_9_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_9_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_9_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_9_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_9_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_0__1__8_chany_top_out[0:19]),
		.bottom_left_grid_pin_1_(grid_io_left_8_right_width_0_height_0__pin_1_upper[0]),
		.ccff_head(cbx_1__1__8_ccff_tail[0]),
		.chany_top_out(sb_0__1__8_chany_top_out[0:19]),
		.chanx_right_out(sb_0__1__8_chanx_right_out[0:19]),
		.chany_bottom_out(sb_0__1__8_chany_bottom_out[0:19]),
		.ccff_tail(sb_0__1__8_ccff_tail[0]));

	sb_0__1_ sb_0__10_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_0__1__10_chany_bottom_out[0:19]),
		.top_left_grid_pin_1_(grid_io_left_10_right_width_0_height_0__pin_1_lower[0]),
		.chanx_right_in(cbx_1__1__9_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_10_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_10_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_10_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_10_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_10_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_10_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_10_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_10_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_0__1__9_chany_top_out[0:19]),
		.bottom_left_grid_pin_1_(grid_io_left_9_right_width_0_height_0__pin_1_upper[0]),
		.ccff_head(cbx_1__1__9_ccff_tail[0]),
		.chany_top_out(sb_0__1__9_chany_top_out[0:19]),
		.chanx_right_out(sb_0__1__9_chanx_right_out[0:19]),
		.chany_bottom_out(sb_0__1__9_chany_bottom_out[0:19]),
		.ccff_tail(sb_0__1__9_ccff_tail[0]));

	sb_0__1_ sb_0__11_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_0__1__11_chany_bottom_out[0:19]),
		.top_left_grid_pin_1_(grid_io_left_11_right_width_0_height_0__pin_1_lower[0]),
		.chanx_right_in(cbx_1__1__10_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_11_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_11_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_11_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_11_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_11_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_11_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_11_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_11_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_0__1__10_chany_top_out[0:19]),
		.bottom_left_grid_pin_1_(grid_io_left_10_right_width_0_height_0__pin_1_upper[0]),
		.ccff_head(cbx_1__1__10_ccff_tail[0]),
		.chany_top_out(sb_0__1__10_chany_top_out[0:19]),
		.chanx_right_out(sb_0__1__10_chanx_right_out[0:19]),
		.chany_bottom_out(sb_0__1__10_chany_bottom_out[0:19]),
		.ccff_tail(sb_0__1__10_ccff_tail[0]));

	sb_0__2_ sb_0__12_ (
		.prog_clk(prog_clk[0]),
		.chanx_right_in(cbx_1__12__0_chanx_left_out[0:19]),
		.right_top_grid_pin_1_(grid_io_top_0_bottom_width_0_height_0__pin_1_upper[0]),
		.chany_bottom_in(cby_0__1__11_chany_top_out[0:19]),
		.bottom_left_grid_pin_1_(grid_io_left_11_right_width_0_height_0__pin_1_upper[0]),
		.ccff_head(grid_io_top_0_ccff_tail[0]),
		.chanx_right_out(sb_0__12__0_chanx_right_out[0:19]),
		.chany_bottom_out(sb_0__12__0_chany_bottom_out[0:19]),
		.ccff_tail(sb_0__12__0_ccff_tail[0]));

	sb_1__0_ sb_1__0_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__0_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_0_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_0_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_0_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_0_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_0_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_0_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_0_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_0_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__0__1_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_12_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_12_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_12_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_12_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_12_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_12_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_12_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_12_bottom_width_0_height_0__pin_49_upper[0]),
		.right_bottom_grid_pin_1_(grid_io_bottom_1_top_width_0_height_0__pin_1_upper[0]),
		.chanx_left_in(cbx_1__0__0_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_0_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_0_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_0_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_0_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_0_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_0_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_0_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_0_bottom_width_0_height_0__pin_49_lower[0]),
		.left_bottom_grid_pin_1_(grid_io_bottom_0_top_width_0_height_0__pin_1_lower[0]),
		.ccff_head(grid_io_bottom_1_ccff_tail[0]),
		.chany_top_out(sb_1__0__0_chany_top_out[0:19]),
		.chanx_right_out(sb_1__0__0_chanx_right_out[0:19]),
		.chanx_left_out(sb_1__0__0_chanx_left_out[0:19]),
		.ccff_tail(sb_1__0__0_ccff_tail[0]));

	sb_1__0_ sb_2__0_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__12_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_12_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_12_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_12_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_12_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_12_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_12_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_12_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_12_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__0__2_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_24_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_24_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_24_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_24_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_24_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_24_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_24_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_24_bottom_width_0_height_0__pin_49_upper[0]),
		.right_bottom_grid_pin_1_(grid_io_bottom_2_top_width_0_height_0__pin_1_upper[0]),
		.chanx_left_in(cbx_1__0__1_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_12_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_12_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_12_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_12_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_12_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_12_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_12_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_12_bottom_width_0_height_0__pin_49_lower[0]),
		.left_bottom_grid_pin_1_(grid_io_bottom_1_top_width_0_height_0__pin_1_lower[0]),
		.ccff_head(grid_io_bottom_2_ccff_tail[0]),
		.chany_top_out(sb_1__0__1_chany_top_out[0:19]),
		.chanx_right_out(sb_1__0__1_chanx_right_out[0:19]),
		.chanx_left_out(sb_1__0__1_chanx_left_out[0:19]),
		.ccff_tail(sb_1__0__1_ccff_tail[0]));

	sb_1__0_ sb_3__0_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__24_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_24_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_24_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_24_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_24_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_24_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_24_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_24_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_24_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__0__3_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_36_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_36_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_36_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_36_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_36_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_36_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_36_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_36_bottom_width_0_height_0__pin_49_upper[0]),
		.right_bottom_grid_pin_1_(grid_io_bottom_3_top_width_0_height_0__pin_1_upper[0]),
		.chanx_left_in(cbx_1__0__2_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_24_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_24_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_24_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_24_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_24_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_24_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_24_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_24_bottom_width_0_height_0__pin_49_lower[0]),
		.left_bottom_grid_pin_1_(grid_io_bottom_2_top_width_0_height_0__pin_1_lower[0]),
		.ccff_head(grid_io_bottom_3_ccff_tail[0]),
		.chany_top_out(sb_1__0__2_chany_top_out[0:19]),
		.chanx_right_out(sb_1__0__2_chanx_right_out[0:19]),
		.chanx_left_out(sb_1__0__2_chanx_left_out[0:19]),
		.ccff_tail(sb_1__0__2_ccff_tail[0]));

	sb_1__0_ sb_4__0_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__36_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_36_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_36_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_36_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_36_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_36_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_36_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_36_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_36_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__0__4_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_48_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_48_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_48_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_48_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_48_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_48_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_48_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_48_bottom_width_0_height_0__pin_49_upper[0]),
		.right_bottom_grid_pin_1_(grid_io_bottom_4_top_width_0_height_0__pin_1_upper[0]),
		.chanx_left_in(cbx_1__0__3_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_36_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_36_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_36_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_36_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_36_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_36_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_36_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_36_bottom_width_0_height_0__pin_49_lower[0]),
		.left_bottom_grid_pin_1_(grid_io_bottom_3_top_width_0_height_0__pin_1_lower[0]),
		.ccff_head(grid_io_bottom_4_ccff_tail[0]),
		.chany_top_out(sb_1__0__3_chany_top_out[0:19]),
		.chanx_right_out(sb_1__0__3_chanx_right_out[0:19]),
		.chanx_left_out(sb_1__0__3_chanx_left_out[0:19]),
		.ccff_tail(sb_1__0__3_ccff_tail[0]));

	sb_1__0_ sb_5__0_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__48_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_48_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_48_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_48_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_48_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_48_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_48_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_48_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_48_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__0__5_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_60_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_60_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_60_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_60_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_60_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_60_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_60_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_60_bottom_width_0_height_0__pin_49_upper[0]),
		.right_bottom_grid_pin_1_(grid_io_bottom_5_top_width_0_height_0__pin_1_upper[0]),
		.chanx_left_in(cbx_1__0__4_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_48_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_48_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_48_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_48_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_48_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_48_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_48_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_48_bottom_width_0_height_0__pin_49_lower[0]),
		.left_bottom_grid_pin_1_(grid_io_bottom_4_top_width_0_height_0__pin_1_lower[0]),
		.ccff_head(grid_io_bottom_5_ccff_tail[0]),
		.chany_top_out(sb_1__0__4_chany_top_out[0:19]),
		.chanx_right_out(sb_1__0__4_chanx_right_out[0:19]),
		.chanx_left_out(sb_1__0__4_chanx_left_out[0:19]),
		.ccff_tail(sb_1__0__4_ccff_tail[0]));

	sb_1__0_ sb_6__0_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__60_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_60_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_60_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_60_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_60_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_60_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_60_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_60_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_60_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__0__6_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_72_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_72_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_72_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_72_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_72_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_72_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_72_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_72_bottom_width_0_height_0__pin_49_upper[0]),
		.right_bottom_grid_pin_1_(grid_io_bottom_6_top_width_0_height_0__pin_1_upper[0]),
		.chanx_left_in(cbx_1__0__5_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_60_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_60_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_60_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_60_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_60_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_60_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_60_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_60_bottom_width_0_height_0__pin_49_lower[0]),
		.left_bottom_grid_pin_1_(grid_io_bottom_5_top_width_0_height_0__pin_1_lower[0]),
		.ccff_head(grid_io_bottom_6_ccff_tail[0]),
		.chany_top_out(sb_1__0__5_chany_top_out[0:19]),
		.chanx_right_out(sb_1__0__5_chanx_right_out[0:19]),
		.chanx_left_out(sb_1__0__5_chanx_left_out[0:19]),
		.ccff_tail(sb_1__0__5_ccff_tail[0]));

	sb_1__0_ sb_7__0_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__72_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_72_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_72_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_72_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_72_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_72_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_72_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_72_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_72_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__0__7_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_84_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_84_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_84_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_84_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_84_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_84_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_84_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_84_bottom_width_0_height_0__pin_49_upper[0]),
		.right_bottom_grid_pin_1_(grid_io_bottom_7_top_width_0_height_0__pin_1_upper[0]),
		.chanx_left_in(cbx_1__0__6_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_72_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_72_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_72_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_72_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_72_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_72_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_72_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_72_bottom_width_0_height_0__pin_49_lower[0]),
		.left_bottom_grid_pin_1_(grid_io_bottom_6_top_width_0_height_0__pin_1_lower[0]),
		.ccff_head(grid_io_bottom_7_ccff_tail[0]),
		.chany_top_out(sb_1__0__6_chany_top_out[0:19]),
		.chanx_right_out(sb_1__0__6_chanx_right_out[0:19]),
		.chanx_left_out(sb_1__0__6_chanx_left_out[0:19]),
		.ccff_tail(sb_1__0__6_ccff_tail[0]));

	sb_1__0_ sb_8__0_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__84_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_84_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_84_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_84_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_84_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_84_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_84_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_84_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_84_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__0__8_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_96_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_96_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_96_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_96_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_96_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_96_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_96_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_96_bottom_width_0_height_0__pin_49_upper[0]),
		.right_bottom_grid_pin_1_(grid_io_bottom_8_top_width_0_height_0__pin_1_upper[0]),
		.chanx_left_in(cbx_1__0__7_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_84_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_84_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_84_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_84_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_84_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_84_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_84_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_84_bottom_width_0_height_0__pin_49_lower[0]),
		.left_bottom_grid_pin_1_(grid_io_bottom_7_top_width_0_height_0__pin_1_lower[0]),
		.ccff_head(grid_io_bottom_8_ccff_tail[0]),
		.chany_top_out(sb_1__0__7_chany_top_out[0:19]),
		.chanx_right_out(sb_1__0__7_chanx_right_out[0:19]),
		.chanx_left_out(sb_1__0__7_chanx_left_out[0:19]),
		.ccff_tail(sb_1__0__7_ccff_tail[0]));

	sb_1__0_ sb_9__0_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__96_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_96_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_96_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_96_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_96_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_96_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_96_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_96_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_96_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__0__9_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_108_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_108_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_108_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_108_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_108_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_108_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_108_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_108_bottom_width_0_height_0__pin_49_upper[0]),
		.right_bottom_grid_pin_1_(grid_io_bottom_9_top_width_0_height_0__pin_1_upper[0]),
		.chanx_left_in(cbx_1__0__8_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_96_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_96_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_96_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_96_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_96_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_96_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_96_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_96_bottom_width_0_height_0__pin_49_lower[0]),
		.left_bottom_grid_pin_1_(grid_io_bottom_8_top_width_0_height_0__pin_1_lower[0]),
		.ccff_head(grid_io_bottom_9_ccff_tail[0]),
		.chany_top_out(sb_1__0__8_chany_top_out[0:19]),
		.chanx_right_out(sb_1__0__8_chanx_right_out[0:19]),
		.chanx_left_out(sb_1__0__8_chanx_left_out[0:19]),
		.ccff_tail(sb_1__0__8_ccff_tail[0]));

	sb_1__0_ sb_10__0_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__108_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_108_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_108_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_108_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_108_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_108_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_108_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_108_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_108_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__0__10_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_120_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_120_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_120_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_120_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_120_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_120_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_120_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_120_bottom_width_0_height_0__pin_49_upper[0]),
		.right_bottom_grid_pin_1_(grid_io_bottom_10_top_width_0_height_0__pin_1_upper[0]),
		.chanx_left_in(cbx_1__0__9_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_108_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_108_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_108_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_108_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_108_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_108_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_108_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_108_bottom_width_0_height_0__pin_49_lower[0]),
		.left_bottom_grid_pin_1_(grid_io_bottom_9_top_width_0_height_0__pin_1_lower[0]),
		.ccff_head(grid_io_bottom_10_ccff_tail[0]),
		.chany_top_out(sb_1__0__9_chany_top_out[0:19]),
		.chanx_right_out(sb_1__0__9_chanx_right_out[0:19]),
		.chanx_left_out(sb_1__0__9_chanx_left_out[0:19]),
		.ccff_tail(sb_1__0__9_ccff_tail[0]));

	sb_1__0_ sb_11__0_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__120_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_120_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_120_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_120_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_120_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_120_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_120_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_120_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_120_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__0__11_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_132_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_132_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_132_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_132_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_132_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_132_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_132_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_132_bottom_width_0_height_0__pin_49_upper[0]),
		.right_bottom_grid_pin_1_(grid_io_bottom_11_top_width_0_height_0__pin_1_upper[0]),
		.chanx_left_in(cbx_1__0__10_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_120_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_120_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_120_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_120_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_120_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_120_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_120_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_120_bottom_width_0_height_0__pin_49_lower[0]),
		.left_bottom_grid_pin_1_(grid_io_bottom_10_top_width_0_height_0__pin_1_lower[0]),
		.ccff_head(grid_io_bottom_11_ccff_tail[0]),
		.chany_top_out(sb_1__0__10_chany_top_out[0:19]),
		.chanx_right_out(sb_1__0__10_chanx_right_out[0:19]),
		.chanx_left_out(sb_1__0__10_chanx_left_out[0:19]),
		.ccff_tail(sb_1__0__10_ccff_tail[0]));

	sb_1__1_ sb_1__1_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__1_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_1_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_1_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_1_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_1_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_1_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_1_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_1_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_1_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__1__11_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_13_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_13_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_13_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_13_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_13_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_13_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_13_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_13_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_1__1__0_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_0_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_0_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_0_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_0_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_0_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_0_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_0_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_0_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__0_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_1_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_1_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_1_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_1_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_1_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_1_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_1_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_1_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(cbx_1__1__11_ccff_tail[0]),
		.chany_top_out(sb_1__1__0_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__0_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__0_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__0_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__0_ccff_tail[0]));

	sb_1__1_ sb_1__2_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__2_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_2_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_2_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_2_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_2_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_2_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_2_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_2_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_2_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__1__12_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_14_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_14_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_14_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_14_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_14_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_14_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_14_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_14_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_1__1__1_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_1_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_1_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_1_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_1_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_1_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_1_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_1_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_1_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__1_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_2_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_2_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_2_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_2_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_2_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_2_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_2_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_2_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(cbx_1__1__12_ccff_tail[0]),
		.chany_top_out(sb_1__1__1_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__1_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__1_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__1_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__1_ccff_tail[0]));

	sb_1__1_ sb_1__3_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__3_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_3_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_3_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_3_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_3_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_3_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_3_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_3_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_3_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__1__13_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_15_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_15_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_15_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_15_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_15_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_15_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_15_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_15_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_1__1__2_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_2_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_2_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_2_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_2_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_2_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_2_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_2_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_2_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__2_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_3_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_3_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_3_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_3_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_3_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_3_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_3_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_3_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(cbx_1__1__13_ccff_tail[0]),
		.chany_top_out(sb_1__1__2_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__2_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__2_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__2_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__2_ccff_tail[0]));

	sb_1__1_ sb_1__4_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__4_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_4_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_4_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_4_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_4_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_4_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_4_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_4_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_4_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__1__14_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_16_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_16_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_16_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_16_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_16_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_16_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_16_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_16_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_1__1__3_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_3_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_3_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_3_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_3_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_3_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_3_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_3_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_3_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__3_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_4_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_4_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_4_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_4_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_4_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_4_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_4_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_4_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(cbx_1__1__14_ccff_tail[0]),
		.chany_top_out(sb_1__1__3_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__3_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__3_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__3_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__3_ccff_tail[0]));

	sb_1__1_ sb_1__5_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__5_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_5_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_5_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_5_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_5_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_5_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_5_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_5_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_5_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__1__15_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_17_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_17_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_17_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_17_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_17_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_17_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_17_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_17_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_1__1__4_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_4_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_4_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_4_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_4_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_4_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_4_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_4_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_4_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__4_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_5_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_5_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_5_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_5_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_5_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_5_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_5_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_5_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(cbx_1__1__15_ccff_tail[0]),
		.chany_top_out(sb_1__1__4_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__4_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__4_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__4_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__4_ccff_tail[0]));

	sb_1__1_ sb_1__6_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__6_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_6_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_6_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_6_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_6_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_6_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_6_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_6_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_6_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__1__16_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_18_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_18_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_18_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_18_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_18_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_18_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_18_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_18_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_1__1__5_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_5_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_5_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_5_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_5_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_5_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_5_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_5_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_5_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__5_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_6_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_6_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_6_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_6_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_6_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_6_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_6_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_6_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(cbx_1__1__16_ccff_tail[0]),
		.chany_top_out(sb_1__1__5_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__5_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__5_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__5_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__5_ccff_tail[0]));

	sb_1__1_ sb_1__7_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__7_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_7_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_7_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_7_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_7_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_7_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_7_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_7_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_7_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__1__17_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_19_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_19_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_19_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_19_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_19_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_19_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_19_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_19_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_1__1__6_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_6_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_6_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_6_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_6_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_6_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_6_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_6_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_6_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__6_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_7_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_7_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_7_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_7_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_7_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_7_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_7_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_7_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(cbx_1__1__17_ccff_tail[0]),
		.chany_top_out(sb_1__1__6_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__6_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__6_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__6_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__6_ccff_tail[0]));

	sb_1__1_ sb_1__8_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__8_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_8_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_8_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_8_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_8_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_8_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_8_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_8_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_8_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__1__18_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_20_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_20_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_20_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_20_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_20_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_20_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_20_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_20_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_1__1__7_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_7_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_7_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_7_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_7_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_7_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_7_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_7_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_7_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__7_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_8_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_8_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_8_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_8_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_8_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_8_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_8_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_8_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(cbx_1__1__18_ccff_tail[0]),
		.chany_top_out(sb_1__1__7_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__7_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__7_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__7_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__7_ccff_tail[0]));

	sb_1__1_ sb_1__9_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__9_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_9_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_9_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_9_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_9_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_9_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_9_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_9_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_9_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__1__19_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_21_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_21_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_21_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_21_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_21_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_21_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_21_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_21_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_1__1__8_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_8_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_8_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_8_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_8_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_8_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_8_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_8_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_8_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__8_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_9_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_9_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_9_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_9_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_9_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_9_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_9_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_9_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(cbx_1__1__19_ccff_tail[0]),
		.chany_top_out(sb_1__1__8_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__8_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__8_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__8_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__8_ccff_tail[0]));

	sb_1__1_ sb_1__10_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__10_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_10_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_10_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_10_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_10_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_10_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_10_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_10_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_10_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__1__20_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_22_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_22_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_22_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_22_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_22_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_22_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_22_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_22_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_1__1__9_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_9_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_9_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_9_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_9_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_9_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_9_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_9_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_9_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__9_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_10_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_10_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_10_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_10_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_10_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_10_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_10_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_10_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(cbx_1__1__20_ccff_tail[0]),
		.chany_top_out(sb_1__1__9_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__9_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__9_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__9_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__9_ccff_tail[0]));

	sb_1__1_ sb_1__11_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__11_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_11_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_11_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_11_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_11_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_11_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_11_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_11_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_11_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__1__21_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_23_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_23_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_23_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_23_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_23_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_23_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_23_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_23_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_1__1__10_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_10_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_10_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_10_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_10_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_10_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_10_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_10_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_10_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__10_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_11_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_11_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_11_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_11_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_11_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_11_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_11_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_11_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(cbx_1__1__21_ccff_tail[0]),
		.chany_top_out(sb_1__1__10_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__10_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__10_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__10_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__10_ccff_tail[0]));

	sb_1__1_ sb_2__1_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__13_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_13_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_13_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_13_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_13_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_13_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_13_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_13_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_13_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__1__22_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_25_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_25_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_25_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_25_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_25_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_25_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_25_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_25_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_1__1__12_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_12_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_12_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_12_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_12_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_12_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_12_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_12_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_12_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__11_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_13_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_13_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_13_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_13_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_13_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_13_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_13_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_13_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(cbx_1__1__22_ccff_tail[0]),
		.chany_top_out(sb_1__1__11_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__11_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__11_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__11_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__11_ccff_tail[0]));

	sb_1__1_ sb_2__2_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__14_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_14_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_14_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_14_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_14_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_14_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_14_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_14_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_14_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__1__23_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_26_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_26_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_26_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_26_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_26_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_26_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_26_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_26_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_1__1__13_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_13_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_13_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_13_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_13_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_13_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_13_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_13_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_13_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__12_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_14_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_14_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_14_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_14_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_14_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_14_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_14_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_14_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(cbx_1__1__23_ccff_tail[0]),
		.chany_top_out(sb_1__1__12_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__12_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__12_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__12_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__12_ccff_tail[0]));

	sb_1__1_ sb_2__3_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__15_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_15_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_15_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_15_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_15_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_15_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_15_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_15_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_15_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__1__24_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_27_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_27_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_27_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_27_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_27_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_27_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_27_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_27_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_1__1__14_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_14_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_14_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_14_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_14_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_14_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_14_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_14_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_14_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__13_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_15_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_15_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_15_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_15_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_15_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_15_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_15_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_15_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(cbx_1__1__24_ccff_tail[0]),
		.chany_top_out(sb_1__1__13_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__13_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__13_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__13_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__13_ccff_tail[0]));

	sb_1__1_ sb_2__4_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__16_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_16_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_16_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_16_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_16_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_16_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_16_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_16_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_16_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__1__25_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_28_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_28_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_28_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_28_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_28_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_28_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_28_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_28_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_1__1__15_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_15_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_15_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_15_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_15_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_15_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_15_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_15_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_15_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__14_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_16_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_16_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_16_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_16_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_16_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_16_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_16_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_16_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(cbx_1__1__25_ccff_tail[0]),
		.chany_top_out(sb_1__1__14_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__14_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__14_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__14_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__14_ccff_tail[0]));

	sb_1__1_ sb_2__5_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__17_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_17_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_17_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_17_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_17_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_17_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_17_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_17_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_17_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__1__26_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_29_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_29_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_29_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_29_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_29_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_29_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_29_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_29_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_1__1__16_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_16_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_16_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_16_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_16_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_16_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_16_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_16_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_16_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__15_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_17_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_17_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_17_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_17_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_17_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_17_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_17_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_17_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(cbx_1__1__26_ccff_tail[0]),
		.chany_top_out(sb_1__1__15_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__15_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__15_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__15_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__15_ccff_tail[0]));

	sb_1__1_ sb_2__6_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__18_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_18_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_18_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_18_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_18_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_18_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_18_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_18_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_18_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__1__27_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_30_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_30_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_30_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_30_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_30_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_30_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_30_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_30_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_1__1__17_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_17_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_17_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_17_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_17_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_17_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_17_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_17_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_17_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__16_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_18_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_18_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_18_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_18_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_18_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_18_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_18_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_18_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(cbx_1__1__27_ccff_tail[0]),
		.chany_top_out(sb_1__1__16_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__16_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__16_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__16_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__16_ccff_tail[0]));

	sb_1__1_ sb_2__7_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__19_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_19_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_19_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_19_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_19_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_19_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_19_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_19_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_19_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__1__28_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_31_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_31_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_31_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_31_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_31_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_31_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_31_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_31_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_1__1__18_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_18_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_18_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_18_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_18_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_18_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_18_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_18_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_18_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__17_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_19_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_19_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_19_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_19_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_19_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_19_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_19_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_19_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(cbx_1__1__28_ccff_tail[0]),
		.chany_top_out(sb_1__1__17_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__17_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__17_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__17_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__17_ccff_tail[0]));

	sb_1__1_ sb_2__8_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__20_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_20_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_20_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_20_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_20_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_20_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_20_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_20_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_20_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__1__29_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_32_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_32_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_32_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_32_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_32_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_32_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_32_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_32_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_1__1__19_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_19_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_19_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_19_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_19_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_19_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_19_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_19_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_19_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__18_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_20_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_20_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_20_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_20_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_20_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_20_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_20_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_20_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(cbx_1__1__29_ccff_tail[0]),
		.chany_top_out(sb_1__1__18_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__18_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__18_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__18_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__18_ccff_tail[0]));

	sb_1__1_ sb_2__9_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__21_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_21_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_21_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_21_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_21_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_21_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_21_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_21_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_21_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__1__30_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_33_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_33_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_33_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_33_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_33_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_33_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_33_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_33_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_1__1__20_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_20_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_20_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_20_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_20_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_20_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_20_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_20_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_20_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__19_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_21_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_21_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_21_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_21_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_21_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_21_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_21_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_21_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(cbx_1__1__30_ccff_tail[0]),
		.chany_top_out(sb_1__1__19_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__19_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__19_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__19_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__19_ccff_tail[0]));

	sb_1__1_ sb_2__10_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__22_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_22_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_22_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_22_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_22_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_22_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_22_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_22_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_22_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__1__31_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_34_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_34_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_34_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_34_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_34_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_34_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_34_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_34_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_1__1__21_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_21_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_21_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_21_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_21_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_21_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_21_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_21_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_21_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__20_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_22_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_22_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_22_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_22_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_22_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_22_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_22_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_22_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(cbx_1__1__31_ccff_tail[0]),
		.chany_top_out(sb_1__1__20_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__20_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__20_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__20_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__20_ccff_tail[0]));

	sb_1__1_ sb_2__11_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__23_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_23_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_23_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_23_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_23_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_23_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_23_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_23_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_23_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__1__32_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_35_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_35_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_35_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_35_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_35_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_35_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_35_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_35_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_1__1__22_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_22_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_22_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_22_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_22_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_22_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_22_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_22_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_22_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__21_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_23_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_23_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_23_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_23_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_23_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_23_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_23_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_23_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(cbx_1__1__32_ccff_tail[0]),
		.chany_top_out(sb_1__1__21_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__21_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__21_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__21_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__21_ccff_tail[0]));

	sb_1__1_ sb_3__1_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__25_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_25_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_25_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_25_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_25_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_25_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_25_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_25_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_25_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__1__33_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_37_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_37_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_37_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_37_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_37_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_37_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_37_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_37_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_1__1__24_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_24_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_24_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_24_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_24_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_24_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_24_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_24_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_24_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__22_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_25_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_25_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_25_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_25_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_25_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_25_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_25_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_25_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(cbx_1__1__33_ccff_tail[0]),
		.chany_top_out(sb_1__1__22_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__22_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__22_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__22_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__22_ccff_tail[0]));

	sb_1__1_ sb_3__2_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__26_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_26_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_26_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_26_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_26_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_26_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_26_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_26_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_26_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__1__34_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_38_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_38_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_38_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_38_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_38_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_38_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_38_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_38_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_1__1__25_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_25_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_25_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_25_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_25_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_25_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_25_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_25_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_25_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__23_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_26_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_26_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_26_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_26_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_26_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_26_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_26_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_26_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(cbx_1__1__34_ccff_tail[0]),
		.chany_top_out(sb_1__1__23_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__23_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__23_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__23_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__23_ccff_tail[0]));

	sb_1__1_ sb_3__3_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__27_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_27_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_27_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_27_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_27_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_27_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_27_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_27_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_27_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__1__35_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_39_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_39_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_39_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_39_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_39_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_39_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_39_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_39_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_1__1__26_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_26_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_26_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_26_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_26_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_26_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_26_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_26_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_26_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__24_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_27_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_27_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_27_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_27_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_27_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_27_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_27_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_27_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(cbx_1__1__35_ccff_tail[0]),
		.chany_top_out(sb_1__1__24_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__24_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__24_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__24_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__24_ccff_tail[0]));

	sb_1__1_ sb_3__4_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__28_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_28_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_28_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_28_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_28_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_28_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_28_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_28_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_28_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__1__36_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_40_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_40_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_40_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_40_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_40_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_40_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_40_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_40_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_1__1__27_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_27_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_27_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_27_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_27_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_27_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_27_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_27_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_27_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__25_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_28_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_28_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_28_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_28_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_28_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_28_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_28_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_28_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(cbx_1__1__36_ccff_tail[0]),
		.chany_top_out(sb_1__1__25_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__25_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__25_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__25_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__25_ccff_tail[0]));

	sb_1__1_ sb_3__5_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__29_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_29_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_29_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_29_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_29_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_29_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_29_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_29_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_29_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__1__37_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_41_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_41_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_41_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_41_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_41_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_41_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_41_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_41_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_1__1__28_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_28_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_28_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_28_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_28_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_28_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_28_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_28_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_28_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__26_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_29_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_29_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_29_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_29_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_29_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_29_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_29_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_29_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(cbx_1__1__37_ccff_tail[0]),
		.chany_top_out(sb_1__1__26_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__26_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__26_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__26_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__26_ccff_tail[0]));

	sb_1__1_ sb_3__6_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__30_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_30_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_30_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_30_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_30_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_30_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_30_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_30_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_30_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__1__38_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_42_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_42_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_42_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_42_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_42_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_42_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_42_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_42_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_1__1__29_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_29_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_29_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_29_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_29_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_29_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_29_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_29_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_29_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__27_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_30_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_30_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_30_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_30_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_30_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_30_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_30_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_30_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(cbx_1__1__38_ccff_tail[0]),
		.chany_top_out(sb_1__1__27_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__27_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__27_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__27_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__27_ccff_tail[0]));

	sb_1__1_ sb_3__7_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__31_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_31_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_31_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_31_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_31_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_31_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_31_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_31_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_31_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__1__39_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_43_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_43_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_43_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_43_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_43_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_43_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_43_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_43_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_1__1__30_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_30_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_30_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_30_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_30_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_30_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_30_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_30_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_30_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__28_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_31_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_31_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_31_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_31_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_31_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_31_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_31_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_31_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(cbx_1__1__39_ccff_tail[0]),
		.chany_top_out(sb_1__1__28_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__28_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__28_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__28_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__28_ccff_tail[0]));

	sb_1__1_ sb_3__8_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__32_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_32_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_32_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_32_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_32_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_32_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_32_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_32_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_32_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__1__40_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_44_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_44_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_44_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_44_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_44_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_44_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_44_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_44_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_1__1__31_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_31_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_31_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_31_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_31_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_31_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_31_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_31_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_31_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__29_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_32_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_32_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_32_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_32_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_32_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_32_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_32_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_32_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(cbx_1__1__40_ccff_tail[0]),
		.chany_top_out(sb_1__1__29_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__29_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__29_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__29_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__29_ccff_tail[0]));

	sb_1__1_ sb_3__9_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__33_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_33_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_33_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_33_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_33_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_33_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_33_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_33_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_33_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__1__41_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_45_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_45_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_45_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_45_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_45_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_45_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_45_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_45_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_1__1__32_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_32_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_32_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_32_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_32_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_32_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_32_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_32_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_32_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__30_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_33_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_33_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_33_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_33_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_33_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_33_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_33_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_33_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(cbx_1__1__41_ccff_tail[0]),
		.chany_top_out(sb_1__1__30_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__30_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__30_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__30_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__30_ccff_tail[0]));

	sb_1__1_ sb_3__10_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__34_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_34_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_34_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_34_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_34_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_34_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_34_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_34_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_34_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__1__42_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_46_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_46_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_46_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_46_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_46_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_46_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_46_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_46_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_1__1__33_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_33_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_33_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_33_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_33_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_33_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_33_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_33_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_33_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__31_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_34_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_34_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_34_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_34_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_34_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_34_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_34_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_34_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(cbx_1__1__42_ccff_tail[0]),
		.chany_top_out(sb_1__1__31_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__31_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__31_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__31_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__31_ccff_tail[0]));

	sb_1__1_ sb_3__11_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__35_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_35_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_35_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_35_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_35_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_35_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_35_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_35_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_35_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__1__43_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_47_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_47_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_47_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_47_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_47_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_47_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_47_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_47_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_1__1__34_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_34_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_34_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_34_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_34_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_34_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_34_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_34_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_34_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__32_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_35_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_35_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_35_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_35_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_35_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_35_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_35_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_35_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(cbx_1__1__43_ccff_tail[0]),
		.chany_top_out(sb_1__1__32_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__32_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__32_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__32_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__32_ccff_tail[0]));

	sb_1__1_ sb_4__1_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__37_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_37_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_37_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_37_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_37_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_37_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_37_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_37_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_37_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__1__44_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_49_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_49_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_49_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_49_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_49_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_49_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_49_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_49_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_1__1__36_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_36_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_36_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_36_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_36_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_36_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_36_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_36_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_36_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__33_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_37_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_37_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_37_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_37_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_37_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_37_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_37_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_37_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(cbx_1__1__44_ccff_tail[0]),
		.chany_top_out(sb_1__1__33_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__33_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__33_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__33_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__33_ccff_tail[0]));

	sb_1__1_ sb_4__2_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__38_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_38_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_38_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_38_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_38_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_38_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_38_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_38_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_38_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__1__45_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_50_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_50_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_50_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_50_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_50_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_50_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_50_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_50_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_1__1__37_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_37_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_37_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_37_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_37_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_37_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_37_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_37_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_37_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__34_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_38_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_38_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_38_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_38_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_38_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_38_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_38_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_38_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(cbx_1__1__45_ccff_tail[0]),
		.chany_top_out(sb_1__1__34_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__34_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__34_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__34_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__34_ccff_tail[0]));

	sb_1__1_ sb_4__3_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__39_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_39_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_39_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_39_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_39_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_39_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_39_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_39_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_39_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__1__46_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_51_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_51_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_51_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_51_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_51_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_51_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_51_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_51_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_1__1__38_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_38_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_38_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_38_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_38_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_38_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_38_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_38_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_38_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__35_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_39_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_39_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_39_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_39_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_39_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_39_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_39_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_39_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(cbx_1__1__46_ccff_tail[0]),
		.chany_top_out(sb_1__1__35_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__35_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__35_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__35_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__35_ccff_tail[0]));

	sb_1__1_ sb_4__4_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__40_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_40_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_40_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_40_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_40_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_40_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_40_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_40_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_40_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__1__47_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_52_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_52_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_52_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_52_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_52_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_52_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_52_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_52_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_1__1__39_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_39_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_39_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_39_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_39_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_39_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_39_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_39_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_39_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__36_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_40_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_40_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_40_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_40_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_40_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_40_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_40_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_40_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(cbx_1__1__47_ccff_tail[0]),
		.chany_top_out(sb_1__1__36_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__36_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__36_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__36_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__36_ccff_tail[0]));

	sb_1__1_ sb_4__5_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__41_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_41_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_41_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_41_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_41_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_41_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_41_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_41_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_41_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__1__48_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_53_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_53_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_53_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_53_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_53_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_53_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_53_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_53_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_1__1__40_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_40_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_40_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_40_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_40_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_40_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_40_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_40_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_40_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__37_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_41_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_41_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_41_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_41_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_41_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_41_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_41_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_41_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(cbx_1__1__48_ccff_tail[0]),
		.chany_top_out(sb_1__1__37_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__37_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__37_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__37_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__37_ccff_tail[0]));

	sb_1__1_ sb_4__6_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__42_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_42_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_42_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_42_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_42_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_42_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_42_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_42_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_42_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__1__49_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_54_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_54_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_54_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_54_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_54_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_54_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_54_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_54_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_1__1__41_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_41_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_41_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_41_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_41_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_41_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_41_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_41_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_41_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__38_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_42_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_42_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_42_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_42_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_42_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_42_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_42_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_42_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(cbx_1__1__49_ccff_tail[0]),
		.chany_top_out(sb_1__1__38_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__38_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__38_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__38_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__38_ccff_tail[0]));

	sb_1__1_ sb_4__7_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__43_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_43_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_43_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_43_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_43_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_43_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_43_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_43_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_43_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__1__50_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_55_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_55_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_55_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_55_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_55_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_55_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_55_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_55_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_1__1__42_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_42_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_42_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_42_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_42_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_42_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_42_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_42_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_42_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__39_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_43_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_43_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_43_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_43_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_43_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_43_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_43_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_43_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(cbx_1__1__50_ccff_tail[0]),
		.chany_top_out(sb_1__1__39_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__39_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__39_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__39_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__39_ccff_tail[0]));

	sb_1__1_ sb_4__8_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__44_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_44_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_44_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_44_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_44_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_44_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_44_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_44_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_44_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__1__51_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_56_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_56_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_56_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_56_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_56_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_56_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_56_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_56_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_1__1__43_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_43_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_43_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_43_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_43_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_43_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_43_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_43_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_43_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__40_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_44_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_44_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_44_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_44_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_44_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_44_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_44_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_44_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(cbx_1__1__51_ccff_tail[0]),
		.chany_top_out(sb_1__1__40_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__40_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__40_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__40_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__40_ccff_tail[0]));

	sb_1__1_ sb_4__9_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__45_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_45_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_45_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_45_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_45_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_45_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_45_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_45_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_45_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__1__52_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_57_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_57_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_57_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_57_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_57_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_57_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_57_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_57_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_1__1__44_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_44_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_44_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_44_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_44_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_44_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_44_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_44_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_44_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__41_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_45_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_45_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_45_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_45_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_45_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_45_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_45_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_45_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(cbx_1__1__52_ccff_tail[0]),
		.chany_top_out(sb_1__1__41_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__41_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__41_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__41_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__41_ccff_tail[0]));

	sb_1__1_ sb_4__10_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__46_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_46_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_46_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_46_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_46_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_46_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_46_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_46_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_46_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__1__53_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_58_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_58_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_58_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_58_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_58_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_58_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_58_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_58_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_1__1__45_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_45_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_45_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_45_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_45_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_45_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_45_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_45_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_45_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__42_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_46_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_46_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_46_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_46_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_46_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_46_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_46_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_46_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(cbx_1__1__53_ccff_tail[0]),
		.chany_top_out(sb_1__1__42_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__42_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__42_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__42_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__42_ccff_tail[0]));

	sb_1__1_ sb_4__11_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__47_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_47_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_47_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_47_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_47_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_47_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_47_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_47_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_47_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__1__54_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_59_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_59_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_59_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_59_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_59_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_59_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_59_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_59_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_1__1__46_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_46_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_46_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_46_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_46_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_46_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_46_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_46_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_46_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__43_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_47_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_47_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_47_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_47_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_47_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_47_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_47_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_47_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(cbx_1__1__54_ccff_tail[0]),
		.chany_top_out(sb_1__1__43_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__43_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__43_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__43_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__43_ccff_tail[0]));

	sb_1__1_ sb_5__1_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__49_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_49_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_49_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_49_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_49_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_49_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_49_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_49_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_49_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__1__55_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_61_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_61_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_61_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_61_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_61_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_61_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_61_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_61_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_1__1__48_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_48_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_48_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_48_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_48_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_48_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_48_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_48_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_48_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__44_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_49_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_49_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_49_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_49_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_49_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_49_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_49_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_49_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(cbx_1__1__55_ccff_tail[0]),
		.chany_top_out(sb_1__1__44_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__44_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__44_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__44_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__44_ccff_tail[0]));

	sb_1__1_ sb_5__2_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__50_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_50_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_50_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_50_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_50_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_50_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_50_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_50_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_50_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__1__56_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_62_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_62_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_62_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_62_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_62_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_62_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_62_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_62_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_1__1__49_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_49_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_49_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_49_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_49_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_49_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_49_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_49_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_49_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__45_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_50_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_50_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_50_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_50_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_50_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_50_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_50_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_50_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(cbx_1__1__56_ccff_tail[0]),
		.chany_top_out(sb_1__1__45_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__45_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__45_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__45_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__45_ccff_tail[0]));

	sb_1__1_ sb_5__3_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__51_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_51_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_51_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_51_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_51_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_51_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_51_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_51_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_51_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__1__57_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_63_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_63_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_63_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_63_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_63_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_63_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_63_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_63_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_1__1__50_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_50_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_50_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_50_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_50_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_50_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_50_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_50_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_50_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__46_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_51_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_51_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_51_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_51_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_51_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_51_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_51_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_51_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(cbx_1__1__57_ccff_tail[0]),
		.chany_top_out(sb_1__1__46_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__46_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__46_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__46_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__46_ccff_tail[0]));

	sb_1__1_ sb_5__4_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__52_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_52_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_52_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_52_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_52_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_52_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_52_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_52_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_52_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__1__58_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_64_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_64_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_64_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_64_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_64_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_64_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_64_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_64_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_1__1__51_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_51_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_51_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_51_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_51_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_51_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_51_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_51_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_51_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__47_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_52_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_52_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_52_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_52_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_52_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_52_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_52_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_52_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(cbx_1__1__58_ccff_tail[0]),
		.chany_top_out(sb_1__1__47_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__47_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__47_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__47_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__47_ccff_tail[0]));

	sb_1__1_ sb_5__5_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__53_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_53_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_53_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_53_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_53_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_53_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_53_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_53_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_53_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__1__59_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_65_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_65_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_65_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_65_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_65_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_65_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_65_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_65_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_1__1__52_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_52_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_52_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_52_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_52_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_52_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_52_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_52_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_52_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__48_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_53_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_53_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_53_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_53_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_53_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_53_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_53_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_53_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(cbx_1__1__59_ccff_tail[0]),
		.chany_top_out(sb_1__1__48_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__48_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__48_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__48_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__48_ccff_tail[0]));

	sb_1__1_ sb_5__6_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__54_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_54_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_54_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_54_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_54_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_54_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_54_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_54_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_54_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__1__60_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_66_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_66_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_66_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_66_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_66_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_66_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_66_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_66_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_1__1__53_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_53_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_53_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_53_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_53_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_53_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_53_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_53_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_53_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__49_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_54_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_54_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_54_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_54_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_54_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_54_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_54_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_54_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(cbx_1__1__60_ccff_tail[0]),
		.chany_top_out(sb_1__1__49_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__49_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__49_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__49_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__49_ccff_tail[0]));

	sb_1__1_ sb_5__7_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__55_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_55_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_55_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_55_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_55_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_55_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_55_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_55_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_55_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__1__61_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_67_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_67_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_67_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_67_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_67_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_67_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_67_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_67_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_1__1__54_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_54_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_54_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_54_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_54_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_54_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_54_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_54_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_54_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__50_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_55_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_55_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_55_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_55_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_55_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_55_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_55_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_55_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(cbx_1__1__61_ccff_tail[0]),
		.chany_top_out(sb_1__1__50_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__50_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__50_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__50_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__50_ccff_tail[0]));

	sb_1__1_ sb_5__8_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__56_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_56_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_56_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_56_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_56_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_56_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_56_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_56_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_56_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__1__62_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_68_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_68_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_68_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_68_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_68_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_68_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_68_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_68_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_1__1__55_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_55_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_55_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_55_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_55_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_55_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_55_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_55_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_55_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__51_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_56_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_56_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_56_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_56_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_56_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_56_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_56_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_56_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(cbx_1__1__62_ccff_tail[0]),
		.chany_top_out(sb_1__1__51_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__51_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__51_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__51_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__51_ccff_tail[0]));

	sb_1__1_ sb_5__9_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__57_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_57_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_57_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_57_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_57_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_57_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_57_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_57_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_57_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__1__63_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_69_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_69_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_69_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_69_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_69_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_69_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_69_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_69_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_1__1__56_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_56_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_56_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_56_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_56_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_56_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_56_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_56_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_56_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__52_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_57_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_57_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_57_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_57_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_57_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_57_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_57_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_57_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(cbx_1__1__63_ccff_tail[0]),
		.chany_top_out(sb_1__1__52_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__52_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__52_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__52_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__52_ccff_tail[0]));

	sb_1__1_ sb_5__10_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__58_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_58_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_58_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_58_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_58_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_58_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_58_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_58_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_58_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__1__64_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_70_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_70_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_70_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_70_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_70_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_70_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_70_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_70_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_1__1__57_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_57_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_57_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_57_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_57_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_57_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_57_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_57_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_57_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__53_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_58_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_58_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_58_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_58_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_58_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_58_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_58_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_58_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(cbx_1__1__64_ccff_tail[0]),
		.chany_top_out(sb_1__1__53_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__53_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__53_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__53_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__53_ccff_tail[0]));

	sb_1__1_ sb_5__11_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__59_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_59_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_59_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_59_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_59_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_59_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_59_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_59_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_59_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__1__65_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_71_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_71_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_71_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_71_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_71_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_71_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_71_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_71_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_1__1__58_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_58_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_58_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_58_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_58_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_58_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_58_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_58_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_58_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__54_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_59_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_59_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_59_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_59_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_59_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_59_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_59_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_59_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(cbx_1__1__65_ccff_tail[0]),
		.chany_top_out(sb_1__1__54_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__54_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__54_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__54_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__54_ccff_tail[0]));

	sb_1__1_ sb_6__1_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__61_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_61_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_61_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_61_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_61_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_61_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_61_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_61_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_61_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__1__66_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_73_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_73_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_73_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_73_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_73_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_73_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_73_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_73_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_1__1__60_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_60_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_60_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_60_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_60_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_60_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_60_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_60_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_60_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__55_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_61_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_61_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_61_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_61_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_61_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_61_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_61_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_61_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(cbx_1__1__66_ccff_tail[0]),
		.chany_top_out(sb_1__1__55_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__55_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__55_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__55_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__55_ccff_tail[0]));

	sb_1__1_ sb_6__2_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__62_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_62_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_62_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_62_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_62_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_62_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_62_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_62_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_62_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__1__67_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_74_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_74_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_74_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_74_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_74_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_74_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_74_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_74_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_1__1__61_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_61_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_61_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_61_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_61_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_61_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_61_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_61_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_61_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__56_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_62_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_62_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_62_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_62_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_62_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_62_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_62_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_62_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(cbx_1__1__67_ccff_tail[0]),
		.chany_top_out(sb_1__1__56_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__56_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__56_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__56_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__56_ccff_tail[0]));

	sb_1__1_ sb_6__3_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__63_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_63_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_63_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_63_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_63_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_63_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_63_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_63_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_63_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__1__68_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_75_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_75_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_75_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_75_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_75_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_75_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_75_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_75_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_1__1__62_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_62_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_62_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_62_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_62_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_62_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_62_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_62_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_62_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__57_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_63_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_63_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_63_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_63_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_63_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_63_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_63_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_63_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(cbx_1__1__68_ccff_tail[0]),
		.chany_top_out(sb_1__1__57_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__57_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__57_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__57_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__57_ccff_tail[0]));

	sb_1__1_ sb_6__4_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__64_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_64_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_64_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_64_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_64_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_64_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_64_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_64_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_64_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__1__69_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_76_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_76_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_76_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_76_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_76_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_76_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_76_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_76_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_1__1__63_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_63_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_63_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_63_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_63_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_63_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_63_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_63_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_63_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__58_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_64_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_64_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_64_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_64_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_64_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_64_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_64_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_64_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(cbx_1__1__69_ccff_tail[0]),
		.chany_top_out(sb_1__1__58_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__58_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__58_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__58_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__58_ccff_tail[0]));

	sb_1__1_ sb_6__5_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__65_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_65_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_65_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_65_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_65_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_65_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_65_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_65_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_65_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__1__70_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_77_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_77_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_77_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_77_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_77_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_77_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_77_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_77_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_1__1__64_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_64_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_64_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_64_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_64_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_64_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_64_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_64_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_64_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__59_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_65_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_65_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_65_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_65_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_65_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_65_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_65_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_65_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(cbx_1__1__70_ccff_tail[0]),
		.chany_top_out(sb_1__1__59_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__59_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__59_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__59_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__59_ccff_tail[0]));

	sb_1__1_ sb_6__6_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__66_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_66_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_66_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_66_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_66_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_66_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_66_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_66_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_66_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__1__71_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_78_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_78_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_78_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_78_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_78_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_78_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_78_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_78_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_1__1__65_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_65_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_65_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_65_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_65_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_65_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_65_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_65_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_65_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__60_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_66_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_66_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_66_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_66_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_66_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_66_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_66_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_66_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(cbx_1__1__71_ccff_tail[0]),
		.chany_top_out(sb_1__1__60_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__60_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__60_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__60_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__60_ccff_tail[0]));

	sb_1__1_ sb_6__7_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__67_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_67_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_67_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_67_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_67_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_67_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_67_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_67_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_67_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__1__72_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_79_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_79_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_79_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_79_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_79_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_79_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_79_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_79_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_1__1__66_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_66_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_66_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_66_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_66_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_66_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_66_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_66_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_66_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__61_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_67_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_67_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_67_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_67_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_67_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_67_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_67_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_67_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(cbx_1__1__72_ccff_tail[0]),
		.chany_top_out(sb_1__1__61_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__61_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__61_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__61_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__61_ccff_tail[0]));

	sb_1__1_ sb_6__8_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__68_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_68_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_68_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_68_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_68_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_68_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_68_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_68_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_68_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__1__73_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_80_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_80_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_80_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_80_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_80_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_80_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_80_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_80_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_1__1__67_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_67_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_67_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_67_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_67_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_67_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_67_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_67_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_67_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__62_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_68_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_68_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_68_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_68_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_68_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_68_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_68_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_68_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(cbx_1__1__73_ccff_tail[0]),
		.chany_top_out(sb_1__1__62_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__62_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__62_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__62_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__62_ccff_tail[0]));

	sb_1__1_ sb_6__9_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__69_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_69_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_69_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_69_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_69_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_69_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_69_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_69_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_69_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__1__74_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_81_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_81_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_81_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_81_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_81_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_81_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_81_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_81_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_1__1__68_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_68_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_68_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_68_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_68_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_68_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_68_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_68_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_68_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__63_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_69_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_69_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_69_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_69_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_69_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_69_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_69_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_69_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(cbx_1__1__74_ccff_tail[0]),
		.chany_top_out(sb_1__1__63_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__63_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__63_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__63_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__63_ccff_tail[0]));

	sb_1__1_ sb_6__10_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__70_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_70_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_70_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_70_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_70_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_70_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_70_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_70_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_70_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__1__75_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_82_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_82_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_82_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_82_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_82_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_82_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_82_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_82_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_1__1__69_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_69_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_69_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_69_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_69_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_69_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_69_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_69_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_69_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__64_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_70_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_70_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_70_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_70_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_70_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_70_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_70_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_70_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(cbx_1__1__75_ccff_tail[0]),
		.chany_top_out(sb_1__1__64_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__64_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__64_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__64_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__64_ccff_tail[0]));

	sb_1__1_ sb_6__11_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__71_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_71_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_71_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_71_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_71_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_71_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_71_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_71_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_71_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__1__76_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_83_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_83_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_83_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_83_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_83_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_83_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_83_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_83_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_1__1__70_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_70_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_70_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_70_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_70_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_70_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_70_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_70_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_70_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__65_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_71_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_71_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_71_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_71_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_71_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_71_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_71_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_71_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(cbx_1__1__76_ccff_tail[0]),
		.chany_top_out(sb_1__1__65_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__65_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__65_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__65_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__65_ccff_tail[0]));

	sb_1__1_ sb_7__1_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__73_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_73_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_73_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_73_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_73_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_73_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_73_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_73_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_73_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__1__77_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_85_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_85_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_85_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_85_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_85_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_85_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_85_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_85_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_1__1__72_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_72_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_72_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_72_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_72_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_72_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_72_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_72_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_72_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__66_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_73_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_73_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_73_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_73_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_73_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_73_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_73_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_73_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(cbx_1__1__77_ccff_tail[0]),
		.chany_top_out(sb_1__1__66_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__66_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__66_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__66_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__66_ccff_tail[0]));

	sb_1__1_ sb_7__2_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__74_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_74_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_74_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_74_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_74_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_74_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_74_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_74_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_74_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__1__78_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_86_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_86_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_86_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_86_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_86_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_86_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_86_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_86_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_1__1__73_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_73_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_73_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_73_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_73_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_73_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_73_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_73_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_73_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__67_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_74_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_74_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_74_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_74_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_74_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_74_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_74_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_74_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(cbx_1__1__78_ccff_tail[0]),
		.chany_top_out(sb_1__1__67_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__67_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__67_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__67_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__67_ccff_tail[0]));

	sb_1__1_ sb_7__3_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__75_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_75_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_75_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_75_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_75_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_75_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_75_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_75_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_75_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__1__79_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_87_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_87_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_87_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_87_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_87_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_87_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_87_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_87_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_1__1__74_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_74_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_74_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_74_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_74_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_74_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_74_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_74_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_74_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__68_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_75_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_75_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_75_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_75_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_75_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_75_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_75_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_75_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(cbx_1__1__79_ccff_tail[0]),
		.chany_top_out(sb_1__1__68_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__68_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__68_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__68_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__68_ccff_tail[0]));

	sb_1__1_ sb_7__4_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__76_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_76_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_76_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_76_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_76_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_76_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_76_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_76_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_76_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__1__80_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_88_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_88_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_88_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_88_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_88_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_88_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_88_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_88_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_1__1__75_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_75_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_75_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_75_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_75_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_75_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_75_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_75_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_75_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__69_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_76_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_76_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_76_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_76_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_76_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_76_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_76_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_76_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(cbx_1__1__80_ccff_tail[0]),
		.chany_top_out(sb_1__1__69_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__69_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__69_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__69_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__69_ccff_tail[0]));

	sb_1__1_ sb_7__5_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__77_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_77_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_77_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_77_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_77_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_77_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_77_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_77_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_77_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__1__81_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_89_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_89_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_89_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_89_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_89_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_89_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_89_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_89_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_1__1__76_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_76_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_76_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_76_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_76_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_76_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_76_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_76_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_76_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__70_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_77_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_77_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_77_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_77_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_77_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_77_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_77_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_77_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(cbx_1__1__81_ccff_tail[0]),
		.chany_top_out(sb_1__1__70_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__70_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__70_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__70_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__70_ccff_tail[0]));

	sb_1__1_ sb_7__6_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__78_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_78_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_78_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_78_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_78_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_78_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_78_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_78_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_78_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__1__82_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_90_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_90_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_90_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_90_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_90_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_90_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_90_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_90_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_1__1__77_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_77_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_77_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_77_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_77_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_77_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_77_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_77_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_77_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__71_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_78_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_78_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_78_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_78_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_78_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_78_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_78_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_78_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(cbx_1__1__82_ccff_tail[0]),
		.chany_top_out(sb_1__1__71_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__71_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__71_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__71_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__71_ccff_tail[0]));

	sb_1__1_ sb_7__7_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__79_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_79_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_79_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_79_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_79_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_79_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_79_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_79_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_79_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__1__83_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_91_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_91_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_91_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_91_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_91_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_91_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_91_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_91_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_1__1__78_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_78_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_78_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_78_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_78_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_78_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_78_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_78_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_78_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__72_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_79_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_79_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_79_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_79_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_79_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_79_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_79_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_79_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(cbx_1__1__83_ccff_tail[0]),
		.chany_top_out(sb_1__1__72_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__72_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__72_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__72_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__72_ccff_tail[0]));

	sb_1__1_ sb_7__8_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__80_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_80_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_80_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_80_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_80_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_80_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_80_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_80_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_80_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__1__84_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_92_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_92_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_92_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_92_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_92_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_92_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_92_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_92_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_1__1__79_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_79_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_79_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_79_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_79_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_79_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_79_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_79_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_79_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__73_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_80_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_80_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_80_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_80_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_80_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_80_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_80_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_80_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(cbx_1__1__84_ccff_tail[0]),
		.chany_top_out(sb_1__1__73_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__73_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__73_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__73_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__73_ccff_tail[0]));

	sb_1__1_ sb_7__9_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__81_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_81_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_81_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_81_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_81_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_81_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_81_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_81_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_81_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__1__85_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_93_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_93_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_93_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_93_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_93_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_93_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_93_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_93_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_1__1__80_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_80_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_80_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_80_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_80_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_80_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_80_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_80_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_80_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__74_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_81_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_81_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_81_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_81_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_81_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_81_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_81_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_81_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(cbx_1__1__85_ccff_tail[0]),
		.chany_top_out(sb_1__1__74_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__74_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__74_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__74_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__74_ccff_tail[0]));

	sb_1__1_ sb_7__10_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__82_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_82_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_82_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_82_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_82_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_82_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_82_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_82_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_82_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__1__86_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_94_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_94_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_94_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_94_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_94_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_94_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_94_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_94_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_1__1__81_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_81_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_81_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_81_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_81_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_81_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_81_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_81_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_81_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__75_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_82_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_82_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_82_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_82_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_82_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_82_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_82_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_82_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(cbx_1__1__86_ccff_tail[0]),
		.chany_top_out(sb_1__1__75_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__75_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__75_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__75_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__75_ccff_tail[0]));

	sb_1__1_ sb_7__11_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__83_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_83_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_83_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_83_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_83_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_83_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_83_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_83_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_83_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__1__87_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_95_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_95_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_95_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_95_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_95_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_95_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_95_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_95_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_1__1__82_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_82_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_82_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_82_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_82_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_82_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_82_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_82_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_82_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__76_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_83_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_83_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_83_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_83_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_83_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_83_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_83_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_83_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(cbx_1__1__87_ccff_tail[0]),
		.chany_top_out(sb_1__1__76_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__76_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__76_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__76_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__76_ccff_tail[0]));

	sb_1__1_ sb_8__1_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__85_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_85_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_85_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_85_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_85_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_85_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_85_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_85_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_85_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__1__88_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_97_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_97_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_97_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_97_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_97_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_97_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_97_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_97_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_1__1__84_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_84_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_84_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_84_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_84_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_84_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_84_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_84_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_84_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__77_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_85_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_85_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_85_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_85_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_85_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_85_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_85_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_85_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(cbx_1__1__88_ccff_tail[0]),
		.chany_top_out(sb_1__1__77_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__77_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__77_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__77_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__77_ccff_tail[0]));

	sb_1__1_ sb_8__2_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__86_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_86_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_86_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_86_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_86_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_86_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_86_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_86_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_86_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__1__89_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_98_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_98_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_98_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_98_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_98_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_98_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_98_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_98_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_1__1__85_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_85_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_85_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_85_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_85_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_85_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_85_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_85_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_85_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__78_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_86_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_86_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_86_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_86_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_86_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_86_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_86_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_86_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(cbx_1__1__89_ccff_tail[0]),
		.chany_top_out(sb_1__1__78_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__78_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__78_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__78_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__78_ccff_tail[0]));

	sb_1__1_ sb_8__3_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__87_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_87_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_87_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_87_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_87_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_87_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_87_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_87_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_87_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__1__90_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_99_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_99_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_99_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_99_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_99_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_99_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_99_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_99_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_1__1__86_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_86_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_86_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_86_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_86_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_86_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_86_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_86_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_86_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__79_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_87_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_87_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_87_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_87_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_87_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_87_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_87_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_87_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(cbx_1__1__90_ccff_tail[0]),
		.chany_top_out(sb_1__1__79_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__79_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__79_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__79_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__79_ccff_tail[0]));

	sb_1__1_ sb_8__4_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__88_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_88_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_88_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_88_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_88_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_88_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_88_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_88_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_88_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__1__91_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_100_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_100_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_100_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_100_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_100_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_100_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_100_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_100_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_1__1__87_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_87_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_87_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_87_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_87_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_87_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_87_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_87_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_87_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__80_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_88_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_88_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_88_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_88_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_88_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_88_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_88_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_88_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(cbx_1__1__91_ccff_tail[0]),
		.chany_top_out(sb_1__1__80_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__80_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__80_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__80_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__80_ccff_tail[0]));

	sb_1__1_ sb_8__5_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__89_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_89_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_89_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_89_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_89_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_89_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_89_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_89_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_89_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__1__92_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_101_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_101_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_101_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_101_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_101_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_101_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_101_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_101_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_1__1__88_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_88_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_88_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_88_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_88_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_88_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_88_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_88_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_88_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__81_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_89_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_89_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_89_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_89_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_89_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_89_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_89_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_89_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(cbx_1__1__92_ccff_tail[0]),
		.chany_top_out(sb_1__1__81_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__81_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__81_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__81_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__81_ccff_tail[0]));

	sb_1__1_ sb_8__6_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__90_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_90_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_90_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_90_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_90_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_90_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_90_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_90_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_90_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__1__93_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_102_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_102_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_102_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_102_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_102_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_102_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_102_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_102_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_1__1__89_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_89_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_89_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_89_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_89_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_89_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_89_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_89_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_89_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__82_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_90_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_90_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_90_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_90_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_90_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_90_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_90_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_90_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(cbx_1__1__93_ccff_tail[0]),
		.chany_top_out(sb_1__1__82_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__82_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__82_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__82_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__82_ccff_tail[0]));

	sb_1__1_ sb_8__7_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__91_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_91_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_91_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_91_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_91_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_91_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_91_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_91_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_91_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__1__94_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_103_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_103_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_103_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_103_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_103_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_103_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_103_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_103_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_1__1__90_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_90_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_90_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_90_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_90_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_90_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_90_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_90_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_90_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__83_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_91_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_91_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_91_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_91_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_91_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_91_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_91_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_91_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(cbx_1__1__94_ccff_tail[0]),
		.chany_top_out(sb_1__1__83_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__83_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__83_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__83_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__83_ccff_tail[0]));

	sb_1__1_ sb_8__8_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__92_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_92_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_92_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_92_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_92_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_92_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_92_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_92_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_92_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__1__95_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_104_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_104_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_104_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_104_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_104_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_104_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_104_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_104_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_1__1__91_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_91_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_91_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_91_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_91_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_91_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_91_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_91_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_91_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__84_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_92_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_92_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_92_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_92_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_92_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_92_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_92_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_92_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(cbx_1__1__95_ccff_tail[0]),
		.chany_top_out(sb_1__1__84_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__84_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__84_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__84_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__84_ccff_tail[0]));

	sb_1__1_ sb_8__9_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__93_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_93_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_93_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_93_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_93_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_93_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_93_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_93_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_93_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__1__96_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_105_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_105_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_105_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_105_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_105_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_105_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_105_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_105_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_1__1__92_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_92_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_92_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_92_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_92_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_92_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_92_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_92_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_92_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__85_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_93_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_93_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_93_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_93_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_93_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_93_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_93_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_93_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(cbx_1__1__96_ccff_tail[0]),
		.chany_top_out(sb_1__1__85_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__85_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__85_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__85_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__85_ccff_tail[0]));

	sb_1__1_ sb_8__10_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__94_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_94_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_94_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_94_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_94_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_94_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_94_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_94_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_94_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__1__97_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_106_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_106_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_106_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_106_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_106_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_106_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_106_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_106_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_1__1__93_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_93_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_93_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_93_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_93_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_93_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_93_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_93_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_93_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__86_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_94_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_94_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_94_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_94_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_94_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_94_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_94_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_94_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(cbx_1__1__97_ccff_tail[0]),
		.chany_top_out(sb_1__1__86_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__86_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__86_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__86_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__86_ccff_tail[0]));

	sb_1__1_ sb_8__11_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__95_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_95_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_95_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_95_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_95_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_95_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_95_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_95_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_95_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__1__98_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_107_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_107_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_107_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_107_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_107_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_107_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_107_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_107_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_1__1__94_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_94_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_94_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_94_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_94_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_94_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_94_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_94_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_94_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__87_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_95_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_95_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_95_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_95_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_95_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_95_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_95_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_95_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(cbx_1__1__98_ccff_tail[0]),
		.chany_top_out(sb_1__1__87_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__87_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__87_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__87_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__87_ccff_tail[0]));

	sb_1__1_ sb_9__1_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__97_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_97_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_97_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_97_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_97_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_97_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_97_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_97_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_97_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__1__99_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_109_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_109_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_109_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_109_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_109_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_109_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_109_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_109_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_1__1__96_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_96_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_96_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_96_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_96_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_96_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_96_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_96_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_96_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__88_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_97_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_97_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_97_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_97_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_97_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_97_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_97_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_97_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(cbx_1__1__99_ccff_tail[0]),
		.chany_top_out(sb_1__1__88_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__88_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__88_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__88_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__88_ccff_tail[0]));

	sb_1__1_ sb_9__2_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__98_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_98_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_98_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_98_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_98_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_98_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_98_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_98_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_98_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__1__100_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_110_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_110_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_110_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_110_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_110_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_110_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_110_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_110_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_1__1__97_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_97_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_97_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_97_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_97_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_97_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_97_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_97_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_97_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__89_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_98_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_98_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_98_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_98_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_98_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_98_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_98_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_98_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(cbx_1__1__100_ccff_tail[0]),
		.chany_top_out(sb_1__1__89_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__89_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__89_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__89_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__89_ccff_tail[0]));

	sb_1__1_ sb_9__3_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__99_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_99_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_99_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_99_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_99_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_99_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_99_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_99_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_99_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__1__101_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_111_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_111_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_111_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_111_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_111_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_111_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_111_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_111_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_1__1__98_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_98_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_98_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_98_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_98_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_98_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_98_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_98_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_98_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__90_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_99_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_99_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_99_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_99_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_99_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_99_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_99_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_99_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(cbx_1__1__101_ccff_tail[0]),
		.chany_top_out(sb_1__1__90_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__90_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__90_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__90_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__90_ccff_tail[0]));

	sb_1__1_ sb_9__4_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__100_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_100_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_100_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_100_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_100_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_100_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_100_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_100_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_100_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__1__102_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_112_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_112_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_112_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_112_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_112_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_112_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_112_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_112_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_1__1__99_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_99_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_99_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_99_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_99_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_99_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_99_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_99_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_99_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__91_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_100_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_100_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_100_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_100_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_100_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_100_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_100_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_100_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(cbx_1__1__102_ccff_tail[0]),
		.chany_top_out(sb_1__1__91_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__91_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__91_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__91_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__91_ccff_tail[0]));

	sb_1__1_ sb_9__5_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__101_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_101_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_101_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_101_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_101_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_101_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_101_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_101_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_101_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__1__103_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_113_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_113_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_113_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_113_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_113_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_113_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_113_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_113_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_1__1__100_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_100_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_100_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_100_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_100_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_100_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_100_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_100_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_100_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__92_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_101_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_101_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_101_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_101_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_101_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_101_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_101_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_101_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(cbx_1__1__103_ccff_tail[0]),
		.chany_top_out(sb_1__1__92_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__92_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__92_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__92_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__92_ccff_tail[0]));

	sb_1__1_ sb_9__6_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__102_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_102_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_102_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_102_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_102_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_102_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_102_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_102_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_102_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__1__104_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_114_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_114_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_114_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_114_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_114_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_114_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_114_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_114_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_1__1__101_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_101_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_101_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_101_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_101_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_101_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_101_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_101_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_101_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__93_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_102_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_102_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_102_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_102_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_102_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_102_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_102_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_102_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(cbx_1__1__104_ccff_tail[0]),
		.chany_top_out(sb_1__1__93_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__93_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__93_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__93_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__93_ccff_tail[0]));

	sb_1__1_ sb_9__7_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__103_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_103_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_103_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_103_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_103_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_103_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_103_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_103_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_103_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__1__105_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_115_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_115_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_115_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_115_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_115_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_115_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_115_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_115_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_1__1__102_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_102_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_102_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_102_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_102_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_102_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_102_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_102_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_102_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__94_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_103_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_103_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_103_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_103_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_103_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_103_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_103_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_103_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(cbx_1__1__105_ccff_tail[0]),
		.chany_top_out(sb_1__1__94_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__94_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__94_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__94_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__94_ccff_tail[0]));

	sb_1__1_ sb_9__8_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__104_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_104_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_104_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_104_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_104_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_104_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_104_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_104_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_104_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__1__106_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_116_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_116_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_116_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_116_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_116_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_116_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_116_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_116_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_1__1__103_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_103_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_103_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_103_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_103_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_103_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_103_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_103_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_103_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__95_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_104_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_104_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_104_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_104_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_104_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_104_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_104_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_104_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(cbx_1__1__106_ccff_tail[0]),
		.chany_top_out(sb_1__1__95_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__95_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__95_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__95_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__95_ccff_tail[0]));

	sb_1__1_ sb_9__9_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__105_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_105_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_105_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_105_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_105_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_105_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_105_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_105_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_105_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__1__107_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_117_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_117_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_117_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_117_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_117_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_117_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_117_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_117_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_1__1__104_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_104_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_104_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_104_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_104_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_104_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_104_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_104_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_104_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__96_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_105_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_105_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_105_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_105_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_105_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_105_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_105_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_105_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(cbx_1__1__107_ccff_tail[0]),
		.chany_top_out(sb_1__1__96_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__96_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__96_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__96_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__96_ccff_tail[0]));

	sb_1__1_ sb_9__10_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__106_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_106_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_106_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_106_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_106_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_106_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_106_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_106_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_106_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__1__108_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_118_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_118_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_118_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_118_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_118_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_118_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_118_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_118_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_1__1__105_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_105_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_105_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_105_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_105_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_105_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_105_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_105_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_105_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__97_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_106_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_106_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_106_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_106_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_106_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_106_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_106_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_106_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(cbx_1__1__108_ccff_tail[0]),
		.chany_top_out(sb_1__1__97_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__97_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__97_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__97_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__97_ccff_tail[0]));

	sb_1__1_ sb_9__11_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__107_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_107_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_107_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_107_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_107_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_107_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_107_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_107_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_107_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__1__109_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_119_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_119_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_119_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_119_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_119_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_119_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_119_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_119_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_1__1__106_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_106_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_106_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_106_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_106_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_106_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_106_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_106_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_106_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__98_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_107_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_107_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_107_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_107_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_107_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_107_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_107_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_107_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(cbx_1__1__109_ccff_tail[0]),
		.chany_top_out(sb_1__1__98_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__98_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__98_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__98_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__98_ccff_tail[0]));

	sb_1__1_ sb_10__1_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__109_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_109_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_109_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_109_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_109_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_109_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_109_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_109_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_109_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__1__110_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_121_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_121_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_121_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_121_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_121_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_121_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_121_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_121_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_1__1__108_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_108_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_108_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_108_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_108_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_108_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_108_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_108_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_108_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__99_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_109_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_109_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_109_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_109_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_109_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_109_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_109_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_109_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(cbx_1__1__110_ccff_tail[0]),
		.chany_top_out(sb_1__1__99_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__99_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__99_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__99_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__99_ccff_tail[0]));

	sb_1__1_ sb_10__2_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__110_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_110_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_110_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_110_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_110_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_110_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_110_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_110_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_110_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__1__111_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_122_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_122_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_122_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_122_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_122_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_122_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_122_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_122_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_1__1__109_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_109_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_109_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_109_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_109_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_109_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_109_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_109_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_109_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__100_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_110_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_110_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_110_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_110_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_110_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_110_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_110_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_110_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(cbx_1__1__111_ccff_tail[0]),
		.chany_top_out(sb_1__1__100_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__100_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__100_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__100_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__100_ccff_tail[0]));

	sb_1__1_ sb_10__3_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__111_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_111_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_111_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_111_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_111_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_111_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_111_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_111_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_111_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__1__112_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_123_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_123_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_123_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_123_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_123_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_123_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_123_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_123_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_1__1__110_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_110_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_110_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_110_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_110_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_110_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_110_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_110_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_110_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__101_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_111_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_111_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_111_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_111_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_111_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_111_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_111_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_111_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(cbx_1__1__112_ccff_tail[0]),
		.chany_top_out(sb_1__1__101_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__101_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__101_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__101_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__101_ccff_tail[0]));

	sb_1__1_ sb_10__4_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__112_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_112_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_112_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_112_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_112_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_112_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_112_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_112_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_112_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__1__113_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_124_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_124_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_124_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_124_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_124_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_124_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_124_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_124_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_1__1__111_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_111_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_111_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_111_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_111_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_111_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_111_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_111_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_111_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__102_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_112_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_112_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_112_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_112_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_112_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_112_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_112_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_112_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(cbx_1__1__113_ccff_tail[0]),
		.chany_top_out(sb_1__1__102_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__102_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__102_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__102_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__102_ccff_tail[0]));

	sb_1__1_ sb_10__5_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__113_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_113_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_113_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_113_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_113_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_113_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_113_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_113_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_113_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__1__114_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_125_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_125_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_125_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_125_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_125_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_125_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_125_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_125_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_1__1__112_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_112_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_112_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_112_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_112_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_112_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_112_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_112_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_112_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__103_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_113_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_113_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_113_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_113_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_113_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_113_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_113_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_113_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(cbx_1__1__114_ccff_tail[0]),
		.chany_top_out(sb_1__1__103_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__103_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__103_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__103_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__103_ccff_tail[0]));

	sb_1__1_ sb_10__6_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__114_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_114_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_114_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_114_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_114_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_114_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_114_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_114_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_114_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__1__115_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_126_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_126_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_126_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_126_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_126_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_126_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_126_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_126_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_1__1__113_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_113_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_113_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_113_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_113_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_113_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_113_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_113_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_113_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__104_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_114_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_114_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_114_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_114_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_114_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_114_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_114_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_114_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(cbx_1__1__115_ccff_tail[0]),
		.chany_top_out(sb_1__1__104_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__104_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__104_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__104_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__104_ccff_tail[0]));

	sb_1__1_ sb_10__7_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__115_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_115_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_115_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_115_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_115_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_115_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_115_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_115_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_115_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__1__116_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_127_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_127_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_127_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_127_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_127_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_127_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_127_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_127_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_1__1__114_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_114_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_114_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_114_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_114_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_114_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_114_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_114_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_114_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__105_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_115_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_115_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_115_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_115_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_115_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_115_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_115_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_115_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(cbx_1__1__116_ccff_tail[0]),
		.chany_top_out(sb_1__1__105_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__105_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__105_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__105_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__105_ccff_tail[0]));

	sb_1__1_ sb_10__8_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__116_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_116_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_116_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_116_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_116_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_116_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_116_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_116_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_116_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__1__117_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_128_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_128_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_128_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_128_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_128_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_128_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_128_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_128_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_1__1__115_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_115_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_115_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_115_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_115_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_115_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_115_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_115_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_115_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__106_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_116_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_116_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_116_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_116_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_116_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_116_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_116_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_116_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(cbx_1__1__117_ccff_tail[0]),
		.chany_top_out(sb_1__1__106_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__106_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__106_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__106_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__106_ccff_tail[0]));

	sb_1__1_ sb_10__9_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__117_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_117_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_117_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_117_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_117_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_117_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_117_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_117_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_117_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__1__118_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_129_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_129_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_129_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_129_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_129_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_129_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_129_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_129_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_1__1__116_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_116_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_116_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_116_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_116_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_116_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_116_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_116_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_116_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__107_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_117_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_117_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_117_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_117_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_117_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_117_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_117_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_117_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(cbx_1__1__118_ccff_tail[0]),
		.chany_top_out(sb_1__1__107_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__107_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__107_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__107_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__107_ccff_tail[0]));

	sb_1__1_ sb_10__10_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__118_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_118_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_118_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_118_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_118_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_118_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_118_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_118_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_118_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__1__119_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_130_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_130_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_130_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_130_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_130_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_130_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_130_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_130_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_1__1__117_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_117_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_117_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_117_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_117_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_117_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_117_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_117_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_117_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__108_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_118_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_118_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_118_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_118_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_118_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_118_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_118_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_118_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(cbx_1__1__119_ccff_tail[0]),
		.chany_top_out(sb_1__1__108_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__108_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__108_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__108_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__108_ccff_tail[0]));

	sb_1__1_ sb_10__11_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__119_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_119_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_119_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_119_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_119_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_119_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_119_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_119_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_119_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__1__120_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_131_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_131_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_131_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_131_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_131_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_131_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_131_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_131_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_1__1__118_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_118_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_118_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_118_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_118_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_118_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_118_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_118_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_118_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__109_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_119_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_119_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_119_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_119_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_119_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_119_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_119_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_119_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(cbx_1__1__120_ccff_tail[0]),
		.chany_top_out(sb_1__1__109_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__109_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__109_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__109_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__109_ccff_tail[0]));

	sb_1__1_ sb_11__1_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__121_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_121_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_121_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_121_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_121_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_121_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_121_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_121_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_121_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__1__121_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_133_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_133_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_133_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_133_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_133_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_133_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_133_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_133_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_1__1__120_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_120_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_120_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_120_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_120_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_120_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_120_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_120_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_120_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__110_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_121_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_121_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_121_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_121_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_121_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_121_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_121_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_121_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(cbx_1__1__121_ccff_tail[0]),
		.chany_top_out(sb_1__1__110_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__110_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__110_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__110_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__110_ccff_tail[0]));

	sb_1__1_ sb_11__2_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__122_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_122_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_122_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_122_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_122_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_122_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_122_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_122_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_122_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__1__122_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_134_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_134_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_134_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_134_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_134_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_134_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_134_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_134_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_1__1__121_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_121_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_121_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_121_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_121_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_121_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_121_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_121_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_121_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__111_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_122_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_122_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_122_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_122_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_122_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_122_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_122_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_122_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(cbx_1__1__122_ccff_tail[0]),
		.chany_top_out(sb_1__1__111_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__111_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__111_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__111_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__111_ccff_tail[0]));

	sb_1__1_ sb_11__3_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__123_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_123_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_123_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_123_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_123_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_123_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_123_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_123_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_123_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__1__123_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_135_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_135_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_135_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_135_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_135_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_135_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_135_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_135_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_1__1__122_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_122_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_122_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_122_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_122_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_122_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_122_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_122_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_122_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__112_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_123_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_123_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_123_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_123_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_123_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_123_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_123_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_123_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(cbx_1__1__123_ccff_tail[0]),
		.chany_top_out(sb_1__1__112_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__112_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__112_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__112_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__112_ccff_tail[0]));

	sb_1__1_ sb_11__4_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__124_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_124_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_124_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_124_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_124_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_124_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_124_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_124_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_124_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__1__124_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_136_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_136_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_136_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_136_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_136_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_136_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_136_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_136_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_1__1__123_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_123_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_123_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_123_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_123_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_123_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_123_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_123_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_123_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__113_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_124_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_124_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_124_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_124_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_124_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_124_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_124_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_124_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(cbx_1__1__124_ccff_tail[0]),
		.chany_top_out(sb_1__1__113_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__113_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__113_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__113_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__113_ccff_tail[0]));

	sb_1__1_ sb_11__5_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__125_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_125_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_125_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_125_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_125_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_125_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_125_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_125_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_125_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__1__125_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_137_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_137_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_137_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_137_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_137_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_137_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_137_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_137_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_1__1__124_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_124_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_124_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_124_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_124_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_124_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_124_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_124_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_124_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__114_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_125_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_125_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_125_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_125_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_125_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_125_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_125_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_125_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(cbx_1__1__125_ccff_tail[0]),
		.chany_top_out(sb_1__1__114_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__114_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__114_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__114_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__114_ccff_tail[0]));

	sb_1__1_ sb_11__6_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__126_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_126_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_126_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_126_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_126_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_126_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_126_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_126_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_126_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__1__126_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_138_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_138_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_138_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_138_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_138_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_138_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_138_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_138_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_1__1__125_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_125_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_125_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_125_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_125_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_125_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_125_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_125_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_125_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__115_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_126_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_126_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_126_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_126_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_126_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_126_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_126_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_126_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(cbx_1__1__126_ccff_tail[0]),
		.chany_top_out(sb_1__1__115_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__115_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__115_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__115_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__115_ccff_tail[0]));

	sb_1__1_ sb_11__7_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__127_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_127_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_127_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_127_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_127_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_127_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_127_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_127_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_127_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__1__127_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_139_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_139_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_139_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_139_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_139_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_139_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_139_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_139_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_1__1__126_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_126_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_126_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_126_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_126_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_126_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_126_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_126_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_126_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__116_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_127_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_127_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_127_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_127_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_127_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_127_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_127_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_127_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(cbx_1__1__127_ccff_tail[0]),
		.chany_top_out(sb_1__1__116_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__116_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__116_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__116_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__116_ccff_tail[0]));

	sb_1__1_ sb_11__8_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__128_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_128_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_128_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_128_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_128_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_128_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_128_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_128_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_128_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__1__128_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_140_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_140_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_140_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_140_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_140_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_140_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_140_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_140_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_1__1__127_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_127_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_127_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_127_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_127_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_127_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_127_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_127_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_127_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__117_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_128_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_128_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_128_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_128_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_128_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_128_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_128_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_128_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(cbx_1__1__128_ccff_tail[0]),
		.chany_top_out(sb_1__1__117_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__117_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__117_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__117_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__117_ccff_tail[0]));

	sb_1__1_ sb_11__9_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__129_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_129_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_129_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_129_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_129_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_129_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_129_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_129_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_129_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__1__129_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_141_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_141_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_141_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_141_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_141_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_141_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_141_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_141_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_1__1__128_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_128_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_128_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_128_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_128_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_128_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_128_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_128_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_128_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__118_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_129_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_129_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_129_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_129_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_129_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_129_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_129_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_129_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(cbx_1__1__129_ccff_tail[0]),
		.chany_top_out(sb_1__1__118_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__118_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__118_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__118_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__118_ccff_tail[0]));

	sb_1__1_ sb_11__10_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__130_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_130_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_130_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_130_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_130_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_130_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_130_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_130_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_130_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__1__130_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_142_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_142_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_142_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_142_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_142_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_142_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_142_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_142_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_1__1__129_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_129_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_129_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_129_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_129_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_129_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_129_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_129_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_129_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__119_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_130_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_130_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_130_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_130_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_130_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_130_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_130_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_130_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(cbx_1__1__130_ccff_tail[0]),
		.chany_top_out(sb_1__1__119_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__119_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__119_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__119_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__119_ccff_tail[0]));

	sb_1__1_ sb_11__11_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__131_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_131_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_131_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_131_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_131_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_131_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_131_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_131_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_131_right_width_0_height_0__pin_41_lower[0]),
		.chanx_right_in(cbx_1__1__131_chanx_left_out[0:19]),
		.right_top_grid_pin_42_(grid_clb_143_bottom_width_0_height_0__pin_42_upper[0]),
		.right_top_grid_pin_43_(grid_clb_143_bottom_width_0_height_0__pin_43_upper[0]),
		.right_top_grid_pin_44_(grid_clb_143_bottom_width_0_height_0__pin_44_upper[0]),
		.right_top_grid_pin_45_(grid_clb_143_bottom_width_0_height_0__pin_45_upper[0]),
		.right_top_grid_pin_46_(grid_clb_143_bottom_width_0_height_0__pin_46_upper[0]),
		.right_top_grid_pin_47_(grid_clb_143_bottom_width_0_height_0__pin_47_upper[0]),
		.right_top_grid_pin_48_(grid_clb_143_bottom_width_0_height_0__pin_48_upper[0]),
		.right_top_grid_pin_49_(grid_clb_143_bottom_width_0_height_0__pin_49_upper[0]),
		.chany_bottom_in(cby_1__1__130_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_130_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_130_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_130_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_130_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_130_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_130_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_130_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_130_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__120_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_131_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_131_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_131_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_131_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_131_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_131_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_131_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_131_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(cbx_1__1__131_ccff_tail[0]),
		.chany_top_out(sb_1__1__120_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__120_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__120_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__120_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__120_ccff_tail[0]));

	sb_1__2_ sb_1__12_ (
		.prog_clk(prog_clk[0]),
		.chanx_right_in(cbx_1__12__1_chanx_left_out[0:19]),
		.right_top_grid_pin_1_(grid_io_top_1_bottom_width_0_height_0__pin_1_upper[0]),
		.chany_bottom_in(cby_1__1__11_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_11_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_11_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_11_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_11_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_11_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_11_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_11_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_11_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__12__0_chanx_right_out[0:19]),
		.left_top_grid_pin_1_(grid_io_top_0_bottom_width_0_height_0__pin_1_lower[0]),
		.ccff_head(grid_io_top_1_ccff_tail[0]),
		.chanx_right_out(sb_1__12__0_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__12__0_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__12__0_chanx_left_out[0:19]),
		.ccff_tail(sb_1__12__0_ccff_tail[0]));

	sb_1__2_ sb_2__12_ (
		.prog_clk(prog_clk[0]),
		.chanx_right_in(cbx_1__12__2_chanx_left_out[0:19]),
		.right_top_grid_pin_1_(grid_io_top_2_bottom_width_0_height_0__pin_1_upper[0]),
		.chany_bottom_in(cby_1__1__23_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_23_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_23_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_23_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_23_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_23_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_23_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_23_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_23_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__12__1_chanx_right_out[0:19]),
		.left_top_grid_pin_1_(grid_io_top_1_bottom_width_0_height_0__pin_1_lower[0]),
		.ccff_head(grid_io_top_2_ccff_tail[0]),
		.chanx_right_out(sb_1__12__1_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__12__1_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__12__1_chanx_left_out[0:19]),
		.ccff_tail(sb_1__12__1_ccff_tail[0]));

	sb_1__2_ sb_3__12_ (
		.prog_clk(prog_clk[0]),
		.chanx_right_in(cbx_1__12__3_chanx_left_out[0:19]),
		.right_top_grid_pin_1_(grid_io_top_3_bottom_width_0_height_0__pin_1_upper[0]),
		.chany_bottom_in(cby_1__1__35_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_35_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_35_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_35_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_35_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_35_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_35_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_35_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_35_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__12__2_chanx_right_out[0:19]),
		.left_top_grid_pin_1_(grid_io_top_2_bottom_width_0_height_0__pin_1_lower[0]),
		.ccff_head(grid_io_top_3_ccff_tail[0]),
		.chanx_right_out(sb_1__12__2_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__12__2_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__12__2_chanx_left_out[0:19]),
		.ccff_tail(sb_1__12__2_ccff_tail[0]));

	sb_1__2_ sb_4__12_ (
		.prog_clk(prog_clk[0]),
		.chanx_right_in(cbx_1__12__4_chanx_left_out[0:19]),
		.right_top_grid_pin_1_(grid_io_top_4_bottom_width_0_height_0__pin_1_upper[0]),
		.chany_bottom_in(cby_1__1__47_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_47_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_47_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_47_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_47_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_47_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_47_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_47_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_47_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__12__3_chanx_right_out[0:19]),
		.left_top_grid_pin_1_(grid_io_top_3_bottom_width_0_height_0__pin_1_lower[0]),
		.ccff_head(grid_io_top_4_ccff_tail[0]),
		.chanx_right_out(sb_1__12__3_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__12__3_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__12__3_chanx_left_out[0:19]),
		.ccff_tail(sb_1__12__3_ccff_tail[0]));

	sb_1__2_ sb_5__12_ (
		.prog_clk(prog_clk[0]),
		.chanx_right_in(cbx_1__12__5_chanx_left_out[0:19]),
		.right_top_grid_pin_1_(grid_io_top_5_bottom_width_0_height_0__pin_1_upper[0]),
		.chany_bottom_in(cby_1__1__59_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_59_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_59_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_59_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_59_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_59_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_59_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_59_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_59_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__12__4_chanx_right_out[0:19]),
		.left_top_grid_pin_1_(grid_io_top_4_bottom_width_0_height_0__pin_1_lower[0]),
		.ccff_head(grid_io_top_5_ccff_tail[0]),
		.chanx_right_out(sb_1__12__4_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__12__4_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__12__4_chanx_left_out[0:19]),
		.ccff_tail(sb_1__12__4_ccff_tail[0]));

	sb_1__2_ sb_6__12_ (
		.prog_clk(prog_clk[0]),
		.chanx_right_in(cbx_1__12__6_chanx_left_out[0:19]),
		.right_top_grid_pin_1_(grid_io_top_6_bottom_width_0_height_0__pin_1_upper[0]),
		.chany_bottom_in(cby_1__1__71_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_71_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_71_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_71_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_71_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_71_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_71_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_71_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_71_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__12__5_chanx_right_out[0:19]),
		.left_top_grid_pin_1_(grid_io_top_5_bottom_width_0_height_0__pin_1_lower[0]),
		.ccff_head(grid_io_top_6_ccff_tail[0]),
		.chanx_right_out(sb_1__12__5_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__12__5_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__12__5_chanx_left_out[0:19]),
		.ccff_tail(sb_1__12__5_ccff_tail[0]));

	sb_1__2_ sb_7__12_ (
		.prog_clk(prog_clk[0]),
		.chanx_right_in(cbx_1__12__7_chanx_left_out[0:19]),
		.right_top_grid_pin_1_(grid_io_top_7_bottom_width_0_height_0__pin_1_upper[0]),
		.chany_bottom_in(cby_1__1__83_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_83_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_83_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_83_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_83_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_83_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_83_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_83_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_83_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__12__6_chanx_right_out[0:19]),
		.left_top_grid_pin_1_(grid_io_top_6_bottom_width_0_height_0__pin_1_lower[0]),
		.ccff_head(grid_io_top_7_ccff_tail[0]),
		.chanx_right_out(sb_1__12__6_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__12__6_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__12__6_chanx_left_out[0:19]),
		.ccff_tail(sb_1__12__6_ccff_tail[0]));

	sb_1__2_ sb_8__12_ (
		.prog_clk(prog_clk[0]),
		.chanx_right_in(cbx_1__12__8_chanx_left_out[0:19]),
		.right_top_grid_pin_1_(grid_io_top_8_bottom_width_0_height_0__pin_1_upper[0]),
		.chany_bottom_in(cby_1__1__95_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_95_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_95_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_95_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_95_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_95_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_95_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_95_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_95_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__12__7_chanx_right_out[0:19]),
		.left_top_grid_pin_1_(grid_io_top_7_bottom_width_0_height_0__pin_1_lower[0]),
		.ccff_head(grid_io_top_8_ccff_tail[0]),
		.chanx_right_out(sb_1__12__7_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__12__7_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__12__7_chanx_left_out[0:19]),
		.ccff_tail(sb_1__12__7_ccff_tail[0]));

	sb_1__2_ sb_9__12_ (
		.prog_clk(prog_clk[0]),
		.chanx_right_in(cbx_1__12__9_chanx_left_out[0:19]),
		.right_top_grid_pin_1_(grid_io_top_9_bottom_width_0_height_0__pin_1_upper[0]),
		.chany_bottom_in(cby_1__1__107_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_107_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_107_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_107_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_107_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_107_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_107_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_107_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_107_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__12__8_chanx_right_out[0:19]),
		.left_top_grid_pin_1_(grid_io_top_8_bottom_width_0_height_0__pin_1_lower[0]),
		.ccff_head(grid_io_top_9_ccff_tail[0]),
		.chanx_right_out(sb_1__12__8_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__12__8_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__12__8_chanx_left_out[0:19]),
		.ccff_tail(sb_1__12__8_ccff_tail[0]));

	sb_1__2_ sb_10__12_ (
		.prog_clk(prog_clk[0]),
		.chanx_right_in(cbx_1__12__10_chanx_left_out[0:19]),
		.right_top_grid_pin_1_(grid_io_top_10_bottom_width_0_height_0__pin_1_upper[0]),
		.chany_bottom_in(cby_1__1__119_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_119_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_119_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_119_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_119_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_119_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_119_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_119_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_119_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__12__9_chanx_right_out[0:19]),
		.left_top_grid_pin_1_(grid_io_top_9_bottom_width_0_height_0__pin_1_lower[0]),
		.ccff_head(grid_io_top_10_ccff_tail[0]),
		.chanx_right_out(sb_1__12__9_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__12__9_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__12__9_chanx_left_out[0:19]),
		.ccff_tail(sb_1__12__9_ccff_tail[0]));

	sb_1__2_ sb_11__12_ (
		.prog_clk(prog_clk[0]),
		.chanx_right_in(cbx_1__12__11_chanx_left_out[0:19]),
		.right_top_grid_pin_1_(grid_io_top_11_bottom_width_0_height_0__pin_1_upper[0]),
		.chany_bottom_in(cby_1__1__131_chany_top_out[0:19]),
		.bottom_left_grid_pin_34_(grid_clb_131_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_131_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_131_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_131_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_131_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_131_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_131_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_131_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__12__10_chanx_right_out[0:19]),
		.left_top_grid_pin_1_(grid_io_top_10_bottom_width_0_height_0__pin_1_lower[0]),
		.ccff_head(grid_io_top_11_ccff_tail[0]),
		.chanx_right_out(sb_1__12__10_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__12__10_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__12__10_chanx_left_out[0:19]),
		.ccff_tail(sb_1__12__10_ccff_tail[0]));

    sb_2__0_ sb_12__0_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__132_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_132_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_132_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_132_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_132_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_132_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_132_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_132_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_132_right_width_0_height_0__pin_41_lower[0]),
		.top_right_grid_pin_1_(grid_io_right_0_left_width_0_height_0__pin_1_lower[0]),
		.chanx_left_in(cbx_1__0__11_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_132_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_132_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_132_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_132_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_132_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_132_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_132_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_132_bottom_width_0_height_0__pin_49_lower[0]),
		.left_bottom_grid_pin_1_(grid_io_bottom_11_top_width_0_height_0__pin_1_lower[0]),
		.ccff_head(grid_io_right_0_ccff_tail[0]),
		.chany_top_out(sb_12__0__0_chany_top_out[0:19]),
		.chanx_left_out(sb_12__0__0_chanx_left_out[0:19]),
		.ccff_tail(sb_12__0__0_ccff_tail[0]));

    sb_2__1_ sb_12__1_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__133_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_133_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_133_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_133_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_133_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_133_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_133_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_133_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_133_right_width_0_height_0__pin_41_lower[0]),
		.top_right_grid_pin_1_(grid_io_right_1_left_width_0_height_0__pin_1_lower[0]),
		.chany_bottom_in(cby_1__1__132_chany_top_out[0:19]),
		.bottom_right_grid_pin_1_(grid_io_right_0_left_width_0_height_0__pin_1_upper[0]),
		.bottom_left_grid_pin_34_(grid_clb_132_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_132_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_132_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_132_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_132_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_132_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_132_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_132_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__121_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_133_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_133_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_133_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_133_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_133_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_133_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_133_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_133_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(grid_io_right_1_ccff_tail[0]),
		.chany_top_out(sb_12__1__0_chany_top_out[0:19]),
		.chany_bottom_out(sb_12__1__0_chany_bottom_out[0:19]),
		.chanx_left_out(sb_12__1__0_chanx_left_out[0:19]),
		.ccff_tail(sb_12__1__0_ccff_tail[0]));

    sb_2__1_ sb_12__2_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__134_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_134_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_134_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_134_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_134_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_134_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_134_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_134_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_134_right_width_0_height_0__pin_41_lower[0]),
		.top_right_grid_pin_1_(grid_io_right_2_left_width_0_height_0__pin_1_lower[0]),
		.chany_bottom_in(cby_1__1__133_chany_top_out[0:19]),
		.bottom_right_grid_pin_1_(grid_io_right_1_left_width_0_height_0__pin_1_upper[0]),
		.bottom_left_grid_pin_34_(grid_clb_133_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_133_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_133_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_133_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_133_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_133_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_133_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_133_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__122_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_134_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_134_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_134_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_134_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_134_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_134_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_134_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_134_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(grid_io_right_2_ccff_tail[0]),
		.chany_top_out(sb_12__1__1_chany_top_out[0:19]),
		.chany_bottom_out(sb_12__1__1_chany_bottom_out[0:19]),
		.chanx_left_out(sb_12__1__1_chanx_left_out[0:19]),
		.ccff_tail(sb_12__1__1_ccff_tail[0]));

    sb_2__1_ sb_12__3_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__135_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_135_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_135_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_135_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_135_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_135_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_135_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_135_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_135_right_width_0_height_0__pin_41_lower[0]),
		.top_right_grid_pin_1_(grid_io_right_3_left_width_0_height_0__pin_1_lower[0]),
		.chany_bottom_in(cby_1__1__134_chany_top_out[0:19]),
		.bottom_right_grid_pin_1_(grid_io_right_2_left_width_0_height_0__pin_1_upper[0]),
		.bottom_left_grid_pin_34_(grid_clb_134_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_134_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_134_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_134_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_134_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_134_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_134_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_134_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__123_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_135_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_135_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_135_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_135_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_135_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_135_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_135_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_135_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(grid_io_right_3_ccff_tail[0]),
		.chany_top_out(sb_12__1__2_chany_top_out[0:19]),
		.chany_bottom_out(sb_12__1__2_chany_bottom_out[0:19]),
		.chanx_left_out(sb_12__1__2_chanx_left_out[0:19]),
		.ccff_tail(sb_12__1__2_ccff_tail[0]));

    sb_2__1_ sb_12__4_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__136_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_136_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_136_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_136_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_136_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_136_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_136_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_136_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_136_right_width_0_height_0__pin_41_lower[0]),
		.top_right_grid_pin_1_(grid_io_right_4_left_width_0_height_0__pin_1_lower[0]),
		.chany_bottom_in(cby_1__1__135_chany_top_out[0:19]),
		.bottom_right_grid_pin_1_(grid_io_right_3_left_width_0_height_0__pin_1_upper[0]),
		.bottom_left_grid_pin_34_(grid_clb_135_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_135_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_135_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_135_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_135_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_135_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_135_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_135_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__124_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_136_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_136_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_136_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_136_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_136_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_136_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_136_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_136_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(grid_io_right_4_ccff_tail[0]),
		.chany_top_out(sb_12__1__3_chany_top_out[0:19]),
		.chany_bottom_out(sb_12__1__3_chany_bottom_out[0:19]),
		.chanx_left_out(sb_12__1__3_chanx_left_out[0:19]),
		.ccff_tail(sb_12__1__3_ccff_tail[0]));

    sb_2__1_ sb_12__5_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__137_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_137_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_137_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_137_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_137_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_137_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_137_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_137_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_137_right_width_0_height_0__pin_41_lower[0]),
		.top_right_grid_pin_1_(grid_io_right_5_left_width_0_height_0__pin_1_lower[0]),
		.chany_bottom_in(cby_1__1__136_chany_top_out[0:19]),
		.bottom_right_grid_pin_1_(grid_io_right_4_left_width_0_height_0__pin_1_upper[0]),
		.bottom_left_grid_pin_34_(grid_clb_136_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_136_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_136_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_136_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_136_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_136_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_136_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_136_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__125_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_137_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_137_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_137_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_137_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_137_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_137_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_137_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_137_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(grid_io_right_5_ccff_tail[0]),
		.chany_top_out(sb_12__1__4_chany_top_out[0:19]),
		.chany_bottom_out(sb_12__1__4_chany_bottom_out[0:19]),
		.chanx_left_out(sb_12__1__4_chanx_left_out[0:19]),
		.ccff_tail(sb_12__1__4_ccff_tail[0]));

    sb_2__1_ sb_12__6_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__138_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_138_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_138_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_138_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_138_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_138_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_138_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_138_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_138_right_width_0_height_0__pin_41_lower[0]),
		.top_right_grid_pin_1_(grid_io_right_6_left_width_0_height_0__pin_1_lower[0]),
		.chany_bottom_in(cby_1__1__137_chany_top_out[0:19]),
		.bottom_right_grid_pin_1_(grid_io_right_5_left_width_0_height_0__pin_1_upper[0]),
		.bottom_left_grid_pin_34_(grid_clb_137_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_137_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_137_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_137_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_137_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_137_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_137_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_137_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__126_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_138_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_138_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_138_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_138_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_138_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_138_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_138_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_138_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(grid_io_right_6_ccff_tail[0]),
		.chany_top_out(sb_12__1__5_chany_top_out[0:19]),
		.chany_bottom_out(sb_12__1__5_chany_bottom_out[0:19]),
		.chanx_left_out(sb_12__1__5_chanx_left_out[0:19]),
		.ccff_tail(sb_12__1__5_ccff_tail[0]));

    sb_2__1_ sb_12__7_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__139_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_139_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_139_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_139_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_139_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_139_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_139_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_139_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_139_right_width_0_height_0__pin_41_lower[0]),
		.top_right_grid_pin_1_(grid_io_right_7_left_width_0_height_0__pin_1_lower[0]),
		.chany_bottom_in(cby_1__1__138_chany_top_out[0:19]),
		.bottom_right_grid_pin_1_(grid_io_right_6_left_width_0_height_0__pin_1_upper[0]),
		.bottom_left_grid_pin_34_(grid_clb_138_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_138_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_138_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_138_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_138_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_138_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_138_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_138_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__127_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_139_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_139_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_139_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_139_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_139_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_139_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_139_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_139_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(grid_io_right_7_ccff_tail[0]),
		.chany_top_out(sb_12__1__6_chany_top_out[0:19]),
		.chany_bottom_out(sb_12__1__6_chany_bottom_out[0:19]),
		.chanx_left_out(sb_12__1__6_chanx_left_out[0:19]),
		.ccff_tail(sb_12__1__6_ccff_tail[0]));

    sb_2__1_ sb_12__8_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__140_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_140_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_140_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_140_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_140_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_140_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_140_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_140_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_140_right_width_0_height_0__pin_41_lower[0]),
		.top_right_grid_pin_1_(grid_io_right_8_left_width_0_height_0__pin_1_lower[0]),
		.chany_bottom_in(cby_1__1__139_chany_top_out[0:19]),
		.bottom_right_grid_pin_1_(grid_io_right_7_left_width_0_height_0__pin_1_upper[0]),
		.bottom_left_grid_pin_34_(grid_clb_139_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_139_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_139_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_139_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_139_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_139_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_139_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_139_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__128_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_140_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_140_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_140_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_140_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_140_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_140_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_140_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_140_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(grid_io_right_8_ccff_tail[0]),
		.chany_top_out(sb_12__1__7_chany_top_out[0:19]),
		.chany_bottom_out(sb_12__1__7_chany_bottom_out[0:19]),
		.chanx_left_out(sb_12__1__7_chanx_left_out[0:19]),
		.ccff_tail(sb_12__1__7_ccff_tail[0]));

    sb_2__1_ sb_12__9_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__141_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_141_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_141_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_141_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_141_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_141_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_141_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_141_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_141_right_width_0_height_0__pin_41_lower[0]),
		.top_right_grid_pin_1_(grid_io_right_9_left_width_0_height_0__pin_1_lower[0]),
		.chany_bottom_in(cby_1__1__140_chany_top_out[0:19]),
		.bottom_right_grid_pin_1_(grid_io_right_8_left_width_0_height_0__pin_1_upper[0]),
		.bottom_left_grid_pin_34_(grid_clb_140_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_140_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_140_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_140_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_140_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_140_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_140_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_140_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__129_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_141_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_141_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_141_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_141_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_141_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_141_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_141_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_141_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(grid_io_right_9_ccff_tail[0]),
		.chany_top_out(sb_12__1__8_chany_top_out[0:19]),
		.chany_bottom_out(sb_12__1__8_chany_bottom_out[0:19]),
		.chanx_left_out(sb_12__1__8_chanx_left_out[0:19]),
		.ccff_tail(sb_12__1__8_ccff_tail[0]));

    sb_2__1_ sb_12__10_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__142_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_142_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_142_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_142_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_142_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_142_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_142_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_142_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_142_right_width_0_height_0__pin_41_lower[0]),
		.top_right_grid_pin_1_(grid_io_right_10_left_width_0_height_0__pin_1_lower[0]),
		.chany_bottom_in(cby_1__1__141_chany_top_out[0:19]),
		.bottom_right_grid_pin_1_(grid_io_right_9_left_width_0_height_0__pin_1_upper[0]),
		.bottom_left_grid_pin_34_(grid_clb_141_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_141_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_141_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_141_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_141_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_141_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_141_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_141_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__130_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_142_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_142_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_142_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_142_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_142_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_142_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_142_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_142_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(grid_io_right_10_ccff_tail[0]),
		.chany_top_out(sb_12__1__9_chany_top_out[0:19]),
		.chany_bottom_out(sb_12__1__9_chany_bottom_out[0:19]),
		.chanx_left_out(sb_12__1__9_chanx_left_out[0:19]),
		.ccff_tail(sb_12__1__9_ccff_tail[0]));

    sb_2__1_ sb_12__11_ (
		.prog_clk(prog_clk[0]),
		.chany_top_in(cby_1__1__143_chany_bottom_out[0:19]),
		.top_left_grid_pin_34_(grid_clb_143_right_width_0_height_0__pin_34_lower[0]),
		.top_left_grid_pin_35_(grid_clb_143_right_width_0_height_0__pin_35_lower[0]),
		.top_left_grid_pin_36_(grid_clb_143_right_width_0_height_0__pin_36_lower[0]),
		.top_left_grid_pin_37_(grid_clb_143_right_width_0_height_0__pin_37_lower[0]),
		.top_left_grid_pin_38_(grid_clb_143_right_width_0_height_0__pin_38_lower[0]),
		.top_left_grid_pin_39_(grid_clb_143_right_width_0_height_0__pin_39_lower[0]),
		.top_left_grid_pin_40_(grid_clb_143_right_width_0_height_0__pin_40_lower[0]),
		.top_left_grid_pin_41_(grid_clb_143_right_width_0_height_0__pin_41_lower[0]),
		.top_right_grid_pin_1_(grid_io_right_11_left_width_0_height_0__pin_1_lower[0]),
		.chany_bottom_in(cby_1__1__142_chany_top_out[0:19]),
		.bottom_right_grid_pin_1_(grid_io_right_10_left_width_0_height_0__pin_1_upper[0]),
		.bottom_left_grid_pin_34_(grid_clb_142_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_142_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_142_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_142_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_142_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_142_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_142_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_142_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__1__131_chanx_right_out[0:19]),
		.left_top_grid_pin_42_(grid_clb_143_bottom_width_0_height_0__pin_42_lower[0]),
		.left_top_grid_pin_43_(grid_clb_143_bottom_width_0_height_0__pin_43_lower[0]),
		.left_top_grid_pin_44_(grid_clb_143_bottom_width_0_height_0__pin_44_lower[0]),
		.left_top_grid_pin_45_(grid_clb_143_bottom_width_0_height_0__pin_45_lower[0]),
		.left_top_grid_pin_46_(grid_clb_143_bottom_width_0_height_0__pin_46_lower[0]),
		.left_top_grid_pin_47_(grid_clb_143_bottom_width_0_height_0__pin_47_lower[0]),
		.left_top_grid_pin_48_(grid_clb_143_bottom_width_0_height_0__pin_48_lower[0]),
		.left_top_grid_pin_49_(grid_clb_143_bottom_width_0_height_0__pin_49_lower[0]),
		.ccff_head(grid_io_right_11_ccff_tail[0]),
		.chany_top_out(sb_12__1__10_chany_top_out[0:19]),
		.chany_bottom_out(sb_12__1__10_chany_bottom_out[0:19]),
		.chanx_left_out(sb_12__1__10_chanx_left_out[0:19]),
		.ccff_tail(sb_12__1__10_ccff_tail[0]));

    sb_2__2_ sb_12__12_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(cby_1__1__143_chany_top_out[0:19]),
		.bottom_right_grid_pin_1_(grid_io_right_11_left_width_0_height_0__pin_1_upper[0]),
		.bottom_left_grid_pin_34_(grid_clb_143_right_width_0_height_0__pin_34_upper[0]),
		.bottom_left_grid_pin_35_(grid_clb_143_right_width_0_height_0__pin_35_upper[0]),
		.bottom_left_grid_pin_36_(grid_clb_143_right_width_0_height_0__pin_36_upper[0]),
		.bottom_left_grid_pin_37_(grid_clb_143_right_width_0_height_0__pin_37_upper[0]),
		.bottom_left_grid_pin_38_(grid_clb_143_right_width_0_height_0__pin_38_upper[0]),
		.bottom_left_grid_pin_39_(grid_clb_143_right_width_0_height_0__pin_39_upper[0]),
		.bottom_left_grid_pin_40_(grid_clb_143_right_width_0_height_0__pin_40_upper[0]),
		.bottom_left_grid_pin_41_(grid_clb_143_right_width_0_height_0__pin_41_upper[0]),
		.chanx_left_in(cbx_1__12__11_chanx_right_out[0:19]),
		.left_top_grid_pin_1_(grid_io_top_11_bottom_width_0_height_0__pin_1_lower[0]),
		.ccff_head(ccff_head[0]),
		.chany_bottom_out(sb_12__12__0_chany_bottom_out[0:19]),
		.chanx_left_out(sb_12__12__0_chanx_left_out[0:19]),
		.ccff_tail(sb_12__12__0_ccff_tail[0]));

	cbx_1__0_ cbx_1__0_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_0__0__0_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__0__0_chanx_left_out[0:19]),
		.ccff_head(sb_1__0__0_ccff_tail[0]),
		.chanx_left_out(cbx_1__0__0_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__0__0_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__0__0_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__0__0_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__0__0_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__0__0_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__0__0_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__0__0_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__0__0_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__0__0_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__0__0_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__0__0_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__0__0_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__0__0_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__0__0_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__0__0_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__0__0_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__0__0_top_grid_pin_31_[0]),
		.bottom_grid_pin_0_(cbx_1__0__0_bottom_grid_pin_0_[0]),
		.ccff_tail(cbx_1__0__0_ccff_tail[0]));

	cbx_1__0_ cbx_2__0_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__0__0_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__0__1_chanx_left_out[0:19]),
		.ccff_head(sb_1__0__1_ccff_tail[0]),
		.chanx_left_out(cbx_1__0__1_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__0__1_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__0__1_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__0__1_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__0__1_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__0__1_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__0__1_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__0__1_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__0__1_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__0__1_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__0__1_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__0__1_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__0__1_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__0__1_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__0__1_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__0__1_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__0__1_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__0__1_top_grid_pin_31_[0]),
		.bottom_grid_pin_0_(cbx_1__0__1_bottom_grid_pin_0_[0]),
		.ccff_tail(cbx_1__0__1_ccff_tail[0]));

	cbx_1__0_ cbx_3__0_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__0__1_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__0__2_chanx_left_out[0:19]),
		.ccff_head(sb_1__0__2_ccff_tail[0]),
		.chanx_left_out(cbx_1__0__2_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__0__2_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__0__2_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__0__2_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__0__2_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__0__2_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__0__2_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__0__2_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__0__2_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__0__2_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__0__2_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__0__2_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__0__2_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__0__2_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__0__2_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__0__2_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__0__2_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__0__2_top_grid_pin_31_[0]),
		.bottom_grid_pin_0_(cbx_1__0__2_bottom_grid_pin_0_[0]),
		.ccff_tail(cbx_1__0__2_ccff_tail[0]));

	cbx_1__0_ cbx_4__0_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__0__2_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__0__3_chanx_left_out[0:19]),
		.ccff_head(sb_1__0__3_ccff_tail[0]),
		.chanx_left_out(cbx_1__0__3_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__0__3_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__0__3_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__0__3_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__0__3_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__0__3_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__0__3_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__0__3_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__0__3_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__0__3_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__0__3_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__0__3_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__0__3_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__0__3_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__0__3_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__0__3_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__0__3_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__0__3_top_grid_pin_31_[0]),
		.bottom_grid_pin_0_(cbx_1__0__3_bottom_grid_pin_0_[0]),
		.ccff_tail(cbx_1__0__3_ccff_tail[0]));

	cbx_1__0_ cbx_5__0_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__0__3_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__0__4_chanx_left_out[0:19]),
		.ccff_head(sb_1__0__4_ccff_tail[0]),
		.chanx_left_out(cbx_1__0__4_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__0__4_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__0__4_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__0__4_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__0__4_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__0__4_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__0__4_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__0__4_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__0__4_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__0__4_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__0__4_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__0__4_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__0__4_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__0__4_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__0__4_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__0__4_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__0__4_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__0__4_top_grid_pin_31_[0]),
		.bottom_grid_pin_0_(cbx_1__0__4_bottom_grid_pin_0_[0]),
		.ccff_tail(cbx_1__0__4_ccff_tail[0]));

	cbx_1__0_ cbx_6__0_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__0__4_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__0__5_chanx_left_out[0:19]),
		.ccff_head(sb_1__0__5_ccff_tail[0]),
		.chanx_left_out(cbx_1__0__5_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__0__5_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__0__5_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__0__5_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__0__5_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__0__5_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__0__5_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__0__5_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__0__5_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__0__5_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__0__5_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__0__5_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__0__5_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__0__5_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__0__5_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__0__5_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__0__5_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__0__5_top_grid_pin_31_[0]),
		.bottom_grid_pin_0_(cbx_1__0__5_bottom_grid_pin_0_[0]),
		.ccff_tail(cbx_1__0__5_ccff_tail[0]));

	cbx_1__0_ cbx_7__0_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__0__5_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__0__6_chanx_left_out[0:19]),
		.ccff_head(sb_1__0__6_ccff_tail[0]),
		.chanx_left_out(cbx_1__0__6_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__0__6_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__0__6_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__0__6_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__0__6_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__0__6_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__0__6_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__0__6_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__0__6_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__0__6_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__0__6_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__0__6_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__0__6_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__0__6_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__0__6_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__0__6_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__0__6_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__0__6_top_grid_pin_31_[0]),
		.bottom_grid_pin_0_(cbx_1__0__6_bottom_grid_pin_0_[0]),
		.ccff_tail(cbx_1__0__6_ccff_tail[0]));

	cbx_1__0_ cbx_8__0_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__0__6_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__0__7_chanx_left_out[0:19]),
		.ccff_head(sb_1__0__7_ccff_tail[0]),
		.chanx_left_out(cbx_1__0__7_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__0__7_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__0__7_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__0__7_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__0__7_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__0__7_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__0__7_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__0__7_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__0__7_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__0__7_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__0__7_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__0__7_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__0__7_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__0__7_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__0__7_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__0__7_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__0__7_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__0__7_top_grid_pin_31_[0]),
		.bottom_grid_pin_0_(cbx_1__0__7_bottom_grid_pin_0_[0]),
		.ccff_tail(cbx_1__0__7_ccff_tail[0]));

	cbx_1__0_ cbx_9__0_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__0__7_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__0__8_chanx_left_out[0:19]),
		.ccff_head(sb_1__0__8_ccff_tail[0]),
		.chanx_left_out(cbx_1__0__8_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__0__8_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__0__8_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__0__8_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__0__8_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__0__8_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__0__8_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__0__8_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__0__8_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__0__8_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__0__8_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__0__8_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__0__8_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__0__8_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__0__8_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__0__8_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__0__8_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__0__8_top_grid_pin_31_[0]),
		.bottom_grid_pin_0_(cbx_1__0__8_bottom_grid_pin_0_[0]),
		.ccff_tail(cbx_1__0__8_ccff_tail[0]));

	cbx_1__0_ cbx_10__0_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__0__8_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__0__9_chanx_left_out[0:19]),
		.ccff_head(sb_1__0__9_ccff_tail[0]),
		.chanx_left_out(cbx_1__0__9_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__0__9_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__0__9_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__0__9_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__0__9_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__0__9_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__0__9_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__0__9_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__0__9_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__0__9_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__0__9_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__0__9_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__0__9_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__0__9_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__0__9_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__0__9_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__0__9_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__0__9_top_grid_pin_31_[0]),
		.bottom_grid_pin_0_(cbx_1__0__9_bottom_grid_pin_0_[0]),
		.ccff_tail(cbx_1__0__9_ccff_tail[0]));

	cbx_1__0_ cbx_11__0_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__0__9_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__0__10_chanx_left_out[0:19]),
		.ccff_head(sb_1__0__10_ccff_tail[0]),
		.chanx_left_out(cbx_1__0__10_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__0__10_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__0__10_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__0__10_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__0__10_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__0__10_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__0__10_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__0__10_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__0__10_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__0__10_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__0__10_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__0__10_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__0__10_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__0__10_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__0__10_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__0__10_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__0__10_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__0__10_top_grid_pin_31_[0]),
		.bottom_grid_pin_0_(cbx_1__0__10_bottom_grid_pin_0_[0]),
		.ccff_tail(cbx_1__0__10_ccff_tail[0]));

	cbx_1__0_ cbx_12__0_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__0__10_chanx_right_out[0:19]),
		.chanx_right_in(sb_12__0__0_chanx_left_out[0:19]),
		.ccff_head(sb_12__0__0_ccff_tail[0]),
		.chanx_left_out(cbx_1__0__11_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__0__11_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__0__11_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__0__11_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__0__11_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__0__11_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__0__11_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__0__11_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__0__11_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__0__11_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__0__11_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__0__11_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__0__11_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__0__11_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__0__11_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__0__11_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__0__11_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__0__11_top_grid_pin_31_[0]),
		.bottom_grid_pin_0_(cbx_1__0__11_bottom_grid_pin_0_[0]),
		.ccff_tail(cbx_1__0__11_ccff_tail[0]));

	cbx_1__1_ cbx_1__1_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_0__1__0_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__0_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__0_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__0_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__0_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__0_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__0_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__0_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__0_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__0_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__0_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__0_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__0_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__0_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__0_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__0_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__0_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__0_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__0_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__0_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__0_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__0_ccff_tail[0]));

	cbx_1__1_ cbx_1__2_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_0__1__1_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__1_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__1_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__1_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__1_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__1_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__1_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__1_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__1_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__1_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__1_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__1_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__1_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__1_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__1_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__1_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__1_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__1_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__1_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__1_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__1_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__1_ccff_tail[0]));

	cbx_1__1_ cbx_1__3_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_0__1__2_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__2_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__2_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__2_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__2_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__2_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__2_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__2_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__2_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__2_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__2_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__2_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__2_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__2_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__2_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__2_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__2_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__2_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__2_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__2_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__2_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__2_ccff_tail[0]));

	cbx_1__1_ cbx_1__4_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_0__1__3_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__3_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__3_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__3_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__3_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__3_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__3_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__3_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__3_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__3_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__3_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__3_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__3_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__3_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__3_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__3_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__3_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__3_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__3_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__3_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__3_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__3_ccff_tail[0]));

	cbx_1__1_ cbx_1__5_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_0__1__4_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__4_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__4_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__4_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__4_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__4_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__4_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__4_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__4_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__4_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__4_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__4_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__4_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__4_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__4_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__4_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__4_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__4_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__4_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__4_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__4_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__4_ccff_tail[0]));

	cbx_1__1_ cbx_1__6_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_0__1__5_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__5_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__5_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__5_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__5_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__5_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__5_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__5_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__5_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__5_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__5_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__5_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__5_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__5_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__5_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__5_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__5_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__5_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__5_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__5_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__5_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__5_ccff_tail[0]));

	cbx_1__1_ cbx_1__7_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_0__1__6_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__6_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__6_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__6_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__6_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__6_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__6_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__6_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__6_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__6_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__6_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__6_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__6_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__6_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__6_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__6_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__6_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__6_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__6_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__6_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__6_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__6_ccff_tail[0]));

	cbx_1__1_ cbx_1__8_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_0__1__7_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__7_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__7_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__7_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__7_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__7_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__7_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__7_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__7_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__7_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__7_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__7_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__7_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__7_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__7_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__7_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__7_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__7_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__7_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__7_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__7_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__7_ccff_tail[0]));

	cbx_1__1_ cbx_1__9_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_0__1__8_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__8_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__8_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__8_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__8_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__8_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__8_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__8_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__8_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__8_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__8_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__8_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__8_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__8_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__8_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__8_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__8_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__8_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__8_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__8_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__8_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__8_ccff_tail[0]));

	cbx_1__1_ cbx_1__10_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_0__1__9_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__9_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__9_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__9_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__9_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__9_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__9_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__9_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__9_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__9_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__9_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__9_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__9_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__9_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__9_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__9_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__9_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__9_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__9_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__9_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__9_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__9_ccff_tail[0]));

	cbx_1__1_ cbx_1__11_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_0__1__10_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__10_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__10_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__10_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__10_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__10_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__10_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__10_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__10_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__10_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__10_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__10_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__10_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__10_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__10_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__10_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__10_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__10_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__10_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__10_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__10_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__10_ccff_tail[0]));

	cbx_1__1_ cbx_2__1_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__0_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__11_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__11_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__11_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__11_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__11_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__11_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__11_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__11_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__11_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__11_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__11_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__11_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__11_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__11_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__11_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__11_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__11_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__11_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__11_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__11_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__11_ccff_tail[0]));

	cbx_1__1_ cbx_2__2_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__1_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__12_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__12_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__12_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__12_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__12_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__12_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__12_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__12_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__12_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__12_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__12_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__12_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__12_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__12_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__12_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__12_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__12_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__12_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__12_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__12_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__12_ccff_tail[0]));

	cbx_1__1_ cbx_2__3_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__2_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__13_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__13_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__13_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__13_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__13_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__13_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__13_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__13_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__13_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__13_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__13_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__13_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__13_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__13_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__13_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__13_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__13_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__13_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__13_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__13_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__13_ccff_tail[0]));

	cbx_1__1_ cbx_2__4_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__3_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__14_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__14_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__14_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__14_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__14_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__14_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__14_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__14_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__14_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__14_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__14_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__14_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__14_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__14_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__14_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__14_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__14_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__14_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__14_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__14_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__14_ccff_tail[0]));

	cbx_1__1_ cbx_2__5_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__4_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__15_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__15_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__15_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__15_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__15_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__15_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__15_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__15_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__15_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__15_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__15_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__15_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__15_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__15_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__15_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__15_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__15_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__15_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__15_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__15_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__15_ccff_tail[0]));

	cbx_1__1_ cbx_2__6_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__5_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__16_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__16_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__16_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__16_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__16_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__16_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__16_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__16_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__16_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__16_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__16_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__16_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__16_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__16_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__16_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__16_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__16_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__16_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__16_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__16_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__16_ccff_tail[0]));

	cbx_1__1_ cbx_2__7_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__6_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__17_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__17_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__17_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__17_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__17_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__17_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__17_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__17_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__17_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__17_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__17_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__17_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__17_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__17_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__17_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__17_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__17_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__17_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__17_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__17_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__17_ccff_tail[0]));

	cbx_1__1_ cbx_2__8_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__7_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__18_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__18_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__18_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__18_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__18_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__18_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__18_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__18_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__18_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__18_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__18_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__18_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__18_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__18_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__18_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__18_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__18_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__18_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__18_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__18_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__18_ccff_tail[0]));

	cbx_1__1_ cbx_2__9_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__8_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__19_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__19_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__19_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__19_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__19_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__19_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__19_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__19_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__19_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__19_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__19_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__19_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__19_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__19_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__19_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__19_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__19_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__19_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__19_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__19_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__19_ccff_tail[0]));

	cbx_1__1_ cbx_2__10_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__9_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__20_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__20_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__20_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__20_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__20_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__20_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__20_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__20_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__20_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__20_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__20_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__20_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__20_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__20_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__20_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__20_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__20_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__20_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__20_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__20_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__20_ccff_tail[0]));

	cbx_1__1_ cbx_2__11_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__10_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__21_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__21_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__21_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__21_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__21_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__21_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__21_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__21_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__21_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__21_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__21_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__21_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__21_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__21_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__21_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__21_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__21_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__21_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__21_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__21_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__21_ccff_tail[0]));

	cbx_1__1_ cbx_3__1_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__11_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__22_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__22_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__22_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__22_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__22_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__22_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__22_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__22_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__22_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__22_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__22_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__22_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__22_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__22_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__22_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__22_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__22_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__22_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__22_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__22_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__22_ccff_tail[0]));

	cbx_1__1_ cbx_3__2_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__12_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__23_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__23_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__23_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__23_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__23_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__23_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__23_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__23_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__23_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__23_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__23_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__23_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__23_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__23_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__23_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__23_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__23_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__23_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__23_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__23_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__23_ccff_tail[0]));

	cbx_1__1_ cbx_3__3_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__13_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__24_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__24_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__24_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__24_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__24_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__24_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__24_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__24_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__24_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__24_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__24_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__24_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__24_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__24_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__24_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__24_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__24_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__24_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__24_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__24_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__24_ccff_tail[0]));

	cbx_1__1_ cbx_3__4_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__14_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__25_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__25_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__25_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__25_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__25_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__25_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__25_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__25_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__25_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__25_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__25_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__25_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__25_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__25_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__25_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__25_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__25_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__25_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__25_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__25_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__25_ccff_tail[0]));

	cbx_1__1_ cbx_3__5_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__15_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__26_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__26_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__26_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__26_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__26_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__26_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__26_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__26_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__26_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__26_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__26_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__26_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__26_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__26_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__26_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__26_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__26_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__26_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__26_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__26_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__26_ccff_tail[0]));

	cbx_1__1_ cbx_3__6_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__16_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__27_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__27_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__27_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__27_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__27_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__27_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__27_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__27_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__27_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__27_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__27_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__27_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__27_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__27_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__27_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__27_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__27_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__27_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__27_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__27_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__27_ccff_tail[0]));

	cbx_1__1_ cbx_3__7_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__17_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__28_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__28_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__28_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__28_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__28_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__28_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__28_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__28_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__28_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__28_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__28_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__28_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__28_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__28_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__28_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__28_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__28_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__28_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__28_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__28_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__28_ccff_tail[0]));

	cbx_1__1_ cbx_3__8_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__18_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__29_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__29_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__29_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__29_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__29_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__29_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__29_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__29_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__29_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__29_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__29_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__29_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__29_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__29_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__29_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__29_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__29_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__29_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__29_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__29_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__29_ccff_tail[0]));

	cbx_1__1_ cbx_3__9_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__19_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__30_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__30_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__30_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__30_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__30_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__30_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__30_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__30_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__30_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__30_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__30_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__30_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__30_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__30_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__30_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__30_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__30_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__30_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__30_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__30_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__30_ccff_tail[0]));

	cbx_1__1_ cbx_3__10_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__20_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__31_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__31_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__31_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__31_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__31_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__31_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__31_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__31_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__31_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__31_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__31_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__31_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__31_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__31_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__31_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__31_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__31_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__31_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__31_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__31_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__31_ccff_tail[0]));

	cbx_1__1_ cbx_3__11_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__21_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__32_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__32_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__32_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__32_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__32_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__32_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__32_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__32_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__32_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__32_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__32_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__32_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__32_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__32_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__32_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__32_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__32_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__32_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__32_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__32_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__32_ccff_tail[0]));

	cbx_1__1_ cbx_4__1_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__22_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__33_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__33_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__33_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__33_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__33_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__33_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__33_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__33_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__33_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__33_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__33_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__33_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__33_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__33_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__33_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__33_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__33_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__33_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__33_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__33_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__33_ccff_tail[0]));

	cbx_1__1_ cbx_4__2_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__23_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__34_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__34_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__34_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__34_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__34_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__34_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__34_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__34_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__34_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__34_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__34_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__34_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__34_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__34_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__34_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__34_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__34_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__34_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__34_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__34_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__34_ccff_tail[0]));

	cbx_1__1_ cbx_4__3_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__24_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__35_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__35_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__35_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__35_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__35_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__35_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__35_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__35_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__35_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__35_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__35_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__35_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__35_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__35_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__35_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__35_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__35_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__35_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__35_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__35_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__35_ccff_tail[0]));

	cbx_1__1_ cbx_4__4_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__25_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__36_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__36_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__36_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__36_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__36_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__36_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__36_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__36_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__36_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__36_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__36_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__36_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__36_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__36_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__36_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__36_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__36_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__36_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__36_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__36_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__36_ccff_tail[0]));

	cbx_1__1_ cbx_4__5_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__26_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__37_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__37_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__37_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__37_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__37_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__37_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__37_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__37_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__37_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__37_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__37_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__37_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__37_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__37_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__37_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__37_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__37_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__37_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__37_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__37_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__37_ccff_tail[0]));

	cbx_1__1_ cbx_4__6_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__27_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__38_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__38_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__38_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__38_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__38_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__38_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__38_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__38_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__38_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__38_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__38_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__38_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__38_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__38_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__38_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__38_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__38_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__38_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__38_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__38_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__38_ccff_tail[0]));

	cbx_1__1_ cbx_4__7_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__28_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__39_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__39_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__39_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__39_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__39_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__39_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__39_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__39_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__39_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__39_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__39_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__39_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__39_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__39_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__39_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__39_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__39_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__39_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__39_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__39_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__39_ccff_tail[0]));

	cbx_1__1_ cbx_4__8_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__29_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__40_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__40_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__40_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__40_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__40_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__40_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__40_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__40_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__40_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__40_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__40_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__40_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__40_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__40_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__40_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__40_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__40_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__40_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__40_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__40_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__40_ccff_tail[0]));

	cbx_1__1_ cbx_4__9_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__30_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__41_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__41_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__41_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__41_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__41_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__41_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__41_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__41_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__41_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__41_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__41_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__41_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__41_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__41_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__41_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__41_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__41_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__41_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__41_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__41_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__41_ccff_tail[0]));

	cbx_1__1_ cbx_4__10_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__31_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__42_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__42_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__42_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__42_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__42_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__42_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__42_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__42_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__42_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__42_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__42_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__42_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__42_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__42_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__42_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__42_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__42_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__42_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__42_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__42_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__42_ccff_tail[0]));

	cbx_1__1_ cbx_4__11_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__32_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__43_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__43_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__43_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__43_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__43_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__43_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__43_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__43_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__43_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__43_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__43_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__43_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__43_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__43_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__43_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__43_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__43_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__43_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__43_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__43_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__43_ccff_tail[0]));

	cbx_1__1_ cbx_5__1_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__33_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__44_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__44_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__44_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__44_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__44_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__44_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__44_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__44_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__44_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__44_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__44_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__44_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__44_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__44_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__44_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__44_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__44_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__44_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__44_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__44_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__44_ccff_tail[0]));

	cbx_1__1_ cbx_5__2_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__34_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__45_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__45_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__45_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__45_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__45_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__45_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__45_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__45_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__45_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__45_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__45_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__45_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__45_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__45_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__45_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__45_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__45_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__45_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__45_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__45_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__45_ccff_tail[0]));

	cbx_1__1_ cbx_5__3_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__35_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__46_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__46_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__46_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__46_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__46_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__46_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__46_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__46_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__46_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__46_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__46_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__46_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__46_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__46_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__46_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__46_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__46_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__46_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__46_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__46_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__46_ccff_tail[0]));

	cbx_1__1_ cbx_5__4_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__36_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__47_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__47_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__47_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__47_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__47_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__47_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__47_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__47_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__47_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__47_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__47_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__47_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__47_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__47_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__47_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__47_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__47_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__47_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__47_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__47_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__47_ccff_tail[0]));

	cbx_1__1_ cbx_5__5_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__37_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__48_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__48_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__48_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__48_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__48_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__48_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__48_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__48_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__48_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__48_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__48_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__48_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__48_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__48_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__48_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__48_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__48_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__48_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__48_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__48_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__48_ccff_tail[0]));

	cbx_1__1_ cbx_5__6_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__38_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__49_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__49_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__49_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__49_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__49_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__49_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__49_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__49_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__49_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__49_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__49_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__49_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__49_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__49_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__49_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__49_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__49_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__49_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__49_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__49_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__49_ccff_tail[0]));

	cbx_1__1_ cbx_5__7_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__39_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__50_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__50_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__50_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__50_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__50_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__50_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__50_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__50_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__50_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__50_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__50_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__50_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__50_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__50_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__50_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__50_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__50_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__50_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__50_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__50_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__50_ccff_tail[0]));

	cbx_1__1_ cbx_5__8_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__40_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__51_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__51_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__51_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__51_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__51_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__51_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__51_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__51_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__51_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__51_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__51_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__51_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__51_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__51_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__51_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__51_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__51_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__51_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__51_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__51_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__51_ccff_tail[0]));

	cbx_1__1_ cbx_5__9_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__41_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__52_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__52_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__52_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__52_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__52_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__52_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__52_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__52_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__52_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__52_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__52_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__52_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__52_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__52_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__52_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__52_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__52_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__52_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__52_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__52_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__52_ccff_tail[0]));

	cbx_1__1_ cbx_5__10_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__42_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__53_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__53_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__53_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__53_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__53_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__53_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__53_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__53_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__53_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__53_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__53_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__53_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__53_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__53_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__53_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__53_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__53_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__53_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__53_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__53_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__53_ccff_tail[0]));

	cbx_1__1_ cbx_5__11_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__43_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__54_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__54_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__54_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__54_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__54_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__54_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__54_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__54_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__54_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__54_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__54_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__54_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__54_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__54_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__54_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__54_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__54_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__54_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__54_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__54_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__54_ccff_tail[0]));

	cbx_1__1_ cbx_6__1_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__44_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__55_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__55_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__55_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__55_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__55_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__55_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__55_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__55_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__55_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__55_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__55_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__55_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__55_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__55_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__55_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__55_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__55_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__55_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__55_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__55_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__55_ccff_tail[0]));

	cbx_1__1_ cbx_6__2_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__45_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__56_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__56_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__56_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__56_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__56_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__56_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__56_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__56_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__56_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__56_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__56_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__56_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__56_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__56_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__56_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__56_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__56_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__56_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__56_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__56_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__56_ccff_tail[0]));

	cbx_1__1_ cbx_6__3_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__46_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__57_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__57_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__57_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__57_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__57_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__57_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__57_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__57_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__57_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__57_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__57_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__57_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__57_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__57_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__57_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__57_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__57_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__57_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__57_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__57_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__57_ccff_tail[0]));

	cbx_1__1_ cbx_6__4_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__47_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__58_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__58_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__58_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__58_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__58_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__58_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__58_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__58_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__58_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__58_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__58_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__58_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__58_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__58_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__58_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__58_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__58_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__58_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__58_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__58_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__58_ccff_tail[0]));

	cbx_1__1_ cbx_6__5_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__48_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__59_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__59_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__59_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__59_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__59_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__59_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__59_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__59_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__59_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__59_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__59_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__59_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__59_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__59_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__59_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__59_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__59_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__59_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__59_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__59_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__59_ccff_tail[0]));

	cbx_1__1_ cbx_6__6_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__49_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__60_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__60_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__60_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__60_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__60_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__60_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__60_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__60_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__60_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__60_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__60_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__60_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__60_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__60_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__60_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__60_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__60_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__60_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__60_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__60_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__60_ccff_tail[0]));

	cbx_1__1_ cbx_6__7_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__50_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__61_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__61_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__61_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__61_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__61_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__61_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__61_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__61_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__61_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__61_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__61_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__61_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__61_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__61_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__61_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__61_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__61_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__61_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__61_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__61_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__61_ccff_tail[0]));

	cbx_1__1_ cbx_6__8_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__51_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__62_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__62_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__62_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__62_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__62_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__62_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__62_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__62_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__62_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__62_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__62_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__62_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__62_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__62_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__62_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__62_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__62_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__62_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__62_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__62_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__62_ccff_tail[0]));

	cbx_1__1_ cbx_6__9_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__52_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__63_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__63_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__63_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__63_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__63_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__63_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__63_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__63_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__63_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__63_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__63_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__63_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__63_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__63_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__63_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__63_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__63_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__63_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__63_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__63_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__63_ccff_tail[0]));

	cbx_1__1_ cbx_6__10_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__53_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__64_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__64_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__64_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__64_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__64_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__64_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__64_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__64_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__64_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__64_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__64_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__64_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__64_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__64_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__64_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__64_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__64_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__64_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__64_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__64_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__64_ccff_tail[0]));

	cbx_1__1_ cbx_6__11_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__54_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__65_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__65_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__65_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__65_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__65_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__65_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__65_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__65_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__65_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__65_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__65_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__65_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__65_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__65_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__65_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__65_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__65_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__65_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__65_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__65_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__65_ccff_tail[0]));

	cbx_1__1_ cbx_7__1_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__55_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__66_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__66_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__66_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__66_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__66_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__66_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__66_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__66_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__66_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__66_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__66_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__66_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__66_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__66_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__66_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__66_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__66_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__66_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__66_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__66_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__66_ccff_tail[0]));

	cbx_1__1_ cbx_7__2_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__56_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__67_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__67_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__67_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__67_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__67_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__67_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__67_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__67_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__67_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__67_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__67_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__67_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__67_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__67_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__67_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__67_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__67_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__67_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__67_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__67_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__67_ccff_tail[0]));

	cbx_1__1_ cbx_7__3_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__57_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__68_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__68_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__68_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__68_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__68_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__68_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__68_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__68_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__68_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__68_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__68_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__68_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__68_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__68_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__68_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__68_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__68_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__68_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__68_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__68_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__68_ccff_tail[0]));

	cbx_1__1_ cbx_7__4_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__58_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__69_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__69_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__69_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__69_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__69_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__69_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__69_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__69_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__69_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__69_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__69_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__69_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__69_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__69_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__69_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__69_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__69_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__69_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__69_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__69_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__69_ccff_tail[0]));

	cbx_1__1_ cbx_7__5_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__59_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__70_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__70_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__70_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__70_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__70_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__70_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__70_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__70_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__70_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__70_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__70_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__70_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__70_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__70_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__70_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__70_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__70_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__70_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__70_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__70_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__70_ccff_tail[0]));

	cbx_1__1_ cbx_7__6_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__60_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__71_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__71_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__71_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__71_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__71_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__71_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__71_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__71_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__71_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__71_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__71_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__71_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__71_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__71_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__71_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__71_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__71_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__71_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__71_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__71_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__71_ccff_tail[0]));

	cbx_1__1_ cbx_7__7_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__61_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__72_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__72_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__72_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__72_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__72_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__72_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__72_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__72_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__72_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__72_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__72_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__72_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__72_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__72_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__72_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__72_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__72_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__72_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__72_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__72_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__72_ccff_tail[0]));

	cbx_1__1_ cbx_7__8_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__62_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__73_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__73_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__73_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__73_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__73_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__73_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__73_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__73_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__73_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__73_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__73_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__73_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__73_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__73_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__73_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__73_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__73_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__73_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__73_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__73_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__73_ccff_tail[0]));

	cbx_1__1_ cbx_7__9_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__63_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__74_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__74_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__74_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__74_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__74_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__74_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__74_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__74_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__74_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__74_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__74_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__74_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__74_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__74_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__74_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__74_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__74_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__74_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__74_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__74_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__74_ccff_tail[0]));

	cbx_1__1_ cbx_7__10_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__64_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__75_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__75_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__75_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__75_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__75_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__75_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__75_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__75_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__75_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__75_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__75_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__75_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__75_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__75_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__75_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__75_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__75_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__75_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__75_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__75_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__75_ccff_tail[0]));

	cbx_1__1_ cbx_7__11_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__65_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__76_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__76_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__76_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__76_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__76_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__76_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__76_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__76_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__76_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__76_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__76_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__76_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__76_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__76_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__76_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__76_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__76_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__76_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__76_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__76_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__76_ccff_tail[0]));

	cbx_1__1_ cbx_8__1_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__66_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__77_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__77_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__77_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__77_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__77_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__77_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__77_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__77_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__77_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__77_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__77_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__77_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__77_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__77_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__77_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__77_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__77_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__77_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__77_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__77_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__77_ccff_tail[0]));

	cbx_1__1_ cbx_8__2_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__67_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__78_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__78_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__78_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__78_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__78_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__78_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__78_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__78_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__78_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__78_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__78_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__78_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__78_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__78_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__78_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__78_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__78_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__78_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__78_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__78_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__78_ccff_tail[0]));

	cbx_1__1_ cbx_8__3_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__68_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__79_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__79_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__79_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__79_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__79_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__79_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__79_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__79_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__79_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__79_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__79_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__79_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__79_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__79_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__79_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__79_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__79_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__79_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__79_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__79_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__79_ccff_tail[0]));

	cbx_1__1_ cbx_8__4_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__69_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__80_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__80_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__80_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__80_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__80_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__80_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__80_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__80_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__80_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__80_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__80_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__80_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__80_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__80_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__80_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__80_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__80_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__80_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__80_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__80_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__80_ccff_tail[0]));

	cbx_1__1_ cbx_8__5_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__70_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__81_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__81_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__81_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__81_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__81_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__81_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__81_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__81_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__81_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__81_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__81_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__81_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__81_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__81_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__81_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__81_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__81_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__81_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__81_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__81_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__81_ccff_tail[0]));

	cbx_1__1_ cbx_8__6_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__71_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__82_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__82_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__82_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__82_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__82_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__82_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__82_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__82_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__82_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__82_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__82_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__82_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__82_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__82_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__82_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__82_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__82_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__82_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__82_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__82_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__82_ccff_tail[0]));

	cbx_1__1_ cbx_8__7_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__72_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__83_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__83_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__83_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__83_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__83_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__83_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__83_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__83_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__83_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__83_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__83_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__83_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__83_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__83_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__83_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__83_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__83_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__83_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__83_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__83_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__83_ccff_tail[0]));

	cbx_1__1_ cbx_8__8_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__73_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__84_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__84_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__84_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__84_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__84_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__84_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__84_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__84_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__84_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__84_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__84_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__84_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__84_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__84_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__84_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__84_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__84_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__84_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__84_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__84_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__84_ccff_tail[0]));

	cbx_1__1_ cbx_8__9_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__74_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__85_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__85_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__85_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__85_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__85_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__85_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__85_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__85_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__85_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__85_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__85_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__85_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__85_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__85_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__85_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__85_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__85_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__85_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__85_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__85_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__85_ccff_tail[0]));

	cbx_1__1_ cbx_8__10_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__75_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__86_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__86_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__86_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__86_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__86_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__86_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__86_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__86_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__86_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__86_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__86_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__86_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__86_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__86_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__86_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__86_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__86_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__86_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__86_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__86_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__86_ccff_tail[0]));

	cbx_1__1_ cbx_8__11_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__76_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__87_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__87_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__87_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__87_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__87_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__87_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__87_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__87_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__87_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__87_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__87_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__87_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__87_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__87_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__87_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__87_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__87_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__87_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__87_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__87_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__87_ccff_tail[0]));

	cbx_1__1_ cbx_9__1_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__77_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__88_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__88_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__88_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__88_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__88_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__88_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__88_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__88_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__88_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__88_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__88_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__88_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__88_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__88_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__88_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__88_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__88_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__88_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__88_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__88_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__88_ccff_tail[0]));

	cbx_1__1_ cbx_9__2_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__78_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__89_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__89_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__89_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__89_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__89_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__89_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__89_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__89_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__89_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__89_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__89_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__89_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__89_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__89_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__89_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__89_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__89_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__89_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__89_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__89_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__89_ccff_tail[0]));

	cbx_1__1_ cbx_9__3_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__79_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__90_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__90_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__90_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__90_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__90_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__90_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__90_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__90_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__90_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__90_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__90_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__90_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__90_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__90_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__90_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__90_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__90_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__90_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__90_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__90_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__90_ccff_tail[0]));

	cbx_1__1_ cbx_9__4_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__80_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__91_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__91_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__91_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__91_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__91_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__91_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__91_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__91_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__91_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__91_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__91_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__91_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__91_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__91_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__91_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__91_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__91_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__91_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__91_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__91_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__91_ccff_tail[0]));

	cbx_1__1_ cbx_9__5_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__81_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__92_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__92_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__92_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__92_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__92_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__92_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__92_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__92_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__92_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__92_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__92_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__92_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__92_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__92_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__92_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__92_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__92_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__92_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__92_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__92_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__92_ccff_tail[0]));

	cbx_1__1_ cbx_9__6_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__82_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__93_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__93_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__93_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__93_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__93_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__93_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__93_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__93_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__93_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__93_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__93_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__93_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__93_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__93_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__93_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__93_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__93_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__93_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__93_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__93_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__93_ccff_tail[0]));

	cbx_1__1_ cbx_9__7_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__83_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__94_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__94_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__94_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__94_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__94_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__94_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__94_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__94_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__94_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__94_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__94_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__94_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__94_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__94_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__94_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__94_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__94_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__94_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__94_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__94_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__94_ccff_tail[0]));

	cbx_1__1_ cbx_9__8_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__84_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__95_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__95_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__95_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__95_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__95_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__95_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__95_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__95_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__95_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__95_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__95_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__95_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__95_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__95_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__95_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__95_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__95_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__95_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__95_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__95_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__95_ccff_tail[0]));

	cbx_1__1_ cbx_9__9_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__85_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__96_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__96_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__96_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__96_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__96_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__96_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__96_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__96_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__96_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__96_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__96_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__96_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__96_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__96_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__96_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__96_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__96_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__96_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__96_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__96_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__96_ccff_tail[0]));

	cbx_1__1_ cbx_9__10_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__86_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__97_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__97_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__97_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__97_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__97_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__97_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__97_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__97_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__97_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__97_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__97_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__97_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__97_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__97_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__97_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__97_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__97_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__97_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__97_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__97_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__97_ccff_tail[0]));

	cbx_1__1_ cbx_9__11_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__87_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__98_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__98_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__98_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__98_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__98_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__98_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__98_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__98_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__98_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__98_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__98_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__98_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__98_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__98_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__98_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__98_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__98_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__98_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__98_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__98_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__98_ccff_tail[0]));

	cbx_1__1_ cbx_10__1_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__88_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__99_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__99_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__99_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__99_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__99_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__99_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__99_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__99_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__99_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__99_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__99_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__99_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__99_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__99_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__99_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__99_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__99_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__99_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__99_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__99_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__99_ccff_tail[0]));

	cbx_1__1_ cbx_10__2_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__89_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__100_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__100_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__100_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__100_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__100_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__100_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__100_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__100_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__100_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__100_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__100_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__100_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__100_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__100_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__100_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__100_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__100_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__100_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__100_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__100_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__100_ccff_tail[0]));

	cbx_1__1_ cbx_10__3_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__90_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__101_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__101_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__101_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__101_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__101_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__101_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__101_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__101_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__101_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__101_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__101_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__101_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__101_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__101_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__101_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__101_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__101_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__101_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__101_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__101_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__101_ccff_tail[0]));

	cbx_1__1_ cbx_10__4_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__91_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__102_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__102_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__102_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__102_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__102_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__102_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__102_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__102_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__102_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__102_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__102_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__102_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__102_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__102_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__102_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__102_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__102_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__102_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__102_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__102_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__102_ccff_tail[0]));

	cbx_1__1_ cbx_10__5_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__92_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__103_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__103_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__103_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__103_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__103_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__103_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__103_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__103_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__103_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__103_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__103_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__103_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__103_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__103_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__103_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__103_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__103_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__103_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__103_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__103_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__103_ccff_tail[0]));

	cbx_1__1_ cbx_10__6_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__93_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__104_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__104_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__104_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__104_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__104_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__104_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__104_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__104_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__104_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__104_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__104_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__104_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__104_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__104_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__104_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__104_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__104_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__104_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__104_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__104_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__104_ccff_tail[0]));

	cbx_1__1_ cbx_10__7_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__94_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__105_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__105_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__105_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__105_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__105_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__105_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__105_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__105_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__105_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__105_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__105_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__105_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__105_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__105_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__105_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__105_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__105_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__105_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__105_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__105_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__105_ccff_tail[0]));

	cbx_1__1_ cbx_10__8_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__95_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__106_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__106_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__106_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__106_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__106_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__106_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__106_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__106_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__106_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__106_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__106_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__106_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__106_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__106_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__106_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__106_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__106_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__106_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__106_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__106_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__106_ccff_tail[0]));

	cbx_1__1_ cbx_10__9_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__96_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__107_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__107_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__107_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__107_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__107_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__107_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__107_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__107_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__107_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__107_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__107_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__107_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__107_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__107_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__107_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__107_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__107_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__107_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__107_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__107_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__107_ccff_tail[0]));

	cbx_1__1_ cbx_10__10_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__97_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__108_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__108_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__108_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__108_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__108_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__108_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__108_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__108_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__108_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__108_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__108_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__108_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__108_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__108_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__108_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__108_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__108_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__108_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__108_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__108_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__108_ccff_tail[0]));

	cbx_1__1_ cbx_10__11_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__98_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__109_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__109_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__109_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__109_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__109_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__109_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__109_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__109_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__109_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__109_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__109_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__109_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__109_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__109_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__109_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__109_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__109_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__109_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__109_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__109_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__109_ccff_tail[0]));

	cbx_1__1_ cbx_11__1_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__99_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__110_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__110_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__110_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__110_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__110_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__110_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__110_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__110_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__110_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__110_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__110_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__110_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__110_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__110_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__110_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__110_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__110_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__110_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__110_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__110_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__110_ccff_tail[0]));

	cbx_1__1_ cbx_11__2_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__100_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__111_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__111_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__111_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__111_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__111_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__111_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__111_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__111_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__111_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__111_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__111_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__111_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__111_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__111_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__111_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__111_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__111_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__111_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__111_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__111_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__111_ccff_tail[0]));

	cbx_1__1_ cbx_11__3_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__101_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__112_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__112_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__112_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__112_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__112_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__112_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__112_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__112_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__112_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__112_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__112_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__112_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__112_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__112_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__112_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__112_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__112_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__112_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__112_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__112_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__112_ccff_tail[0]));

	cbx_1__1_ cbx_11__4_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__102_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__113_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__113_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__113_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__113_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__113_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__113_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__113_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__113_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__113_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__113_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__113_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__113_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__113_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__113_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__113_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__113_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__113_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__113_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__113_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__113_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__113_ccff_tail[0]));

	cbx_1__1_ cbx_11__5_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__103_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__114_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__114_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__114_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__114_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__114_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__114_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__114_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__114_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__114_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__114_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__114_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__114_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__114_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__114_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__114_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__114_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__114_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__114_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__114_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__114_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__114_ccff_tail[0]));

	cbx_1__1_ cbx_11__6_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__104_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__115_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__115_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__115_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__115_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__115_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__115_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__115_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__115_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__115_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__115_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__115_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__115_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__115_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__115_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__115_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__115_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__115_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__115_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__115_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__115_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__115_ccff_tail[0]));

	cbx_1__1_ cbx_11__7_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__105_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__116_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__116_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__116_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__116_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__116_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__116_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__116_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__116_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__116_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__116_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__116_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__116_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__116_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__116_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__116_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__116_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__116_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__116_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__116_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__116_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__116_ccff_tail[0]));

	cbx_1__1_ cbx_11__8_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__106_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__117_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__117_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__117_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__117_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__117_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__117_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__117_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__117_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__117_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__117_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__117_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__117_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__117_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__117_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__117_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__117_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__117_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__117_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__117_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__117_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__117_ccff_tail[0]));

	cbx_1__1_ cbx_11__9_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__107_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__118_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__118_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__118_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__118_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__118_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__118_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__118_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__118_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__118_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__118_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__118_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__118_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__118_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__118_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__118_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__118_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__118_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__118_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__118_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__118_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__118_ccff_tail[0]));

	cbx_1__1_ cbx_11__10_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__108_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__119_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__119_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__119_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__119_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__119_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__119_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__119_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__119_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__119_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__119_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__119_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__119_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__119_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__119_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__119_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__119_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__119_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__119_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__119_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__119_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__119_ccff_tail[0]));

	cbx_1__1_ cbx_11__11_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__109_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__120_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__120_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__120_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__120_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__120_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__120_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__120_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__120_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__120_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__120_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__120_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__120_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__120_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__120_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__120_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__120_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__120_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__120_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__120_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__120_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__120_ccff_tail[0]));

	cbx_1__1_ cbx_12__1_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__110_chanx_right_out[0:19]),
		.chanx_right_in(sb_12__1__0_chanx_left_out[0:19]),
		.ccff_head(sb_12__1__0_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__121_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__121_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__121_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__121_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__121_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__121_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__121_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__121_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__121_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__121_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__121_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__121_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__121_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__121_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__121_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__121_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__121_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__121_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__121_ccff_tail[0]));

	cbx_1__1_ cbx_12__2_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__111_chanx_right_out[0:19]),
		.chanx_right_in(sb_12__1__1_chanx_left_out[0:19]),
		.ccff_head(sb_12__1__1_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__122_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__122_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__122_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__122_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__122_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__122_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__122_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__122_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__122_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__122_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__122_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__122_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__122_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__122_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__122_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__122_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__122_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__122_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__122_ccff_tail[0]));

	cbx_1__1_ cbx_12__3_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__112_chanx_right_out[0:19]),
		.chanx_right_in(sb_12__1__2_chanx_left_out[0:19]),
		.ccff_head(sb_12__1__2_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__123_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__123_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__123_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__123_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__123_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__123_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__123_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__123_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__123_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__123_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__123_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__123_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__123_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__123_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__123_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__123_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__123_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__123_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__123_ccff_tail[0]));

	cbx_1__1_ cbx_12__4_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__113_chanx_right_out[0:19]),
		.chanx_right_in(sb_12__1__3_chanx_left_out[0:19]),
		.ccff_head(sb_12__1__3_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__124_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__124_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__124_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__124_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__124_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__124_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__124_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__124_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__124_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__124_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__124_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__124_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__124_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__124_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__124_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__124_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__124_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__124_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__124_ccff_tail[0]));

	cbx_1__1_ cbx_12__5_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__114_chanx_right_out[0:19]),
		.chanx_right_in(sb_12__1__4_chanx_left_out[0:19]),
		.ccff_head(sb_12__1__4_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__125_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__125_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__125_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__125_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__125_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__125_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__125_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__125_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__125_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__125_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__125_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__125_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__125_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__125_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__125_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__125_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__125_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__125_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__125_ccff_tail[0]));

	cbx_1__1_ cbx_12__6_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__115_chanx_right_out[0:19]),
		.chanx_right_in(sb_12__1__5_chanx_left_out[0:19]),
		.ccff_head(sb_12__1__5_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__126_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__126_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__126_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__126_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__126_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__126_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__126_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__126_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__126_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__126_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__126_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__126_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__126_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__126_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__126_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__126_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__126_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__126_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__126_ccff_tail[0]));

	cbx_1__1_ cbx_12__7_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__116_chanx_right_out[0:19]),
		.chanx_right_in(sb_12__1__6_chanx_left_out[0:19]),
		.ccff_head(sb_12__1__6_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__127_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__127_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__127_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__127_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__127_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__127_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__127_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__127_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__127_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__127_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__127_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__127_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__127_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__127_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__127_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__127_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__127_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__127_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__127_ccff_tail[0]));

	cbx_1__1_ cbx_12__8_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__117_chanx_right_out[0:19]),
		.chanx_right_in(sb_12__1__7_chanx_left_out[0:19]),
		.ccff_head(sb_12__1__7_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__128_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__128_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__128_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__128_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__128_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__128_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__128_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__128_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__128_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__128_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__128_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__128_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__128_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__128_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__128_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__128_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__128_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__128_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__128_ccff_tail[0]));

	cbx_1__1_ cbx_12__9_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__118_chanx_right_out[0:19]),
		.chanx_right_in(sb_12__1__8_chanx_left_out[0:19]),
		.ccff_head(sb_12__1__8_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__129_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__129_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__129_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__129_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__129_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__129_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__129_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__129_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__129_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__129_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__129_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__129_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__129_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__129_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__129_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__129_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__129_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__129_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__129_ccff_tail[0]));

	cbx_1__1_ cbx_12__10_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__119_chanx_right_out[0:19]),
		.chanx_right_in(sb_12__1__9_chanx_left_out[0:19]),
		.ccff_head(sb_12__1__9_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__130_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__130_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__130_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__130_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__130_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__130_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__130_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__130_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__130_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__130_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__130_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__130_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__130_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__130_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__130_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__130_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__130_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__130_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__130_ccff_tail[0]));

	cbx_1__1_ cbx_12__11_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__1__120_chanx_right_out[0:19]),
		.chanx_right_in(sb_12__1__10_chanx_left_out[0:19]),
		.ccff_head(sb_12__1__10_ccff_tail[0]),
		.chanx_left_out(cbx_1__1__131_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__131_chanx_right_out[0:19]),
		.top_grid_pin_16_(cbx_1__1__131_top_grid_pin_16_[0]),
		.top_grid_pin_17_(cbx_1__1__131_top_grid_pin_17_[0]),
		.top_grid_pin_18_(cbx_1__1__131_top_grid_pin_18_[0]),
		.top_grid_pin_19_(cbx_1__1__131_top_grid_pin_19_[0]),
		.top_grid_pin_20_(cbx_1__1__131_top_grid_pin_20_[0]),
		.top_grid_pin_21_(cbx_1__1__131_top_grid_pin_21_[0]),
		.top_grid_pin_22_(cbx_1__1__131_top_grid_pin_22_[0]),
		.top_grid_pin_23_(cbx_1__1__131_top_grid_pin_23_[0]),
		.top_grid_pin_24_(cbx_1__1__131_top_grid_pin_24_[0]),
		.top_grid_pin_25_(cbx_1__1__131_top_grid_pin_25_[0]),
		.top_grid_pin_26_(cbx_1__1__131_top_grid_pin_26_[0]),
		.top_grid_pin_27_(cbx_1__1__131_top_grid_pin_27_[0]),
		.top_grid_pin_28_(cbx_1__1__131_top_grid_pin_28_[0]),
		.top_grid_pin_29_(cbx_1__1__131_top_grid_pin_29_[0]),
		.top_grid_pin_30_(cbx_1__1__131_top_grid_pin_30_[0]),
		.top_grid_pin_31_(cbx_1__1__131_top_grid_pin_31_[0]),
		.ccff_tail(cbx_1__1__131_ccff_tail[0]));

	cbx_1__2_ cbx_1__12_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_0__12__0_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__12__0_chanx_left_out[0:19]),
		.ccff_head(sb_1__12__0_ccff_tail[0]),
		.chanx_left_out(cbx_1__12__0_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__12__0_chanx_right_out[0:19]),
		.top_grid_pin_0_(cbx_1__12__0_top_grid_pin_0_[0]),
		.ccff_tail(cbx_1__12__0_ccff_tail[0]));

	cbx_1__2_ cbx_2__12_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__12__0_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__12__1_chanx_left_out[0:19]),
		.ccff_head(sb_1__12__1_ccff_tail[0]),
		.chanx_left_out(cbx_1__12__1_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__12__1_chanx_right_out[0:19]),
		.top_grid_pin_0_(cbx_1__12__1_top_grid_pin_0_[0]),
		.ccff_tail(cbx_1__12__1_ccff_tail[0]));

	cbx_1__2_ cbx_3__12_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__12__1_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__12__2_chanx_left_out[0:19]),
		.ccff_head(sb_1__12__2_ccff_tail[0]),
		.chanx_left_out(cbx_1__12__2_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__12__2_chanx_right_out[0:19]),
		.top_grid_pin_0_(cbx_1__12__2_top_grid_pin_0_[0]),
		.ccff_tail(cbx_1__12__2_ccff_tail[0]));

	cbx_1__2_ cbx_4__12_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__12__2_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__12__3_chanx_left_out[0:19]),
		.ccff_head(sb_1__12__3_ccff_tail[0]),
		.chanx_left_out(cbx_1__12__3_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__12__3_chanx_right_out[0:19]),
		.top_grid_pin_0_(cbx_1__12__3_top_grid_pin_0_[0]),
		.ccff_tail(cbx_1__12__3_ccff_tail[0]));

	cbx_1__2_ cbx_5__12_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__12__3_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__12__4_chanx_left_out[0:19]),
		.ccff_head(sb_1__12__4_ccff_tail[0]),
		.chanx_left_out(cbx_1__12__4_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__12__4_chanx_right_out[0:19]),
		.top_grid_pin_0_(cbx_1__12__4_top_grid_pin_0_[0]),
		.ccff_tail(cbx_1__12__4_ccff_tail[0]));

	cbx_1__2_ cbx_6__12_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__12__4_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__12__5_chanx_left_out[0:19]),
		.ccff_head(sb_1__12__5_ccff_tail[0]),
		.chanx_left_out(cbx_1__12__5_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__12__5_chanx_right_out[0:19]),
		.top_grid_pin_0_(cbx_1__12__5_top_grid_pin_0_[0]),
		.ccff_tail(cbx_1__12__5_ccff_tail[0]));

	cbx_1__2_ cbx_7__12_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__12__5_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__12__6_chanx_left_out[0:19]),
		.ccff_head(sb_1__12__6_ccff_tail[0]),
		.chanx_left_out(cbx_1__12__6_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__12__6_chanx_right_out[0:19]),
		.top_grid_pin_0_(cbx_1__12__6_top_grid_pin_0_[0]),
		.ccff_tail(cbx_1__12__6_ccff_tail[0]));

	cbx_1__2_ cbx_8__12_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__12__6_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__12__7_chanx_left_out[0:19]),
		.ccff_head(sb_1__12__7_ccff_tail[0]),
		.chanx_left_out(cbx_1__12__7_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__12__7_chanx_right_out[0:19]),
		.top_grid_pin_0_(cbx_1__12__7_top_grid_pin_0_[0]),
		.ccff_tail(cbx_1__12__7_ccff_tail[0]));

	cbx_1__2_ cbx_9__12_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__12__7_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__12__8_chanx_left_out[0:19]),
		.ccff_head(sb_1__12__8_ccff_tail[0]),
		.chanx_left_out(cbx_1__12__8_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__12__8_chanx_right_out[0:19]),
		.top_grid_pin_0_(cbx_1__12__8_top_grid_pin_0_[0]),
		.ccff_tail(cbx_1__12__8_ccff_tail[0]));

	cbx_1__2_ cbx_10__12_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__12__8_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__12__9_chanx_left_out[0:19]),
		.ccff_head(sb_1__12__9_ccff_tail[0]),
		.chanx_left_out(cbx_1__12__9_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__12__9_chanx_right_out[0:19]),
		.top_grid_pin_0_(cbx_1__12__9_top_grid_pin_0_[0]),
		.ccff_tail(cbx_1__12__9_ccff_tail[0]));

	cbx_1__2_ cbx_11__12_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__12__9_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__12__10_chanx_left_out[0:19]),
		.ccff_head(sb_1__12__10_ccff_tail[0]),
		.chanx_left_out(cbx_1__12__10_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__12__10_chanx_right_out[0:19]),
		.top_grid_pin_0_(cbx_1__12__10_top_grid_pin_0_[0]),
		.ccff_tail(cbx_1__12__10_ccff_tail[0]));

	cbx_1__2_ cbx_12__12_ (
		.prog_clk(prog_clk[0]),
		.chanx_left_in(sb_1__12__10_chanx_right_out[0:19]),
		.chanx_right_in(sb_12__12__0_chanx_left_out[0:19]),
		.ccff_head(sb_12__12__0_ccff_tail[0]),
		.chanx_left_out(cbx_1__12__11_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__12__11_chanx_right_out[0:19]),
		.top_grid_pin_0_(cbx_1__12__11_top_grid_pin_0_[0]),
		.ccff_tail(cbx_1__12__11_ccff_tail[0]));

	cby_0__1_ cby_0__1_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_0__0__0_chany_top_out[0:19]),
		.chany_top_in(sb_0__1__0_chany_bottom_out[0:19]),
		.ccff_head(sb_0__1__0_ccff_tail[0]),
		.chany_bottom_out(cby_0__1__0_chany_bottom_out[0:19]),
		.chany_top_out(cby_0__1__0_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_0__1__0_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_0__1__0_left_grid_pin_0_[0]),
		.ccff_tail(cby_0__1__0_ccff_tail[0]));

	cby_0__1_ cby_0__2_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_0__1__0_chany_top_out[0:19]),
		.chany_top_in(sb_0__1__1_chany_bottom_out[0:19]),
		.ccff_head(sb_0__1__1_ccff_tail[0]),
		.chany_bottom_out(cby_0__1__1_chany_bottom_out[0:19]),
		.chany_top_out(cby_0__1__1_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_0__1__1_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_0__1__1_left_grid_pin_0_[0]),
		.ccff_tail(cby_0__1__1_ccff_tail[0]));

	cby_0__1_ cby_0__3_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_0__1__1_chany_top_out[0:19]),
		.chany_top_in(sb_0__1__2_chany_bottom_out[0:19]),
		.ccff_head(sb_0__1__2_ccff_tail[0]),
		.chany_bottom_out(cby_0__1__2_chany_bottom_out[0:19]),
		.chany_top_out(cby_0__1__2_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_0__1__2_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_0__1__2_left_grid_pin_0_[0]),
		.ccff_tail(cby_0__1__2_ccff_tail[0]));

	cby_0__1_ cby_0__4_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_0__1__2_chany_top_out[0:19]),
		.chany_top_in(sb_0__1__3_chany_bottom_out[0:19]),
		.ccff_head(sb_0__1__3_ccff_tail[0]),
		.chany_bottom_out(cby_0__1__3_chany_bottom_out[0:19]),
		.chany_top_out(cby_0__1__3_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_0__1__3_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_0__1__3_left_grid_pin_0_[0]),
		.ccff_tail(cby_0__1__3_ccff_tail[0]));

	cby_0__1_ cby_0__5_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_0__1__3_chany_top_out[0:19]),
		.chany_top_in(sb_0__1__4_chany_bottom_out[0:19]),
		.ccff_head(sb_0__1__4_ccff_tail[0]),
		.chany_bottom_out(cby_0__1__4_chany_bottom_out[0:19]),
		.chany_top_out(cby_0__1__4_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_0__1__4_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_0__1__4_left_grid_pin_0_[0]),
		.ccff_tail(cby_0__1__4_ccff_tail[0]));

	cby_0__1_ cby_0__6_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_0__1__4_chany_top_out[0:19]),
		.chany_top_in(sb_0__1__5_chany_bottom_out[0:19]),
		.ccff_head(sb_0__1__5_ccff_tail[0]),
		.chany_bottom_out(cby_0__1__5_chany_bottom_out[0:19]),
		.chany_top_out(cby_0__1__5_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_0__1__5_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_0__1__5_left_grid_pin_0_[0]),
		.ccff_tail(cby_0__1__5_ccff_tail[0]));

	cby_0__1_ cby_0__7_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_0__1__5_chany_top_out[0:19]),
		.chany_top_in(sb_0__1__6_chany_bottom_out[0:19]),
		.ccff_head(sb_0__1__6_ccff_tail[0]),
		.chany_bottom_out(cby_0__1__6_chany_bottom_out[0:19]),
		.chany_top_out(cby_0__1__6_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_0__1__6_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_0__1__6_left_grid_pin_0_[0]),
		.ccff_tail(cby_0__1__6_ccff_tail[0]));

	cby_0__1_ cby_0__8_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_0__1__6_chany_top_out[0:19]),
		.chany_top_in(sb_0__1__7_chany_bottom_out[0:19]),
		.ccff_head(sb_0__1__7_ccff_tail[0]),
		.chany_bottom_out(cby_0__1__7_chany_bottom_out[0:19]),
		.chany_top_out(cby_0__1__7_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_0__1__7_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_0__1__7_left_grid_pin_0_[0]),
		.ccff_tail(cby_0__1__7_ccff_tail[0]));

	cby_0__1_ cby_0__9_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_0__1__7_chany_top_out[0:19]),
		.chany_top_in(sb_0__1__8_chany_bottom_out[0:19]),
		.ccff_head(sb_0__1__8_ccff_tail[0]),
		.chany_bottom_out(cby_0__1__8_chany_bottom_out[0:19]),
		.chany_top_out(cby_0__1__8_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_0__1__8_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_0__1__8_left_grid_pin_0_[0]),
		.ccff_tail(cby_0__1__8_ccff_tail[0]));

	cby_0__1_ cby_0__10_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_0__1__8_chany_top_out[0:19]),
		.chany_top_in(sb_0__1__9_chany_bottom_out[0:19]),
		.ccff_head(sb_0__1__9_ccff_tail[0]),
		.chany_bottom_out(cby_0__1__9_chany_bottom_out[0:19]),
		.chany_top_out(cby_0__1__9_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_0__1__9_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_0__1__9_left_grid_pin_0_[0]),
		.ccff_tail(cby_0__1__9_ccff_tail[0]));

	cby_0__1_ cby_0__11_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_0__1__9_chany_top_out[0:19]),
		.chany_top_in(sb_0__1__10_chany_bottom_out[0:19]),
		.ccff_head(sb_0__1__10_ccff_tail[0]),
		.chany_bottom_out(cby_0__1__10_chany_bottom_out[0:19]),
		.chany_top_out(cby_0__1__10_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_0__1__10_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_0__1__10_left_grid_pin_0_[0]),
		.ccff_tail(cby_0__1__10_ccff_tail[0]));

	cby_0__1_ cby_0__12_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_0__1__10_chany_top_out[0:19]),
		.chany_top_in(sb_0__12__0_chany_bottom_out[0:19]),
		.ccff_head(sb_0__12__0_ccff_tail[0]),
		.chany_bottom_out(cby_0__1__11_chany_bottom_out[0:19]),
		.chany_top_out(cby_0__1__11_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_0__1__11_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_0__1__11_left_grid_pin_0_[0]),
		.ccff_tail(cby_0__1__11_ccff_tail[0]));

	cby_1__1_ cby_1__1_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__0__0_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__0_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_0_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__0_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__0_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__0_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__0_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__0_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__0_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__0_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__0_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__0_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__0_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__0_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__0_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__0_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__0_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__0_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__0_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__0_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__0_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__0_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__0_ccff_tail[0]));

	cby_1__1_ cby_1__2_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__0_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__1_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_1_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__1_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__1_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__1_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__1_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__1_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__1_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__1_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__1_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__1_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__1_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__1_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__1_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__1_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__1_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__1_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__1_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__1_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__1_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__1_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__1_ccff_tail[0]));

	cby_1__1_ cby_1__3_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__1_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__2_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_2_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__2_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__2_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__2_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__2_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__2_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__2_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__2_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__2_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__2_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__2_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__2_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__2_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__2_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__2_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__2_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__2_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__2_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__2_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__2_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__2_ccff_tail[0]));

	cby_1__1_ cby_1__4_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__2_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__3_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_3_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__3_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__3_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__3_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__3_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__3_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__3_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__3_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__3_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__3_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__3_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__3_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__3_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__3_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__3_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__3_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__3_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__3_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__3_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__3_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__3_ccff_tail[0]));

	cby_1__1_ cby_1__5_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__3_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__4_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_4_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__4_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__4_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__4_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__4_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__4_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__4_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__4_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__4_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__4_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__4_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__4_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__4_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__4_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__4_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__4_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__4_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__4_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__4_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__4_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__4_ccff_tail[0]));

	cby_1__1_ cby_1__6_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__4_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__5_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_5_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__5_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__5_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__5_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__5_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__5_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__5_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__5_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__5_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__5_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__5_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__5_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__5_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__5_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__5_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__5_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__5_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__5_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__5_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__5_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__5_ccff_tail[0]));

	cby_1__1_ cby_1__7_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__5_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__6_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_6_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__6_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__6_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__6_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__6_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__6_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__6_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__6_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__6_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__6_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__6_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__6_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__6_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__6_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__6_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__6_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__6_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__6_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__6_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__6_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__6_ccff_tail[0]));

	cby_1__1_ cby_1__8_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__6_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__7_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_7_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__7_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__7_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__7_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__7_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__7_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__7_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__7_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__7_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__7_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__7_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__7_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__7_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__7_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__7_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__7_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__7_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__7_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__7_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__7_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__7_ccff_tail[0]));

	cby_1__1_ cby_1__9_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__7_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__8_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_8_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__8_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__8_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__8_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__8_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__8_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__8_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__8_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__8_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__8_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__8_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__8_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__8_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__8_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__8_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__8_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__8_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__8_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__8_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__8_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__8_ccff_tail[0]));

	cby_1__1_ cby_1__10_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__8_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__9_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_9_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__9_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__9_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__9_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__9_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__9_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__9_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__9_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__9_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__9_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__9_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__9_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__9_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__9_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__9_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__9_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__9_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__9_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__9_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__9_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__9_ccff_tail[0]));

	cby_1__1_ cby_1__11_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__9_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__10_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_10_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__10_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__10_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__10_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__10_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__10_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__10_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__10_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__10_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__10_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__10_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__10_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__10_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__10_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__10_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__10_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__10_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__10_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__10_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__10_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__10_ccff_tail[0]));

	cby_1__1_ cby_1__12_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__10_chany_top_out[0:19]),
		.chany_top_in(sb_1__12__0_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_11_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__11_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__11_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__11_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__11_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__11_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__11_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__11_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__11_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__11_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__11_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__11_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__11_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__11_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__11_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__11_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__11_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__11_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__11_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__11_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__11_ccff_tail[0]));

	cby_1__1_ cby_2__1_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__0__1_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__11_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_12_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__12_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__12_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__12_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__12_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__12_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__12_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__12_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__12_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__12_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__12_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__12_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__12_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__12_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__12_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__12_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__12_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__12_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__12_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__12_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__12_ccff_tail[0]));

	cby_1__1_ cby_2__2_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__11_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__12_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_13_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__13_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__13_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__13_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__13_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__13_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__13_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__13_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__13_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__13_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__13_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__13_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__13_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__13_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__13_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__13_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__13_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__13_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__13_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__13_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__13_ccff_tail[0]));

	cby_1__1_ cby_2__3_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__12_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__13_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_14_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__14_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__14_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__14_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__14_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__14_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__14_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__14_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__14_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__14_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__14_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__14_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__14_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__14_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__14_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__14_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__14_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__14_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__14_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__14_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__14_ccff_tail[0]));

	cby_1__1_ cby_2__4_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__13_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__14_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_15_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__15_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__15_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__15_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__15_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__15_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__15_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__15_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__15_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__15_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__15_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__15_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__15_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__15_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__15_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__15_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__15_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__15_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__15_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__15_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__15_ccff_tail[0]));

	cby_1__1_ cby_2__5_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__14_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__15_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_16_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__16_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__16_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__16_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__16_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__16_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__16_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__16_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__16_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__16_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__16_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__16_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__16_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__16_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__16_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__16_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__16_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__16_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__16_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__16_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__16_ccff_tail[0]));

	cby_1__1_ cby_2__6_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__15_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__16_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_17_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__17_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__17_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__17_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__17_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__17_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__17_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__17_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__17_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__17_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__17_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__17_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__17_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__17_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__17_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__17_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__17_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__17_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__17_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__17_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__17_ccff_tail[0]));

	cby_1__1_ cby_2__7_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__16_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__17_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_18_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__18_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__18_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__18_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__18_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__18_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__18_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__18_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__18_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__18_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__18_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__18_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__18_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__18_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__18_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__18_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__18_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__18_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__18_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__18_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__18_ccff_tail[0]));

	cby_1__1_ cby_2__8_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__17_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__18_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_19_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__19_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__19_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__19_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__19_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__19_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__19_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__19_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__19_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__19_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__19_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__19_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__19_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__19_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__19_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__19_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__19_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__19_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__19_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__19_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__19_ccff_tail[0]));

	cby_1__1_ cby_2__9_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__18_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__19_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_20_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__20_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__20_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__20_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__20_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__20_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__20_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__20_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__20_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__20_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__20_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__20_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__20_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__20_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__20_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__20_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__20_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__20_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__20_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__20_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__20_ccff_tail[0]));

	cby_1__1_ cby_2__10_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__19_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__20_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_21_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__21_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__21_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__21_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__21_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__21_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__21_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__21_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__21_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__21_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__21_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__21_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__21_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__21_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__21_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__21_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__21_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__21_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__21_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__21_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__21_ccff_tail[0]));

	cby_1__1_ cby_2__11_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__20_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__21_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_22_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__22_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__22_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__22_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__22_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__22_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__22_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__22_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__22_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__22_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__22_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__22_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__22_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__22_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__22_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__22_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__22_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__22_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__22_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__22_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__22_ccff_tail[0]));

	cby_1__1_ cby_2__12_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__21_chany_top_out[0:19]),
		.chany_top_in(sb_1__12__1_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_23_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__23_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__23_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__23_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__23_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__23_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__23_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__23_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__23_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__23_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__23_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__23_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__23_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__23_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__23_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__23_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__23_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__23_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__23_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__23_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__23_ccff_tail[0]));

	cby_1__1_ cby_3__1_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__0__2_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__22_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_24_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__24_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__24_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__24_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__24_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__24_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__24_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__24_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__24_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__24_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__24_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__24_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__24_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__24_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__24_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__24_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__24_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__24_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__24_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__24_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__24_ccff_tail[0]));

	cby_1__1_ cby_3__2_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__22_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__23_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_25_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__25_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__25_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__25_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__25_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__25_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__25_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__25_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__25_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__25_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__25_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__25_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__25_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__25_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__25_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__25_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__25_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__25_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__25_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__25_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__25_ccff_tail[0]));

	cby_1__1_ cby_3__3_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__23_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__24_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_26_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__26_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__26_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__26_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__26_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__26_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__26_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__26_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__26_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__26_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__26_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__26_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__26_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__26_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__26_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__26_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__26_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__26_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__26_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__26_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__26_ccff_tail[0]));

	cby_1__1_ cby_3__4_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__24_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__25_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_27_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__27_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__27_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__27_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__27_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__27_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__27_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__27_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__27_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__27_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__27_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__27_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__27_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__27_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__27_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__27_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__27_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__27_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__27_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__27_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__27_ccff_tail[0]));

	cby_1__1_ cby_3__5_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__25_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__26_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_28_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__28_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__28_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__28_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__28_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__28_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__28_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__28_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__28_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__28_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__28_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__28_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__28_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__28_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__28_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__28_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__28_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__28_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__28_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__28_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__28_ccff_tail[0]));

	cby_1__1_ cby_3__6_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__26_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__27_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_29_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__29_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__29_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__29_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__29_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__29_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__29_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__29_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__29_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__29_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__29_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__29_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__29_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__29_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__29_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__29_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__29_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__29_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__29_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__29_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__29_ccff_tail[0]));

	cby_1__1_ cby_3__7_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__27_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__28_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_30_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__30_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__30_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__30_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__30_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__30_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__30_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__30_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__30_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__30_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__30_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__30_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__30_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__30_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__30_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__30_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__30_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__30_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__30_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__30_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__30_ccff_tail[0]));

	cby_1__1_ cby_3__8_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__28_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__29_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_31_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__31_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__31_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__31_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__31_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__31_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__31_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__31_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__31_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__31_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__31_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__31_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__31_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__31_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__31_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__31_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__31_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__31_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__31_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__31_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__31_ccff_tail[0]));

	cby_1__1_ cby_3__9_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__29_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__30_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_32_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__32_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__32_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__32_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__32_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__32_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__32_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__32_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__32_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__32_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__32_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__32_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__32_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__32_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__32_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__32_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__32_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__32_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__32_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__32_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__32_ccff_tail[0]));

	cby_1__1_ cby_3__10_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__30_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__31_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_33_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__33_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__33_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__33_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__33_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__33_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__33_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__33_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__33_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__33_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__33_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__33_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__33_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__33_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__33_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__33_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__33_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__33_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__33_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__33_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__33_ccff_tail[0]));

	cby_1__1_ cby_3__11_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__31_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__32_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_34_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__34_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__34_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__34_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__34_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__34_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__34_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__34_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__34_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__34_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__34_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__34_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__34_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__34_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__34_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__34_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__34_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__34_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__34_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__34_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__34_ccff_tail[0]));

	cby_1__1_ cby_3__12_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__32_chany_top_out[0:19]),
		.chany_top_in(sb_1__12__2_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_35_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__35_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__35_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__35_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__35_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__35_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__35_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__35_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__35_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__35_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__35_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__35_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__35_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__35_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__35_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__35_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__35_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__35_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__35_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__35_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__35_ccff_tail[0]));

	cby_1__1_ cby_4__1_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__0__3_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__33_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_36_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__36_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__36_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__36_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__36_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__36_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__36_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__36_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__36_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__36_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__36_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__36_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__36_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__36_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__36_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__36_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__36_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__36_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__36_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__36_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__36_ccff_tail[0]));

	cby_1__1_ cby_4__2_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__33_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__34_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_37_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__37_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__37_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__37_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__37_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__37_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__37_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__37_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__37_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__37_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__37_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__37_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__37_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__37_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__37_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__37_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__37_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__37_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__37_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__37_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__37_ccff_tail[0]));

	cby_1__1_ cby_4__3_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__34_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__35_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_38_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__38_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__38_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__38_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__38_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__38_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__38_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__38_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__38_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__38_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__38_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__38_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__38_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__38_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__38_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__38_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__38_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__38_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__38_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__38_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__38_ccff_tail[0]));

	cby_1__1_ cby_4__4_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__35_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__36_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_39_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__39_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__39_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__39_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__39_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__39_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__39_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__39_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__39_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__39_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__39_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__39_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__39_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__39_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__39_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__39_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__39_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__39_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__39_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__39_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__39_ccff_tail[0]));

	cby_1__1_ cby_4__5_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__36_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__37_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_40_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__40_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__40_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__40_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__40_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__40_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__40_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__40_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__40_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__40_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__40_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__40_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__40_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__40_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__40_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__40_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__40_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__40_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__40_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__40_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__40_ccff_tail[0]));

	cby_1__1_ cby_4__6_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__37_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__38_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_41_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__41_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__41_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__41_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__41_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__41_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__41_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__41_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__41_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__41_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__41_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__41_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__41_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__41_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__41_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__41_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__41_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__41_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__41_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__41_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__41_ccff_tail[0]));

	cby_1__1_ cby_4__7_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__38_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__39_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_42_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__42_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__42_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__42_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__42_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__42_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__42_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__42_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__42_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__42_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__42_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__42_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__42_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__42_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__42_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__42_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__42_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__42_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__42_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__42_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__42_ccff_tail[0]));

	cby_1__1_ cby_4__8_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__39_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__40_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_43_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__43_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__43_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__43_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__43_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__43_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__43_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__43_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__43_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__43_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__43_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__43_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__43_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__43_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__43_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__43_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__43_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__43_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__43_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__43_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__43_ccff_tail[0]));

	cby_1__1_ cby_4__9_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__40_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__41_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_44_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__44_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__44_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__44_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__44_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__44_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__44_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__44_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__44_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__44_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__44_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__44_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__44_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__44_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__44_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__44_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__44_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__44_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__44_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__44_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__44_ccff_tail[0]));

	cby_1__1_ cby_4__10_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__41_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__42_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_45_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__45_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__45_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__45_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__45_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__45_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__45_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__45_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__45_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__45_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__45_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__45_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__45_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__45_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__45_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__45_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__45_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__45_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__45_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__45_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__45_ccff_tail[0]));

	cby_1__1_ cby_4__11_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__42_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__43_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_46_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__46_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__46_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__46_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__46_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__46_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__46_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__46_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__46_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__46_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__46_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__46_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__46_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__46_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__46_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__46_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__46_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__46_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__46_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__46_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__46_ccff_tail[0]));

	cby_1__1_ cby_4__12_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__43_chany_top_out[0:19]),
		.chany_top_in(sb_1__12__3_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_47_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__47_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__47_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__47_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__47_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__47_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__47_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__47_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__47_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__47_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__47_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__47_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__47_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__47_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__47_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__47_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__47_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__47_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__47_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__47_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__47_ccff_tail[0]));

	cby_1__1_ cby_5__1_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__0__4_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__44_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_48_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__48_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__48_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__48_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__48_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__48_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__48_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__48_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__48_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__48_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__48_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__48_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__48_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__48_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__48_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__48_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__48_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__48_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__48_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__48_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__48_ccff_tail[0]));

	cby_1__1_ cby_5__2_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__44_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__45_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_49_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__49_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__49_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__49_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__49_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__49_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__49_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__49_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__49_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__49_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__49_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__49_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__49_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__49_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__49_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__49_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__49_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__49_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__49_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__49_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__49_ccff_tail[0]));

	cby_1__1_ cby_5__3_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__45_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__46_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_50_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__50_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__50_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__50_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__50_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__50_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__50_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__50_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__50_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__50_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__50_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__50_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__50_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__50_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__50_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__50_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__50_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__50_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__50_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__50_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__50_ccff_tail[0]));

	cby_1__1_ cby_5__4_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__46_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__47_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_51_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__51_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__51_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__51_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__51_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__51_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__51_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__51_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__51_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__51_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__51_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__51_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__51_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__51_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__51_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__51_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__51_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__51_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__51_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__51_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__51_ccff_tail[0]));

	cby_1__1_ cby_5__5_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__47_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__48_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_52_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__52_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__52_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__52_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__52_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__52_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__52_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__52_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__52_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__52_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__52_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__52_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__52_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__52_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__52_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__52_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__52_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__52_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__52_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__52_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__52_ccff_tail[0]));

	cby_1__1_ cby_5__6_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__48_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__49_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_53_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__53_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__53_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__53_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__53_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__53_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__53_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__53_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__53_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__53_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__53_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__53_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__53_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__53_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__53_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__53_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__53_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__53_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__53_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__53_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__53_ccff_tail[0]));

	cby_1__1_ cby_5__7_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__49_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__50_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_54_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__54_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__54_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__54_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__54_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__54_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__54_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__54_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__54_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__54_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__54_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__54_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__54_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__54_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__54_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__54_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__54_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__54_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__54_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__54_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__54_ccff_tail[0]));

	cby_1__1_ cby_5__8_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__50_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__51_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_55_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__55_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__55_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__55_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__55_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__55_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__55_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__55_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__55_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__55_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__55_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__55_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__55_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__55_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__55_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__55_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__55_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__55_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__55_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__55_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__55_ccff_tail[0]));

	cby_1__1_ cby_5__9_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__51_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__52_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_56_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__56_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__56_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__56_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__56_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__56_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__56_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__56_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__56_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__56_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__56_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__56_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__56_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__56_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__56_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__56_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__56_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__56_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__56_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__56_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__56_ccff_tail[0]));

	cby_1__1_ cby_5__10_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__52_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__53_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_57_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__57_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__57_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__57_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__57_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__57_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__57_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__57_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__57_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__57_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__57_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__57_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__57_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__57_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__57_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__57_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__57_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__57_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__57_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__57_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__57_ccff_tail[0]));

	cby_1__1_ cby_5__11_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__53_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__54_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_58_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__58_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__58_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__58_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__58_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__58_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__58_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__58_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__58_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__58_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__58_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__58_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__58_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__58_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__58_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__58_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__58_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__58_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__58_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__58_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__58_ccff_tail[0]));

	cby_1__1_ cby_5__12_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__54_chany_top_out[0:19]),
		.chany_top_in(sb_1__12__4_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_59_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__59_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__59_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__59_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__59_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__59_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__59_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__59_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__59_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__59_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__59_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__59_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__59_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__59_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__59_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__59_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__59_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__59_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__59_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__59_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__59_ccff_tail[0]));

	cby_1__1_ cby_6__1_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__0__5_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__55_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_60_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__60_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__60_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__60_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__60_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__60_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__60_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__60_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__60_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__60_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__60_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__60_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__60_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__60_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__60_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__60_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__60_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__60_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__60_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__60_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__60_ccff_tail[0]));

	cby_1__1_ cby_6__2_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__55_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__56_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_61_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__61_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__61_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__61_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__61_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__61_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__61_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__61_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__61_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__61_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__61_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__61_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__61_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__61_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__61_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__61_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__61_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__61_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__61_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__61_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__61_ccff_tail[0]));

	cby_1__1_ cby_6__3_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__56_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__57_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_62_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__62_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__62_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__62_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__62_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__62_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__62_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__62_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__62_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__62_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__62_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__62_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__62_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__62_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__62_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__62_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__62_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__62_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__62_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__62_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__62_ccff_tail[0]));

	cby_1__1_ cby_6__4_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__57_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__58_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_63_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__63_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__63_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__63_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__63_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__63_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__63_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__63_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__63_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__63_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__63_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__63_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__63_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__63_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__63_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__63_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__63_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__63_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__63_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__63_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__63_ccff_tail[0]));

	cby_1__1_ cby_6__5_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__58_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__59_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_64_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__64_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__64_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__64_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__64_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__64_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__64_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__64_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__64_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__64_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__64_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__64_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__64_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__64_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__64_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__64_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__64_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__64_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__64_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__64_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__64_ccff_tail[0]));

	cby_1__1_ cby_6__6_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__59_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__60_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_65_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__65_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__65_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__65_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__65_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__65_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__65_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__65_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__65_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__65_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__65_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__65_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__65_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__65_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__65_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__65_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__65_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__65_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__65_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__65_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__65_ccff_tail[0]));

	cby_1__1_ cby_6__7_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__60_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__61_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_66_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__66_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__66_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__66_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__66_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__66_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__66_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__66_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__66_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__66_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__66_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__66_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__66_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__66_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__66_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__66_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__66_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__66_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__66_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__66_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__66_ccff_tail[0]));

	cby_1__1_ cby_6__8_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__61_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__62_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_67_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__67_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__67_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__67_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__67_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__67_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__67_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__67_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__67_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__67_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__67_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__67_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__67_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__67_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__67_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__67_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__67_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__67_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__67_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__67_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__67_ccff_tail[0]));

	cby_1__1_ cby_6__9_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__62_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__63_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_68_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__68_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__68_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__68_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__68_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__68_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__68_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__68_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__68_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__68_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__68_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__68_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__68_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__68_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__68_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__68_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__68_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__68_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__68_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__68_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__68_ccff_tail[0]));

	cby_1__1_ cby_6__10_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__63_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__64_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_69_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__69_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__69_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__69_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__69_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__69_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__69_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__69_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__69_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__69_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__69_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__69_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__69_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__69_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__69_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__69_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__69_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__69_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__69_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__69_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__69_ccff_tail[0]));

	cby_1__1_ cby_6__11_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__64_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__65_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_70_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__70_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__70_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__70_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__70_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__70_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__70_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__70_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__70_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__70_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__70_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__70_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__70_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__70_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__70_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__70_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__70_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__70_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__70_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__70_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__70_ccff_tail[0]));

	cby_1__1_ cby_6__12_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__65_chany_top_out[0:19]),
		.chany_top_in(sb_1__12__5_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_71_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__71_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__71_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__71_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__71_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__71_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__71_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__71_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__71_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__71_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__71_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__71_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__71_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__71_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__71_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__71_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__71_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__71_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__71_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__71_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__71_ccff_tail[0]));

	cby_1__1_ cby_7__1_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__0__6_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__66_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_72_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__72_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__72_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__72_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__72_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__72_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__72_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__72_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__72_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__72_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__72_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__72_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__72_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__72_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__72_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__72_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__72_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__72_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__72_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__72_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__72_ccff_tail[0]));

	cby_1__1_ cby_7__2_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__66_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__67_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_73_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__73_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__73_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__73_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__73_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__73_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__73_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__73_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__73_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__73_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__73_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__73_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__73_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__73_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__73_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__73_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__73_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__73_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__73_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__73_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__73_ccff_tail[0]));

	cby_1__1_ cby_7__3_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__67_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__68_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_74_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__74_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__74_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__74_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__74_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__74_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__74_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__74_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__74_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__74_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__74_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__74_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__74_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__74_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__74_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__74_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__74_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__74_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__74_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__74_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__74_ccff_tail[0]));

	cby_1__1_ cby_7__4_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__68_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__69_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_75_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__75_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__75_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__75_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__75_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__75_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__75_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__75_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__75_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__75_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__75_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__75_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__75_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__75_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__75_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__75_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__75_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__75_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__75_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__75_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__75_ccff_tail[0]));

	cby_1__1_ cby_7__5_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__69_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__70_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_76_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__76_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__76_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__76_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__76_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__76_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__76_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__76_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__76_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__76_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__76_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__76_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__76_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__76_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__76_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__76_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__76_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__76_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__76_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__76_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__76_ccff_tail[0]));

	cby_1__1_ cby_7__6_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__70_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__71_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_77_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__77_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__77_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__77_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__77_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__77_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__77_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__77_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__77_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__77_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__77_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__77_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__77_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__77_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__77_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__77_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__77_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__77_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__77_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__77_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__77_ccff_tail[0]));

	cby_1__1_ cby_7__7_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__71_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__72_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_78_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__78_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__78_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__78_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__78_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__78_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__78_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__78_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__78_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__78_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__78_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__78_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__78_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__78_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__78_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__78_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__78_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__78_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__78_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__78_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__78_ccff_tail[0]));

	cby_1__1_ cby_7__8_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__72_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__73_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_79_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__79_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__79_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__79_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__79_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__79_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__79_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__79_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__79_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__79_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__79_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__79_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__79_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__79_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__79_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__79_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__79_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__79_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__79_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__79_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__79_ccff_tail[0]));

	cby_1__1_ cby_7__9_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__73_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__74_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_80_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__80_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__80_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__80_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__80_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__80_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__80_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__80_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__80_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__80_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__80_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__80_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__80_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__80_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__80_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__80_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__80_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__80_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__80_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__80_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__80_ccff_tail[0]));

	cby_1__1_ cby_7__10_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__74_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__75_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_81_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__81_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__81_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__81_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__81_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__81_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__81_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__81_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__81_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__81_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__81_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__81_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__81_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__81_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__81_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__81_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__81_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__81_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__81_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__81_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__81_ccff_tail[0]));

	cby_1__1_ cby_7__11_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__75_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__76_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_82_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__82_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__82_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__82_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__82_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__82_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__82_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__82_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__82_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__82_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__82_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__82_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__82_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__82_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__82_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__82_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__82_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__82_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__82_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__82_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__82_ccff_tail[0]));

	cby_1__1_ cby_7__12_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__76_chany_top_out[0:19]),
		.chany_top_in(sb_1__12__6_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_83_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__83_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__83_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__83_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__83_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__83_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__83_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__83_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__83_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__83_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__83_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__83_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__83_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__83_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__83_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__83_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__83_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__83_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__83_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__83_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__83_ccff_tail[0]));

	cby_1__1_ cby_8__1_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__0__7_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__77_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_84_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__84_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__84_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__84_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__84_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__84_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__84_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__84_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__84_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__84_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__84_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__84_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__84_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__84_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__84_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__84_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__84_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__84_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__84_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__84_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__84_ccff_tail[0]));

	cby_1__1_ cby_8__2_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__77_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__78_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_85_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__85_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__85_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__85_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__85_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__85_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__85_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__85_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__85_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__85_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__85_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__85_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__85_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__85_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__85_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__85_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__85_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__85_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__85_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__85_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__85_ccff_tail[0]));

	cby_1__1_ cby_8__3_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__78_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__79_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_86_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__86_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__86_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__86_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__86_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__86_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__86_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__86_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__86_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__86_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__86_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__86_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__86_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__86_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__86_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__86_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__86_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__86_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__86_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__86_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__86_ccff_tail[0]));

	cby_1__1_ cby_8__4_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__79_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__80_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_87_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__87_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__87_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__87_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__87_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__87_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__87_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__87_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__87_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__87_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__87_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__87_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__87_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__87_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__87_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__87_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__87_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__87_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__87_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__87_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__87_ccff_tail[0]));

	cby_1__1_ cby_8__5_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__80_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__81_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_88_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__88_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__88_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__88_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__88_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__88_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__88_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__88_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__88_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__88_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__88_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__88_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__88_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__88_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__88_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__88_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__88_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__88_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__88_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__88_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__88_ccff_tail[0]));

	cby_1__1_ cby_8__6_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__81_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__82_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_89_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__89_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__89_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__89_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__89_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__89_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__89_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__89_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__89_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__89_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__89_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__89_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__89_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__89_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__89_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__89_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__89_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__89_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__89_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__89_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__89_ccff_tail[0]));

	cby_1__1_ cby_8__7_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__82_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__83_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_90_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__90_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__90_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__90_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__90_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__90_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__90_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__90_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__90_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__90_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__90_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__90_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__90_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__90_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__90_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__90_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__90_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__90_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__90_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__90_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__90_ccff_tail[0]));

	cby_1__1_ cby_8__8_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__83_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__84_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_91_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__91_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__91_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__91_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__91_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__91_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__91_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__91_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__91_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__91_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__91_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__91_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__91_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__91_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__91_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__91_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__91_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__91_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__91_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__91_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__91_ccff_tail[0]));

	cby_1__1_ cby_8__9_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__84_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__85_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_92_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__92_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__92_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__92_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__92_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__92_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__92_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__92_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__92_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__92_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__92_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__92_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__92_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__92_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__92_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__92_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__92_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__92_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__92_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__92_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__92_ccff_tail[0]));

	cby_1__1_ cby_8__10_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__85_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__86_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_93_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__93_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__93_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__93_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__93_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__93_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__93_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__93_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__93_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__93_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__93_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__93_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__93_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__93_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__93_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__93_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__93_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__93_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__93_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__93_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__93_ccff_tail[0]));

	cby_1__1_ cby_8__11_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__86_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__87_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_94_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__94_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__94_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__94_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__94_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__94_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__94_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__94_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__94_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__94_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__94_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__94_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__94_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__94_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__94_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__94_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__94_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__94_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__94_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__94_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__94_ccff_tail[0]));

	cby_1__1_ cby_8__12_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__87_chany_top_out[0:19]),
		.chany_top_in(sb_1__12__7_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_95_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__95_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__95_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__95_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__95_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__95_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__95_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__95_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__95_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__95_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__95_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__95_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__95_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__95_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__95_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__95_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__95_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__95_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__95_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__95_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__95_ccff_tail[0]));

	cby_1__1_ cby_9__1_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__0__8_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__88_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_96_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__96_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__96_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__96_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__96_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__96_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__96_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__96_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__96_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__96_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__96_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__96_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__96_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__96_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__96_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__96_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__96_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__96_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__96_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__96_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__96_ccff_tail[0]));

	cby_1__1_ cby_9__2_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__88_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__89_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_97_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__97_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__97_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__97_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__97_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__97_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__97_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__97_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__97_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__97_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__97_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__97_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__97_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__97_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__97_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__97_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__97_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__97_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__97_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__97_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__97_ccff_tail[0]));

	cby_1__1_ cby_9__3_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__89_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__90_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_98_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__98_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__98_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__98_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__98_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__98_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__98_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__98_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__98_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__98_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__98_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__98_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__98_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__98_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__98_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__98_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__98_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__98_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__98_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__98_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__98_ccff_tail[0]));

	cby_1__1_ cby_9__4_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__90_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__91_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_99_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__99_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__99_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__99_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__99_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__99_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__99_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__99_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__99_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__99_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__99_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__99_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__99_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__99_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__99_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__99_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__99_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__99_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__99_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__99_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__99_ccff_tail[0]));

	cby_1__1_ cby_9__5_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__91_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__92_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_100_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__100_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__100_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__100_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__100_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__100_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__100_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__100_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__100_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__100_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__100_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__100_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__100_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__100_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__100_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__100_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__100_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__100_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__100_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__100_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__100_ccff_tail[0]));

	cby_1__1_ cby_9__6_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__92_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__93_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_101_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__101_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__101_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__101_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__101_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__101_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__101_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__101_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__101_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__101_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__101_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__101_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__101_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__101_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__101_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__101_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__101_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__101_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__101_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__101_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__101_ccff_tail[0]));

	cby_1__1_ cby_9__7_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__93_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__94_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_102_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__102_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__102_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__102_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__102_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__102_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__102_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__102_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__102_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__102_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__102_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__102_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__102_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__102_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__102_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__102_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__102_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__102_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__102_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__102_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__102_ccff_tail[0]));

	cby_1__1_ cby_9__8_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__94_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__95_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_103_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__103_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__103_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__103_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__103_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__103_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__103_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__103_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__103_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__103_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__103_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__103_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__103_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__103_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__103_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__103_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__103_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__103_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__103_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__103_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__103_ccff_tail[0]));

	cby_1__1_ cby_9__9_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__95_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__96_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_104_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__104_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__104_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__104_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__104_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__104_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__104_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__104_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__104_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__104_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__104_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__104_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__104_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__104_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__104_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__104_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__104_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__104_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__104_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__104_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__104_ccff_tail[0]));

	cby_1__1_ cby_9__10_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__96_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__97_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_105_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__105_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__105_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__105_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__105_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__105_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__105_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__105_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__105_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__105_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__105_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__105_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__105_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__105_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__105_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__105_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__105_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__105_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__105_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__105_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__105_ccff_tail[0]));

	cby_1__1_ cby_9__11_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__97_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__98_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_106_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__106_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__106_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__106_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__106_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__106_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__106_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__106_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__106_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__106_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__106_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__106_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__106_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__106_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__106_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__106_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__106_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__106_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__106_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__106_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__106_ccff_tail[0]));

	cby_1__1_ cby_9__12_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__98_chany_top_out[0:19]),
		.chany_top_in(sb_1__12__8_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_107_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__107_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__107_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__107_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__107_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__107_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__107_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__107_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__107_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__107_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__107_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__107_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__107_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__107_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__107_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__107_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__107_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__107_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__107_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__107_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__107_ccff_tail[0]));

	cby_1__1_ cby_10__1_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__0__9_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__99_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_108_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__108_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__108_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__108_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__108_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__108_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__108_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__108_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__108_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__108_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__108_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__108_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__108_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__108_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__108_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__108_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__108_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__108_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__108_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__108_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__108_ccff_tail[0]));

	cby_1__1_ cby_10__2_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__99_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__100_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_109_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__109_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__109_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__109_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__109_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__109_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__109_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__109_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__109_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__109_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__109_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__109_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__109_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__109_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__109_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__109_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__109_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__109_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__109_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__109_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__109_ccff_tail[0]));

	cby_1__1_ cby_10__3_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__100_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__101_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_110_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__110_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__110_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__110_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__110_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__110_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__110_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__110_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__110_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__110_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__110_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__110_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__110_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__110_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__110_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__110_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__110_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__110_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__110_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__110_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__110_ccff_tail[0]));

	cby_1__1_ cby_10__4_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__101_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__102_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_111_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__111_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__111_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__111_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__111_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__111_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__111_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__111_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__111_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__111_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__111_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__111_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__111_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__111_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__111_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__111_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__111_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__111_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__111_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__111_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__111_ccff_tail[0]));

	cby_1__1_ cby_10__5_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__102_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__103_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_112_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__112_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__112_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__112_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__112_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__112_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__112_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__112_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__112_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__112_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__112_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__112_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__112_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__112_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__112_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__112_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__112_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__112_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__112_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__112_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__112_ccff_tail[0]));

	cby_1__1_ cby_10__6_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__103_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__104_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_113_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__113_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__113_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__113_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__113_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__113_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__113_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__113_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__113_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__113_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__113_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__113_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__113_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__113_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__113_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__113_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__113_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__113_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__113_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__113_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__113_ccff_tail[0]));

	cby_1__1_ cby_10__7_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__104_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__105_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_114_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__114_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__114_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__114_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__114_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__114_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__114_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__114_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__114_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__114_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__114_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__114_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__114_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__114_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__114_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__114_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__114_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__114_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__114_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__114_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__114_ccff_tail[0]));

	cby_1__1_ cby_10__8_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__105_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__106_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_115_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__115_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__115_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__115_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__115_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__115_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__115_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__115_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__115_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__115_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__115_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__115_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__115_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__115_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__115_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__115_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__115_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__115_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__115_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__115_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__115_ccff_tail[0]));

	cby_1__1_ cby_10__9_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__106_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__107_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_116_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__116_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__116_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__116_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__116_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__116_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__116_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__116_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__116_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__116_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__116_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__116_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__116_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__116_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__116_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__116_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__116_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__116_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__116_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__116_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__116_ccff_tail[0]));

	cby_1__1_ cby_10__10_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__107_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__108_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_117_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__117_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__117_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__117_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__117_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__117_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__117_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__117_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__117_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__117_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__117_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__117_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__117_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__117_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__117_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__117_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__117_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__117_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__117_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__117_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__117_ccff_tail[0]));

	cby_1__1_ cby_10__11_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__108_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__109_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_118_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__118_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__118_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__118_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__118_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__118_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__118_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__118_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__118_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__118_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__118_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__118_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__118_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__118_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__118_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__118_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__118_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__118_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__118_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__118_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__118_ccff_tail[0]));

	cby_1__1_ cby_10__12_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__109_chany_top_out[0:19]),
		.chany_top_in(sb_1__12__9_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_119_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__119_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__119_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__119_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__119_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__119_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__119_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__119_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__119_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__119_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__119_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__119_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__119_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__119_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__119_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__119_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__119_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__119_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__119_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__119_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__119_ccff_tail[0]));

	cby_1__1_ cby_11__1_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__0__10_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__110_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_120_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__120_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__120_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__120_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__120_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__120_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__120_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__120_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__120_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__120_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__120_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__120_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__120_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__120_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__120_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__120_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__120_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__120_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__120_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__120_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__120_ccff_tail[0]));

	cby_1__1_ cby_11__2_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__110_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__111_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_121_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__121_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__121_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__121_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__121_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__121_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__121_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__121_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__121_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__121_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__121_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__121_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__121_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__121_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__121_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__121_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__121_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__121_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__121_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__121_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__121_ccff_tail[0]));

	cby_1__1_ cby_11__3_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__111_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__112_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_122_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__122_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__122_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__122_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__122_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__122_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__122_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__122_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__122_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__122_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__122_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__122_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__122_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__122_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__122_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__122_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__122_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__122_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__122_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__122_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__122_ccff_tail[0]));

	cby_1__1_ cby_11__4_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__112_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__113_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_123_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__123_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__123_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__123_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__123_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__123_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__123_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__123_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__123_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__123_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__123_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__123_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__123_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__123_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__123_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__123_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__123_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__123_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__123_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__123_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__123_ccff_tail[0]));

	cby_1__1_ cby_11__5_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__113_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__114_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_124_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__124_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__124_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__124_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__124_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__124_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__124_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__124_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__124_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__124_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__124_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__124_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__124_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__124_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__124_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__124_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__124_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__124_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__124_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__124_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__124_ccff_tail[0]));

	cby_1__1_ cby_11__6_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__114_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__115_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_125_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__125_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__125_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__125_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__125_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__125_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__125_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__125_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__125_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__125_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__125_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__125_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__125_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__125_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__125_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__125_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__125_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__125_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__125_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__125_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__125_ccff_tail[0]));

	cby_1__1_ cby_11__7_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__115_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__116_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_126_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__126_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__126_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__126_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__126_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__126_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__126_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__126_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__126_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__126_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__126_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__126_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__126_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__126_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__126_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__126_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__126_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__126_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__126_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__126_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__126_ccff_tail[0]));

	cby_1__1_ cby_11__8_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__116_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__117_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_127_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__127_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__127_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__127_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__127_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__127_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__127_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__127_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__127_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__127_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__127_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__127_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__127_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__127_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__127_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__127_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__127_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__127_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__127_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__127_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__127_ccff_tail[0]));

	cby_1__1_ cby_11__9_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__117_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__118_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_128_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__128_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__128_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__128_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__128_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__128_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__128_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__128_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__128_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__128_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__128_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__128_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__128_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__128_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__128_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__128_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__128_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__128_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__128_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__128_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__128_ccff_tail[0]));

	cby_1__1_ cby_11__10_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__118_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__119_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_129_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__129_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__129_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__129_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__129_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__129_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__129_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__129_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__129_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__129_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__129_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__129_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__129_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__129_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__129_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__129_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__129_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__129_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__129_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__129_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__129_ccff_tail[0]));

	cby_1__1_ cby_11__11_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__119_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__120_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_130_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__130_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__130_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__130_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__130_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__130_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__130_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__130_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__130_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__130_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__130_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__130_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__130_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__130_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__130_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__130_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__130_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__130_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__130_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__130_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__130_ccff_tail[0]));

	cby_1__1_ cby_11__12_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_1__1__120_chany_top_out[0:19]),
		.chany_top_in(sb_1__12__10_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_131_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__131_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__131_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__131_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__131_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__131_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__131_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__131_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__131_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__131_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__131_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__131_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__131_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__131_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__131_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__131_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__131_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__131_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__131_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__131_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__131_ccff_tail[0]));

	cby_1__1_ cby_12__1_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_12__0__0_chany_top_out[0:19]),
		.chany_top_in(sb_12__1__0_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_132_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__132_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__132_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__132_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__132_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__132_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__132_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__132_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__132_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__132_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__132_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__132_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__132_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__132_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__132_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__132_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__132_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__132_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__132_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__132_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__132_ccff_tail[0]));

	cby_1__1_ cby_12__2_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_12__1__0_chany_top_out[0:19]),
		.chany_top_in(sb_12__1__1_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_133_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__133_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__133_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__133_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__133_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__133_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__133_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__133_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__133_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__133_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__133_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__133_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__133_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__133_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__133_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__133_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__133_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__133_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__133_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__133_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__133_ccff_tail[0]));

	cby_1__1_ cby_12__3_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_12__1__1_chany_top_out[0:19]),
		.chany_top_in(sb_12__1__2_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_134_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__134_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__134_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__134_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__134_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__134_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__134_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__134_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__134_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__134_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__134_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__134_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__134_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__134_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__134_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__134_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__134_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__134_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__134_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__134_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__134_ccff_tail[0]));

	cby_1__1_ cby_12__4_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_12__1__2_chany_top_out[0:19]),
		.chany_top_in(sb_12__1__3_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_135_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__135_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__135_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__135_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__135_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__135_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__135_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__135_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__135_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__135_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__135_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__135_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__135_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__135_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__135_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__135_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__135_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__135_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__135_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__135_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__135_ccff_tail[0]));

	cby_1__1_ cby_12__5_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_12__1__3_chany_top_out[0:19]),
		.chany_top_in(sb_12__1__4_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_136_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__136_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__136_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__136_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__136_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__136_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__136_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__136_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__136_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__136_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__136_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__136_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__136_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__136_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__136_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__136_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__136_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__136_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__136_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__136_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__136_ccff_tail[0]));

	cby_1__1_ cby_12__6_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_12__1__4_chany_top_out[0:19]),
		.chany_top_in(sb_12__1__5_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_137_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__137_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__137_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__137_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__137_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__137_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__137_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__137_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__137_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__137_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__137_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__137_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__137_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__137_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__137_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__137_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__137_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__137_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__137_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__137_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__137_ccff_tail[0]));

	cby_1__1_ cby_12__7_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_12__1__5_chany_top_out[0:19]),
		.chany_top_in(sb_12__1__6_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_138_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__138_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__138_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__138_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__138_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__138_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__138_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__138_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__138_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__138_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__138_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__138_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__138_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__138_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__138_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__138_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__138_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__138_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__138_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__138_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__138_ccff_tail[0]));

	cby_1__1_ cby_12__8_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_12__1__6_chany_top_out[0:19]),
		.chany_top_in(sb_12__1__7_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_139_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__139_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__139_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__139_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__139_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__139_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__139_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__139_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__139_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__139_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__139_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__139_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__139_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__139_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__139_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__139_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__139_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__139_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__139_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__139_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__139_ccff_tail[0]));

	cby_1__1_ cby_12__9_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_12__1__7_chany_top_out[0:19]),
		.chany_top_in(sb_12__1__8_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_140_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__140_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__140_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__140_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__140_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__140_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__140_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__140_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__140_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__140_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__140_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__140_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__140_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__140_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__140_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__140_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__140_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__140_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__140_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__140_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__140_ccff_tail[0]));

	cby_1__1_ cby_12__10_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_12__1__8_chany_top_out[0:19]),
		.chany_top_in(sb_12__1__9_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_141_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__141_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__141_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__141_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__141_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__141_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__141_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__141_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__141_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__141_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__141_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__141_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__141_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__141_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__141_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__141_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__141_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__141_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__141_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__141_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__141_ccff_tail[0]));

	cby_1__1_ cby_12__11_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_12__1__9_chany_top_out[0:19]),
		.chany_top_in(sb_12__1__10_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_142_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__142_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__142_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__142_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__142_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__142_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__142_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__142_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__142_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__142_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__142_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__142_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__142_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__142_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__142_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__142_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__142_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__142_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__142_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__142_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__142_ccff_tail[0]));

	cby_1__1_ cby_12__12_ (
		.prog_clk(prog_clk[0]),
		.chany_bottom_in(sb_12__1__10_chany_top_out[0:19]),
		.chany_top_in(sb_12__12__0_chany_bottom_out[0:19]),
		.ccff_head(grid_clb_143_ccff_tail[0]),
		.chany_bottom_out(cby_1__1__143_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__143_chany_top_out[0:19]),
		.right_grid_pin_52_(cby_1__1__143_right_grid_pin_52_[0]),
		.left_grid_pin_0_(cby_1__1__143_left_grid_pin_0_[0]),
		.left_grid_pin_1_(cby_1__1__143_left_grid_pin_1_[0]),
		.left_grid_pin_2_(cby_1__1__143_left_grid_pin_2_[0]),
		.left_grid_pin_3_(cby_1__1__143_left_grid_pin_3_[0]),
		.left_grid_pin_4_(cby_1__1__143_left_grid_pin_4_[0]),
		.left_grid_pin_5_(cby_1__1__143_left_grid_pin_5_[0]),
		.left_grid_pin_6_(cby_1__1__143_left_grid_pin_6_[0]),
		.left_grid_pin_7_(cby_1__1__143_left_grid_pin_7_[0]),
		.left_grid_pin_8_(cby_1__1__143_left_grid_pin_8_[0]),
		.left_grid_pin_9_(cby_1__1__143_left_grid_pin_9_[0]),
		.left_grid_pin_10_(cby_1__1__143_left_grid_pin_10_[0]),
		.left_grid_pin_11_(cby_1__1__143_left_grid_pin_11_[0]),
		.left_grid_pin_12_(cby_1__1__143_left_grid_pin_12_[0]),
		.left_grid_pin_13_(cby_1__1__143_left_grid_pin_13_[0]),
		.left_grid_pin_14_(cby_1__1__143_left_grid_pin_14_[0]),
		.left_grid_pin_15_(cby_1__1__143_left_grid_pin_15_[0]),
		.ccff_tail(cby_1__1__143_ccff_tail[0]));

	direct_interc direct_interc_0_ (
		.in(grid_clb_1_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_0_out[0]));

	direct_interc direct_interc_1_ (
		.in(grid_clb_2_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_1_out[0]));

	direct_interc direct_interc_2_ (
		.in(grid_clb_3_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_2_out[0]));

	direct_interc direct_interc_3_ (
		.in(grid_clb_4_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_3_out[0]));

	direct_interc direct_interc_4_ (
		.in(grid_clb_5_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_4_out[0]));

	direct_interc direct_interc_5_ (
		.in(grid_clb_6_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_5_out[0]));

	direct_interc direct_interc_6_ (
		.in(grid_clb_7_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_6_out[0]));

	direct_interc direct_interc_7_ (
		.in(grid_clb_8_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_7_out[0]));

	direct_interc direct_interc_8_ (
		.in(grid_clb_9_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_8_out[0]));

	direct_interc direct_interc_9_ (
		.in(grid_clb_10_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_9_out[0]));

	direct_interc direct_interc_10_ (
		.in(grid_clb_11_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_10_out[0]));

	direct_interc direct_interc_11_ (
		.in(grid_clb_13_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_11_out[0]));

	direct_interc direct_interc_12_ (
		.in(grid_clb_14_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_12_out[0]));

	direct_interc direct_interc_13_ (
		.in(grid_clb_15_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_13_out[0]));

	direct_interc direct_interc_14_ (
		.in(grid_clb_16_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_14_out[0]));

	direct_interc direct_interc_15_ (
		.in(grid_clb_17_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_15_out[0]));

	direct_interc direct_interc_16_ (
		.in(grid_clb_18_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_16_out[0]));

	direct_interc direct_interc_17_ (
		.in(grid_clb_19_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_17_out[0]));

	direct_interc direct_interc_18_ (
		.in(grid_clb_20_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_18_out[0]));

	direct_interc direct_interc_19_ (
		.in(grid_clb_21_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_19_out[0]));

	direct_interc direct_interc_20_ (
		.in(grid_clb_22_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_20_out[0]));

	direct_interc direct_interc_21_ (
		.in(grid_clb_23_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_21_out[0]));

	direct_interc direct_interc_22_ (
		.in(grid_clb_25_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_22_out[0]));

	direct_interc direct_interc_23_ (
		.in(grid_clb_26_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_23_out[0]));

	direct_interc direct_interc_24_ (
		.in(grid_clb_27_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_24_out[0]));

	direct_interc direct_interc_25_ (
		.in(grid_clb_28_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_25_out[0]));

	direct_interc direct_interc_26_ (
		.in(grid_clb_29_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_26_out[0]));

	direct_interc direct_interc_27_ (
		.in(grid_clb_30_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_27_out[0]));

	direct_interc direct_interc_28_ (
		.in(grid_clb_31_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_28_out[0]));

	direct_interc direct_interc_29_ (
		.in(grid_clb_32_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_29_out[0]));

	direct_interc direct_interc_30_ (
		.in(grid_clb_33_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_30_out[0]));

	direct_interc direct_interc_31_ (
		.in(grid_clb_34_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_31_out[0]));

	direct_interc direct_interc_32_ (
		.in(grid_clb_35_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_32_out[0]));

	direct_interc direct_interc_33_ (
		.in(grid_clb_37_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_33_out[0]));

	direct_interc direct_interc_34_ (
		.in(grid_clb_38_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_34_out[0]));

	direct_interc direct_interc_35_ (
		.in(grid_clb_39_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_35_out[0]));

	direct_interc direct_interc_36_ (
		.in(grid_clb_40_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_36_out[0]));

	direct_interc direct_interc_37_ (
		.in(grid_clb_41_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_37_out[0]));

	direct_interc direct_interc_38_ (
		.in(grid_clb_42_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_38_out[0]));

	direct_interc direct_interc_39_ (
		.in(grid_clb_43_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_39_out[0]));

	direct_interc direct_interc_40_ (
		.in(grid_clb_44_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_40_out[0]));

	direct_interc direct_interc_41_ (
		.in(grid_clb_45_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_41_out[0]));

	direct_interc direct_interc_42_ (
		.in(grid_clb_46_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_42_out[0]));

	direct_interc direct_interc_43_ (
		.in(grid_clb_47_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_43_out[0]));

	direct_interc direct_interc_44_ (
		.in(grid_clb_49_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_44_out[0]));

	direct_interc direct_interc_45_ (
		.in(grid_clb_50_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_45_out[0]));

	direct_interc direct_interc_46_ (
		.in(grid_clb_51_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_46_out[0]));

	direct_interc direct_interc_47_ (
		.in(grid_clb_52_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_47_out[0]));

	direct_interc direct_interc_48_ (
		.in(grid_clb_53_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_48_out[0]));

	direct_interc direct_interc_49_ (
		.in(grid_clb_54_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_49_out[0]));

	direct_interc direct_interc_50_ (
		.in(grid_clb_55_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_50_out[0]));

	direct_interc direct_interc_51_ (
		.in(grid_clb_56_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_51_out[0]));

	direct_interc direct_interc_52_ (
		.in(grid_clb_57_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_52_out[0]));

	direct_interc direct_interc_53_ (
		.in(grid_clb_58_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_53_out[0]));

	direct_interc direct_interc_54_ (
		.in(grid_clb_59_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_54_out[0]));

	direct_interc direct_interc_55_ (
		.in(grid_clb_61_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_55_out[0]));

	direct_interc direct_interc_56_ (
		.in(grid_clb_62_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_56_out[0]));

	direct_interc direct_interc_57_ (
		.in(grid_clb_63_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_57_out[0]));

	direct_interc direct_interc_58_ (
		.in(grid_clb_64_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_58_out[0]));

	direct_interc direct_interc_59_ (
		.in(grid_clb_65_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_59_out[0]));

	direct_interc direct_interc_60_ (
		.in(grid_clb_66_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_60_out[0]));

	direct_interc direct_interc_61_ (
		.in(grid_clb_67_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_61_out[0]));

	direct_interc direct_interc_62_ (
		.in(grid_clb_68_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_62_out[0]));

	direct_interc direct_interc_63_ (
		.in(grid_clb_69_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_63_out[0]));

	direct_interc direct_interc_64_ (
		.in(grid_clb_70_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_64_out[0]));

	direct_interc direct_interc_65_ (
		.in(grid_clb_71_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_65_out[0]));

	direct_interc direct_interc_66_ (
		.in(grid_clb_73_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_66_out[0]));

	direct_interc direct_interc_67_ (
		.in(grid_clb_74_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_67_out[0]));

	direct_interc direct_interc_68_ (
		.in(grid_clb_75_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_68_out[0]));

	direct_interc direct_interc_69_ (
		.in(grid_clb_76_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_69_out[0]));

	direct_interc direct_interc_70_ (
		.in(grid_clb_77_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_70_out[0]));

	direct_interc direct_interc_71_ (
		.in(grid_clb_78_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_71_out[0]));

	direct_interc direct_interc_72_ (
		.in(grid_clb_79_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_72_out[0]));

	direct_interc direct_interc_73_ (
		.in(grid_clb_80_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_73_out[0]));

	direct_interc direct_interc_74_ (
		.in(grid_clb_81_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_74_out[0]));

	direct_interc direct_interc_75_ (
		.in(grid_clb_82_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_75_out[0]));

	direct_interc direct_interc_76_ (
		.in(grid_clb_83_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_76_out[0]));

	direct_interc direct_interc_77_ (
		.in(grid_clb_85_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_77_out[0]));

	direct_interc direct_interc_78_ (
		.in(grid_clb_86_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_78_out[0]));

	direct_interc direct_interc_79_ (
		.in(grid_clb_87_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_79_out[0]));

	direct_interc direct_interc_80_ (
		.in(grid_clb_88_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_80_out[0]));

	direct_interc direct_interc_81_ (
		.in(grid_clb_89_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_81_out[0]));

	direct_interc direct_interc_82_ (
		.in(grid_clb_90_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_82_out[0]));

	direct_interc direct_interc_83_ (
		.in(grid_clb_91_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_83_out[0]));

	direct_interc direct_interc_84_ (
		.in(grid_clb_92_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_84_out[0]));

	direct_interc direct_interc_85_ (
		.in(grid_clb_93_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_85_out[0]));

	direct_interc direct_interc_86_ (
		.in(grid_clb_94_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_86_out[0]));

	direct_interc direct_interc_87_ (
		.in(grid_clb_95_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_87_out[0]));

	direct_interc direct_interc_88_ (
		.in(grid_clb_97_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_88_out[0]));

	direct_interc direct_interc_89_ (
		.in(grid_clb_98_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_89_out[0]));

	direct_interc direct_interc_90_ (
		.in(grid_clb_99_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_90_out[0]));

	direct_interc direct_interc_91_ (
		.in(grid_clb_100_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_91_out[0]));

	direct_interc direct_interc_92_ (
		.in(grid_clb_101_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_92_out[0]));

	direct_interc direct_interc_93_ (
		.in(grid_clb_102_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_93_out[0]));

	direct_interc direct_interc_94_ (
		.in(grid_clb_103_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_94_out[0]));

	direct_interc direct_interc_95_ (
		.in(grid_clb_104_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_95_out[0]));

	direct_interc direct_interc_96_ (
		.in(grid_clb_105_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_96_out[0]));

	direct_interc direct_interc_97_ (
		.in(grid_clb_106_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_97_out[0]));

	direct_interc direct_interc_98_ (
		.in(grid_clb_107_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_98_out[0]));

	direct_interc direct_interc_99_ (
		.in(grid_clb_109_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_99_out[0]));

	direct_interc direct_interc_100_ (
		.in(grid_clb_110_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_100_out[0]));

	direct_interc direct_interc_101_ (
		.in(grid_clb_111_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_101_out[0]));

	direct_interc direct_interc_102_ (
		.in(grid_clb_112_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_102_out[0]));

	direct_interc direct_interc_103_ (
		.in(grid_clb_113_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_103_out[0]));

	direct_interc direct_interc_104_ (
		.in(grid_clb_114_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_104_out[0]));

	direct_interc direct_interc_105_ (
		.in(grid_clb_115_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_105_out[0]));

	direct_interc direct_interc_106_ (
		.in(grid_clb_116_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_106_out[0]));

	direct_interc direct_interc_107_ (
		.in(grid_clb_117_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_107_out[0]));

	direct_interc direct_interc_108_ (
		.in(grid_clb_118_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_108_out[0]));

	direct_interc direct_interc_109_ (
		.in(grid_clb_119_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_109_out[0]));

	direct_interc direct_interc_110_ (
		.in(grid_clb_121_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_110_out[0]));

	direct_interc direct_interc_111_ (
		.in(grid_clb_122_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_111_out[0]));

	direct_interc direct_interc_112_ (
		.in(grid_clb_123_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_112_out[0]));

	direct_interc direct_interc_113_ (
		.in(grid_clb_124_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_113_out[0]));

	direct_interc direct_interc_114_ (
		.in(grid_clb_125_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_114_out[0]));

	direct_interc direct_interc_115_ (
		.in(grid_clb_126_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_115_out[0]));

	direct_interc direct_interc_116_ (
		.in(grid_clb_127_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_116_out[0]));

	direct_interc direct_interc_117_ (
		.in(grid_clb_128_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_117_out[0]));

	direct_interc direct_interc_118_ (
		.in(grid_clb_129_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_118_out[0]));

	direct_interc direct_interc_119_ (
		.in(grid_clb_130_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_119_out[0]));

	direct_interc direct_interc_120_ (
		.in(grid_clb_131_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_120_out[0]));

	direct_interc direct_interc_121_ (
		.in(grid_clb_133_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_121_out[0]));

	direct_interc direct_interc_122_ (
		.in(grid_clb_134_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_122_out[0]));

	direct_interc direct_interc_123_ (
		.in(grid_clb_135_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_123_out[0]));

	direct_interc direct_interc_124_ (
		.in(grid_clb_136_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_124_out[0]));

	direct_interc direct_interc_125_ (
		.in(grid_clb_137_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_125_out[0]));

	direct_interc direct_interc_126_ (
		.in(grid_clb_138_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_126_out[0]));

	direct_interc direct_interc_127_ (
		.in(grid_clb_139_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_127_out[0]));

	direct_interc direct_interc_128_ (
		.in(grid_clb_140_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_128_out[0]));

	direct_interc direct_interc_129_ (
		.in(grid_clb_141_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_129_out[0]));

	direct_interc direct_interc_130_ (
		.in(grid_clb_142_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_130_out[0]));

	direct_interc direct_interc_131_ (
		.in(grid_clb_143_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_131_out[0]));

	direct_interc direct_interc_132_ (
		.in(grid_clb_0_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_132_out[0]));

	direct_interc direct_interc_133_ (
		.in(grid_clb_12_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_133_out[0]));

	direct_interc direct_interc_134_ (
		.in(grid_clb_24_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_134_out[0]));

	direct_interc direct_interc_135_ (
		.in(grid_clb_36_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_135_out[0]));

	direct_interc direct_interc_136_ (
		.in(grid_clb_48_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_136_out[0]));

	direct_interc direct_interc_137_ (
		.in(grid_clb_60_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_137_out[0]));

	direct_interc direct_interc_138_ (
		.in(grid_clb_72_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_138_out[0]));

	direct_interc direct_interc_139_ (
		.in(grid_clb_84_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_139_out[0]));

	direct_interc direct_interc_140_ (
		.in(grid_clb_96_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_140_out[0]));

	direct_interc direct_interc_141_ (
		.in(grid_clb_108_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_141_out[0]));

	direct_interc direct_interc_142_ (
		.in(grid_clb_120_bottom_width_0_height_0__pin_50_[0]),
		.out(direct_interc_142_out[0]));

	direct_interc direct_interc_143_ (
		.in(grid_clb_1_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_143_out[0]));

	direct_interc direct_interc_144_ (
		.in(grid_clb_2_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_144_out[0]));

	direct_interc direct_interc_145_ (
		.in(grid_clb_3_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_145_out[0]));

	direct_interc direct_interc_146_ (
		.in(grid_clb_4_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_146_out[0]));

	direct_interc direct_interc_147_ (
		.in(grid_clb_5_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_147_out[0]));

	direct_interc direct_interc_148_ (
		.in(grid_clb_6_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_148_out[0]));

	direct_interc direct_interc_149_ (
		.in(grid_clb_7_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_149_out[0]));

	direct_interc direct_interc_150_ (
		.in(grid_clb_8_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_150_out[0]));

	direct_interc direct_interc_151_ (
		.in(grid_clb_9_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_151_out[0]));

	direct_interc direct_interc_152_ (
		.in(grid_clb_10_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_152_out[0]));

	direct_interc direct_interc_153_ (
		.in(grid_clb_11_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_153_out[0]));

	direct_interc direct_interc_154_ (
		.in(grid_clb_13_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_154_out[0]));

	direct_interc direct_interc_155_ (
		.in(grid_clb_14_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_155_out[0]));

	direct_interc direct_interc_156_ (
		.in(grid_clb_15_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_156_out[0]));

	direct_interc direct_interc_157_ (
		.in(grid_clb_16_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_157_out[0]));

	direct_interc direct_interc_158_ (
		.in(grid_clb_17_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_158_out[0]));

	direct_interc direct_interc_159_ (
		.in(grid_clb_18_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_159_out[0]));

	direct_interc direct_interc_160_ (
		.in(grid_clb_19_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_160_out[0]));

	direct_interc direct_interc_161_ (
		.in(grid_clb_20_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_161_out[0]));

	direct_interc direct_interc_162_ (
		.in(grid_clb_21_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_162_out[0]));

	direct_interc direct_interc_163_ (
		.in(grid_clb_22_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_163_out[0]));

	direct_interc direct_interc_164_ (
		.in(grid_clb_23_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_164_out[0]));

	direct_interc direct_interc_165_ (
		.in(grid_clb_25_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_165_out[0]));

	direct_interc direct_interc_166_ (
		.in(grid_clb_26_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_166_out[0]));

	direct_interc direct_interc_167_ (
		.in(grid_clb_27_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_167_out[0]));

	direct_interc direct_interc_168_ (
		.in(grid_clb_28_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_168_out[0]));

	direct_interc direct_interc_169_ (
		.in(grid_clb_29_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_169_out[0]));

	direct_interc direct_interc_170_ (
		.in(grid_clb_30_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_170_out[0]));

	direct_interc direct_interc_171_ (
		.in(grid_clb_31_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_171_out[0]));

	direct_interc direct_interc_172_ (
		.in(grid_clb_32_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_172_out[0]));

	direct_interc direct_interc_173_ (
		.in(grid_clb_33_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_173_out[0]));

	direct_interc direct_interc_174_ (
		.in(grid_clb_34_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_174_out[0]));

	direct_interc direct_interc_175_ (
		.in(grid_clb_35_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_175_out[0]));

	direct_interc direct_interc_176_ (
		.in(grid_clb_37_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_176_out[0]));

	direct_interc direct_interc_177_ (
		.in(grid_clb_38_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_177_out[0]));

	direct_interc direct_interc_178_ (
		.in(grid_clb_39_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_178_out[0]));

	direct_interc direct_interc_179_ (
		.in(grid_clb_40_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_179_out[0]));

	direct_interc direct_interc_180_ (
		.in(grid_clb_41_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_180_out[0]));

	direct_interc direct_interc_181_ (
		.in(grid_clb_42_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_181_out[0]));

	direct_interc direct_interc_182_ (
		.in(grid_clb_43_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_182_out[0]));

	direct_interc direct_interc_183_ (
		.in(grid_clb_44_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_183_out[0]));

	direct_interc direct_interc_184_ (
		.in(grid_clb_45_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_184_out[0]));

	direct_interc direct_interc_185_ (
		.in(grid_clb_46_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_185_out[0]));

	direct_interc direct_interc_186_ (
		.in(grid_clb_47_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_186_out[0]));

	direct_interc direct_interc_187_ (
		.in(grid_clb_49_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_187_out[0]));

	direct_interc direct_interc_188_ (
		.in(grid_clb_50_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_188_out[0]));

	direct_interc direct_interc_189_ (
		.in(grid_clb_51_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_189_out[0]));

	direct_interc direct_interc_190_ (
		.in(grid_clb_52_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_190_out[0]));

	direct_interc direct_interc_191_ (
		.in(grid_clb_53_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_191_out[0]));

	direct_interc direct_interc_192_ (
		.in(grid_clb_54_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_192_out[0]));

	direct_interc direct_interc_193_ (
		.in(grid_clb_55_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_193_out[0]));

	direct_interc direct_interc_194_ (
		.in(grid_clb_56_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_194_out[0]));

	direct_interc direct_interc_195_ (
		.in(grid_clb_57_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_195_out[0]));

	direct_interc direct_interc_196_ (
		.in(grid_clb_58_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_196_out[0]));

	direct_interc direct_interc_197_ (
		.in(grid_clb_59_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_197_out[0]));

	direct_interc direct_interc_198_ (
		.in(grid_clb_61_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_198_out[0]));

	direct_interc direct_interc_199_ (
		.in(grid_clb_62_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_199_out[0]));

	direct_interc direct_interc_200_ (
		.in(grid_clb_63_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_200_out[0]));

	direct_interc direct_interc_201_ (
		.in(grid_clb_64_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_201_out[0]));

	direct_interc direct_interc_202_ (
		.in(grid_clb_65_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_202_out[0]));

	direct_interc direct_interc_203_ (
		.in(grid_clb_66_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_203_out[0]));

	direct_interc direct_interc_204_ (
		.in(grid_clb_67_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_204_out[0]));

	direct_interc direct_interc_205_ (
		.in(grid_clb_68_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_205_out[0]));

	direct_interc direct_interc_206_ (
		.in(grid_clb_69_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_206_out[0]));

	direct_interc direct_interc_207_ (
		.in(grid_clb_70_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_207_out[0]));

	direct_interc direct_interc_208_ (
		.in(grid_clb_71_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_208_out[0]));

	direct_interc direct_interc_209_ (
		.in(grid_clb_73_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_209_out[0]));

	direct_interc direct_interc_210_ (
		.in(grid_clb_74_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_210_out[0]));

	direct_interc direct_interc_211_ (
		.in(grid_clb_75_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_211_out[0]));

	direct_interc direct_interc_212_ (
		.in(grid_clb_76_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_212_out[0]));

	direct_interc direct_interc_213_ (
		.in(grid_clb_77_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_213_out[0]));

	direct_interc direct_interc_214_ (
		.in(grid_clb_78_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_214_out[0]));

	direct_interc direct_interc_215_ (
		.in(grid_clb_79_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_215_out[0]));

	direct_interc direct_interc_216_ (
		.in(grid_clb_80_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_216_out[0]));

	direct_interc direct_interc_217_ (
		.in(grid_clb_81_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_217_out[0]));

	direct_interc direct_interc_218_ (
		.in(grid_clb_82_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_218_out[0]));

	direct_interc direct_interc_219_ (
		.in(grid_clb_83_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_219_out[0]));

	direct_interc direct_interc_220_ (
		.in(grid_clb_85_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_220_out[0]));

	direct_interc direct_interc_221_ (
		.in(grid_clb_86_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_221_out[0]));

	direct_interc direct_interc_222_ (
		.in(grid_clb_87_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_222_out[0]));

	direct_interc direct_interc_223_ (
		.in(grid_clb_88_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_223_out[0]));

	direct_interc direct_interc_224_ (
		.in(grid_clb_89_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_224_out[0]));

	direct_interc direct_interc_225_ (
		.in(grid_clb_90_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_225_out[0]));

	direct_interc direct_interc_226_ (
		.in(grid_clb_91_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_226_out[0]));

	direct_interc direct_interc_227_ (
		.in(grid_clb_92_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_227_out[0]));

	direct_interc direct_interc_228_ (
		.in(grid_clb_93_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_228_out[0]));

	direct_interc direct_interc_229_ (
		.in(grid_clb_94_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_229_out[0]));

	direct_interc direct_interc_230_ (
		.in(grid_clb_95_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_230_out[0]));

	direct_interc direct_interc_231_ (
		.in(grid_clb_97_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_231_out[0]));

	direct_interc direct_interc_232_ (
		.in(grid_clb_98_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_232_out[0]));

	direct_interc direct_interc_233_ (
		.in(grid_clb_99_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_233_out[0]));

	direct_interc direct_interc_234_ (
		.in(grid_clb_100_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_234_out[0]));

	direct_interc direct_interc_235_ (
		.in(grid_clb_101_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_235_out[0]));

	direct_interc direct_interc_236_ (
		.in(grid_clb_102_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_236_out[0]));

	direct_interc direct_interc_237_ (
		.in(grid_clb_103_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_237_out[0]));

	direct_interc direct_interc_238_ (
		.in(grid_clb_104_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_238_out[0]));

	direct_interc direct_interc_239_ (
		.in(grid_clb_105_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_239_out[0]));

	direct_interc direct_interc_240_ (
		.in(grid_clb_106_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_240_out[0]));

	direct_interc direct_interc_241_ (
		.in(grid_clb_107_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_241_out[0]));

	direct_interc direct_interc_242_ (
		.in(grid_clb_109_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_242_out[0]));

	direct_interc direct_interc_243_ (
		.in(grid_clb_110_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_243_out[0]));

	direct_interc direct_interc_244_ (
		.in(grid_clb_111_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_244_out[0]));

	direct_interc direct_interc_245_ (
		.in(grid_clb_112_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_245_out[0]));

	direct_interc direct_interc_246_ (
		.in(grid_clb_113_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_246_out[0]));

	direct_interc direct_interc_247_ (
		.in(grid_clb_114_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_247_out[0]));

	direct_interc direct_interc_248_ (
		.in(grid_clb_115_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_248_out[0]));

	direct_interc direct_interc_249_ (
		.in(grid_clb_116_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_249_out[0]));

	direct_interc direct_interc_250_ (
		.in(grid_clb_117_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_250_out[0]));

	direct_interc direct_interc_251_ (
		.in(grid_clb_118_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_251_out[0]));

	direct_interc direct_interc_252_ (
		.in(grid_clb_119_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_252_out[0]));

	direct_interc direct_interc_253_ (
		.in(grid_clb_121_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_253_out[0]));

	direct_interc direct_interc_254_ (
		.in(grid_clb_122_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_254_out[0]));

	direct_interc direct_interc_255_ (
		.in(grid_clb_123_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_255_out[0]));

	direct_interc direct_interc_256_ (
		.in(grid_clb_124_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_256_out[0]));

	direct_interc direct_interc_257_ (
		.in(grid_clb_125_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_257_out[0]));

	direct_interc direct_interc_258_ (
		.in(grid_clb_126_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_258_out[0]));

	direct_interc direct_interc_259_ (
		.in(grid_clb_127_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_259_out[0]));

	direct_interc direct_interc_260_ (
		.in(grid_clb_128_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_260_out[0]));

	direct_interc direct_interc_261_ (
		.in(grid_clb_129_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_261_out[0]));

	direct_interc direct_interc_262_ (
		.in(grid_clb_130_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_262_out[0]));

	direct_interc direct_interc_263_ (
		.in(grid_clb_131_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_263_out[0]));

	direct_interc direct_interc_264_ (
		.in(grid_clb_133_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_264_out[0]));

	direct_interc direct_interc_265_ (
		.in(grid_clb_134_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_265_out[0]));

	direct_interc direct_interc_266_ (
		.in(grid_clb_135_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_266_out[0]));

	direct_interc direct_interc_267_ (
		.in(grid_clb_136_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_267_out[0]));

	direct_interc direct_interc_268_ (
		.in(grid_clb_137_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_268_out[0]));

	direct_interc direct_interc_269_ (
		.in(grid_clb_138_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_269_out[0]));

	direct_interc direct_interc_270_ (
		.in(grid_clb_139_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_270_out[0]));

	direct_interc direct_interc_271_ (
		.in(grid_clb_140_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_271_out[0]));

	direct_interc direct_interc_272_ (
		.in(grid_clb_141_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_272_out[0]));

	direct_interc direct_interc_273_ (
		.in(grid_clb_142_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_273_out[0]));

	direct_interc direct_interc_274_ (
		.in(grid_clb_143_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_274_out[0]));

	direct_interc direct_interc_275_ (
		.in(grid_clb_0_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_275_out[0]));

	direct_interc direct_interc_276_ (
		.in(grid_clb_12_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_276_out[0]));

	direct_interc direct_interc_277_ (
		.in(grid_clb_24_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_277_out[0]));

	direct_interc direct_interc_278_ (
		.in(grid_clb_36_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_278_out[0]));

	direct_interc direct_interc_279_ (
		.in(grid_clb_48_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_279_out[0]));

	direct_interc direct_interc_280_ (
		.in(grid_clb_60_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_280_out[0]));

	direct_interc direct_interc_281_ (
		.in(grid_clb_72_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_281_out[0]));

	direct_interc direct_interc_282_ (
		.in(grid_clb_84_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_282_out[0]));

	direct_interc direct_interc_283_ (
		.in(grid_clb_96_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_283_out[0]));

	direct_interc direct_interc_284_ (
		.in(grid_clb_108_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_284_out[0]));

	direct_interc direct_interc_285_ (
		.in(grid_clb_120_bottom_width_0_height_0__pin_51_[0]),
		.out(direct_interc_285_out[0]));

endmodule
//



