//
//
//
//
//
//
module mux_tree_tapbuf_size2_mem_15 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb , VDD , VSS ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;
input  VDD ;
input  VSS ;

supply1 VDD ;
supply0 VSS ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) , 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) , 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dlygate4sd1_1 FTB_24__39 ( .A ( mem_out[1] ) , 
    .X ( net_net_59 ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_86 ( .A ( net_net_59 ) , 
    .X ( ccff_tail[0] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb , VDD , VSS ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;
input  VDD ;
input  VSS ;

supply1 VDD ;
supply0 VSS ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) , 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) , 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_23__38 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_16 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb , VDD , VSS ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;
input  VDD ;
input  VSS ;

supply1 VDD ;
supply0 VSS ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) , 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) , 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_22__37 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_14 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb , VDD , VSS ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;
input  VDD ;
input  VSS ;

supply1 VDD ;
supply0 VSS ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) , 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) , 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_21__36 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_13 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb , VDD , VSS ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;
input  VDD ;
input  VSS ;

supply1 VDD ;
supply0 VSS ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) , 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) , 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_20__35 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_12 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb , VDD , VSS ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;
input  VDD ;
input  VSS ;

supply1 VDD ;
supply0 VSS ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) , 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) , 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_19__34 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_11 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb , VDD , VSS ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;
input  VDD ;
input  VSS ;

supply1 VDD ;
supply0 VSS ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) , 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) , 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_18__33 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_10 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb , VDD , VSS ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;
input  VDD ;
input  VSS ;

supply1 VDD ;
supply0 VSS ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) , 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) , 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_17__32 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_9 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb , VDD , VSS ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;
input  VDD ;
input  VSS ;

supply1 VDD ;
supply0 VSS ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) , 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) , 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_16__31 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_8 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb , VDD , VSS ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;
input  VDD ;
input  VSS ;

supply1 VDD ;
supply0 VSS ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) , 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) , 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_15__30 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_7 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb , VDD , VSS ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;
input  VDD ;
input  VSS ;

supply1 VDD ;
supply0 VSS ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) , 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) , 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_14__29 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_6 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb , VDD , VSS ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;
input  VDD ;
input  VSS ;

supply1 VDD ;
supply0 VSS ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) , 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) , 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_13__28 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_5 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb , VDD , VSS ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;
input  VDD ;
input  VSS ;

supply1 VDD ;
supply0 VSS ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) , 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) , 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_12__27 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_4 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb , VDD , VSS ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;
input  VDD ;
input  VSS ;

supply1 VDD ;
supply0 VSS ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) , 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) , 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_11__26 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_3 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb , VDD , VSS ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;
input  VDD ;
input  VSS ;

supply1 VDD ;
supply0 VSS ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) , 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) , 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_10__25 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_2 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb , VDD , VSS ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;
input  VDD ;
input  VSS ;

supply1 VDD ;
supply0 VSS ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) , 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) , 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_9__24 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb , VDD , VSS ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;
input  VDD ;
input  VSS ;

supply1 VDD ;
supply0 VSS ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) , 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) , 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_8__23 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_0 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb , VDD , VSS ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;
input  VDD ;
input  VSS ;

supply1 VDD ;
supply0 VSS ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) , 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) , 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_7__22 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
endmodule


module mux_tree_tapbuf_size2_15 ( in , sram , sram_inv , out , VDD , VSS , 
    p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  VDD ;
input  VSS ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
supply1 VDD ;
supply0 VSS ;

sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) , .VPWR ( VDD ) , 
    .VGND ( VSS ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .VPWR ( VDD ) , 
    .VGND ( VSS ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
endmodule


module mux_tree_tapbuf_size2 ( in , sram , sram_inv , out , VDD , VSS , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  VDD ;
input  VSS ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
supply1 VDD ;
supply0 VSS ;

sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) , .VPWR ( VDD ) , 
    .VGND ( VSS ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .VPWR ( VDD ) , 
    .VGND ( VSS ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
endmodule


module mux_tree_tapbuf_size2_16 ( in , sram , sram_inv , out , VDD , VSS , 
    p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  VDD ;
input  VSS ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
supply1 VDD ;
supply0 VSS ;

sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) , .VPWR ( VDD ) , 
    .VGND ( VSS ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .VPWR ( VDD ) , 
    .VGND ( VSS ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
endmodule


module mux_tree_tapbuf_size2_14 ( in , sram , sram_inv , out , VDD , VSS , 
    p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  VDD ;
input  VSS ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
supply1 VDD ;
supply0 VSS ;

sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) , .VPWR ( VDD ) , 
    .VGND ( VSS ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .VPWR ( VDD ) , 
    .VGND ( VSS ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
endmodule


module mux_tree_tapbuf_size2_13 ( in , sram , sram_inv , out , VDD , VSS , 
    p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  VDD ;
input  VSS ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
supply1 VDD ;
supply0 VSS ;

sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) , .VPWR ( VDD ) , 
    .VGND ( VSS ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .VPWR ( VDD ) , 
    .VGND ( VSS ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
endmodule


module mux_tree_tapbuf_size2_12 ( in , sram , sram_inv , out , VDD , VSS , 
    p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  VDD ;
input  VSS ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
supply1 VDD ;
supply0 VSS ;

sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .VPWR ( VDD ) , 
    .VGND ( VSS ) ) ;
sky130_fd_sc_hd__mux2_8 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , .X ( out[0] ) , 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
endmodule


module mux_tree_tapbuf_size2_11 ( in , sram , sram_inv , out , VDD , VSS , 
    p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  VDD ;
input  VSS ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
supply1 VDD ;
supply0 VSS ;

sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) , .VPWR ( VDD ) , 
    .VGND ( VSS ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .VPWR ( VDD ) , 
    .VGND ( VSS ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
endmodule


module mux_tree_tapbuf_size2_10 ( in , sram , sram_inv , out , VDD , VSS , 
    p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  VDD ;
input  VSS ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
supply1 VDD ;
supply0 VSS ;

sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) , .VPWR ( VDD ) , 
    .VGND ( VSS ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .VPWR ( VDD ) , 
    .VGND ( VSS ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
endmodule


module mux_tree_tapbuf_size2_9 ( in , sram , sram_inv , out , VDD , VSS , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  VDD ;
input  VSS ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
supply1 VDD ;
supply0 VSS ;

sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .VPWR ( VDD ) , 
    .VGND ( VSS ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_42 ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) , .VPWR ( VDD ) , 
    .VGND ( VSS ) ) ;
endmodule


module mux_tree_tapbuf_size2_8 ( in , sram , sram_inv , out , VDD , VSS , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  VDD ;
input  VSS ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
supply1 VDD ;
supply0 VSS ;

sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) , .VPWR ( VDD ) , 
    .VGND ( VSS ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .VPWR ( VDD ) , 
    .VGND ( VSS ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
endmodule


module mux_tree_tapbuf_size2_7 ( in , sram , sram_inv , out , VDD , VSS , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  VDD ;
input  VSS ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
supply1 VDD ;
supply0 VSS ;

sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) , .VPWR ( VDD ) , 
    .VGND ( VSS ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .VPWR ( VDD ) , 
    .VGND ( VSS ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
endmodule


module mux_tree_tapbuf_size2_6 ( in , sram , sram_inv , out , VDD , VSS , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  VDD ;
input  VSS ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
supply1 VDD ;
supply0 VSS ;

sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) , .VPWR ( VDD ) , 
    .VGND ( VSS ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .VPWR ( VDD ) , 
    .VGND ( VSS ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
endmodule


module mux_tree_tapbuf_size2_5 ( in , sram , sram_inv , out , VDD , VSS , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  VDD ;
input  VSS ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
supply1 VDD ;
supply0 VSS ;

sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) , .VPWR ( VDD ) , 
    .VGND ( VSS ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .VPWR ( VDD ) , 
    .VGND ( VSS ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
endmodule


module mux_tree_tapbuf_size2_4 ( in , sram , sram_inv , out , VDD , VSS , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  VDD ;
input  VSS ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
supply1 VDD ;
supply0 VSS ;

sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) , .VPWR ( VDD ) , 
    .VGND ( VSS ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .VPWR ( VDD ) , 
    .VGND ( VSS ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
endmodule


module mux_tree_tapbuf_size2_3 ( in , sram , sram_inv , out , VDD , VSS , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  VDD ;
input  VSS ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
supply1 VDD ;
supply0 VSS ;

sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) , .VPWR ( VDD ) , 
    .VGND ( VSS ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .VPWR ( VDD ) , 
    .VGND ( VSS ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
endmodule


module mux_tree_tapbuf_size2_2 ( in , sram , sram_inv , out , VDD , VSS , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  VDD ;
input  VSS ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
supply1 VDD ;
supply0 VSS ;

sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) , .VPWR ( VDD ) , 
    .VGND ( VSS ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .VPWR ( VDD ) , 
    .VGND ( VSS ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
endmodule


module mux_tree_tapbuf_size2_1 ( in , sram , sram_inv , out , VDD , VSS , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  VDD ;
input  VSS ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
supply1 VDD ;
supply0 VSS ;

sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) , .VPWR ( VDD ) , 
    .VGND ( VSS ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .VPWR ( VDD ) , 
    .VGND ( VSS ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
endmodule


module mux_tree_tapbuf_size2_0 ( in , sram , sram_inv , out , VDD , VSS , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  VDD ;
input  VSS ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
supply1 VDD ;
supply0 VSS ;

sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) , .VPWR ( VDD ) , 
    .VGND ( VSS ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .VPWR ( VDD ) , 
    .VGND ( VSS ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
endmodule


module mux_tree_tapbuf_size3_mem_0 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb , VDD , VSS ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;
input  VDD ;
input  VSS ;

supply1 VDD ;
supply0 VSS ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) , 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) , 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_6__21 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
endmodule


module mux_tree_tapbuf_size3_mem ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb , VDD , VSS ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;
input  VDD ;
input  VSS ;

supply1 VDD ;
supply0 VSS ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) , 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) , 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_5__20 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
endmodule


module mux_tree_tapbuf_size3_0 ( in , sram , sram_inv , out , VDD , VSS , p0 ) ;
input  [0:2] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  VDD ;
input  VSS ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
supply1 VDD ;
supply0 VSS ;

sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .VPWR ( VDD ) , 
    .VGND ( VSS ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( p0 ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .VPWR ( VDD ) , 
    .VGND ( VSS ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_41 ( 
    .A ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .X ( BUF_net_41 ) , 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_P_88 ( .A ( BUF_net_41 ) , 
    .X ( out[0] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
endmodule


module mux_tree_tapbuf_size3 ( in , sram , sram_inv , out , VDD , VSS , p0 ) ;
input  [0:2] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  VDD ;
input  VSS ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
supply1 VDD ;
supply0 VSS ;

sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .X ( out[0] ) , .VPWR ( VDD ) , 
    .VGND ( VSS ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .VPWR ( VDD ) , 
    .VGND ( VSS ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( p0 ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .VPWR ( VDD ) , 
    .VGND ( VSS ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
endmodule


module mux_tree_tapbuf_size5_mem ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb , VDD , VSS ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;
input  VDD ;
input  VSS ;

supply1 VDD ;
supply0 VSS ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) , 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) , 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) , 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_4__19 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
endmodule


module mux_tree_tapbuf_size5_mem_0 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb , VDD , VSS ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;
input  VDD ;
input  VSS ;

supply1 VDD ;
supply0 VSS ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) , 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) , 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) , 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_3__18 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
endmodule


module mux_tree_tapbuf_size5 ( in , sram , sram_inv , out , VDD , VSS , p0 ) ;
input  [0:4] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  VDD ;
input  VSS ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
supply1 VDD ;
supply0 VSS ;

sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .X ( out[0] ) , .VPWR ( VDD ) , 
    .VGND ( VSS ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .VPWR ( VDD ) , 
    .VGND ( VSS ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .VPWR ( VDD ) , 
    .VGND ( VSS ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , .A1 ( in[4] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .VPWR ( VDD ) , 
    .VGND ( VSS ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
endmodule


module mux_tree_tapbuf_size5_0 ( in , sram , sram_inv , out , VDD , VSS , p0 ) ;
input  [0:4] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  VDD ;
input  VSS ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
supply1 VDD ;
supply0 VSS ;

sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .VPWR ( VDD ) , 
    .VGND ( VSS ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .VPWR ( VDD ) , 
    .VGND ( VSS ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , .A1 ( in[4] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .VPWR ( VDD ) , 
    .VGND ( VSS ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_P_87 ( 
    .A ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .X ( out[0] ) , .VPWR ( VDD ) , 
    .VGND ( VSS ) ) ;
endmodule


module mux_tree_tapbuf_size6_mem ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb , VDD , VSS ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;
input  VDD ;
input  VSS ;

supply1 VDD ;
supply0 VSS ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) , 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) , 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) , 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_2__17 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
endmodule


module mux_tree_tapbuf_size6_mem_0 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb , VDD , VSS ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;
input  VDD ;
input  VSS ;

supply1 VDD ;
supply0 VSS ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) , 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) , 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) , 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_1__16 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
endmodule


module mux_tree_tapbuf_size6 ( in , sram , sram_inv , out , VDD , VSS , p0 ) ;
input  [0:5] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  VDD ;
input  VSS ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
supply1 VDD ;
supply0 VSS ;

sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .X ( out[0] ) , .VPWR ( VDD ) , 
    .VGND ( VSS ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .VPWR ( VDD ) , 
    .VGND ( VSS ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .VPWR ( VDD ) , 
    .VGND ( VSS ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .VPWR ( VDD ) , 
    .VGND ( VSS ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
endmodule


module mux_tree_tapbuf_size6_0 ( in , sram , sram_inv , out , VDD , VSS , p0 ) ;
input  [0:5] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  VDD ;
input  VSS ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
supply1 VDD ;
supply0 VSS ;

sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .X ( out[0] ) , .VPWR ( VDD ) , 
    .VGND ( VSS ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .VPWR ( VDD ) , 
    .VGND ( VSS ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .VPWR ( VDD ) , 
    .VGND ( VSS ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .VPWR ( VDD ) , 
    .VGND ( VSS ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
endmodule


module sb_2__2_ ( prog_clk , chany_bottom_in , bottom_right_grid_pin_1_ , 
    bottom_left_grid_pin_34_ , bottom_left_grid_pin_35_ , 
    bottom_left_grid_pin_36_ , bottom_left_grid_pin_37_ , 
    bottom_left_grid_pin_38_ , bottom_left_grid_pin_39_ , 
    bottom_left_grid_pin_40_ , bottom_left_grid_pin_41_ , chanx_left_in , 
    left_top_grid_pin_1_ , ccff_head , chany_bottom_out , chanx_left_out , 
    ccff_tail , VDD , VSS ) ;
input  [0:0] prog_clk ;
input  [0:19] chany_bottom_in ;
input  [0:0] bottom_right_grid_pin_1_ ;
input  [0:0] bottom_left_grid_pin_34_ ;
input  [0:0] bottom_left_grid_pin_35_ ;
input  [0:0] bottom_left_grid_pin_36_ ;
input  [0:0] bottom_left_grid_pin_37_ ;
input  [0:0] bottom_left_grid_pin_38_ ;
input  [0:0] bottom_left_grid_pin_39_ ;
input  [0:0] bottom_left_grid_pin_40_ ;
input  [0:0] bottom_left_grid_pin_41_ ;
input  [0:19] chanx_left_in ;
input  [0:0] left_top_grid_pin_1_ ;
input  [0:0] ccff_head ;
output [0:19] chany_bottom_out ;
output [0:19] chanx_left_out ;
output [0:0] ccff_tail ;
input  VDD ;
input  VSS ;

wire [0:1] mux_tree_tapbuf_size2_0_sram ;
wire [0:1] mux_tree_tapbuf_size2_0_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_10_sram ;
wire [0:1] mux_tree_tapbuf_size2_10_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_11_sram ;
wire [0:1] mux_tree_tapbuf_size2_11_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_12_sram ;
wire [0:1] mux_tree_tapbuf_size2_12_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_13_sram ;
wire [0:1] mux_tree_tapbuf_size2_13_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_14_sram ;
wire [0:1] mux_tree_tapbuf_size2_14_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_15_sram ;
wire [0:1] mux_tree_tapbuf_size2_15_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_16_sram ;
wire [0:1] mux_tree_tapbuf_size2_16_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_17_sram ;
wire [0:1] mux_tree_tapbuf_size2_17_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_1_sram ;
wire [0:1] mux_tree_tapbuf_size2_1_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_2_sram ;
wire [0:1] mux_tree_tapbuf_size2_2_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_3_sram ;
wire [0:1] mux_tree_tapbuf_size2_3_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_4_sram ;
wire [0:1] mux_tree_tapbuf_size2_4_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_5_sram ;
wire [0:1] mux_tree_tapbuf_size2_5_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_6_sram ;
wire [0:1] mux_tree_tapbuf_size2_6_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_7_sram ;
wire [0:1] mux_tree_tapbuf_size2_7_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_8_sram ;
wire [0:1] mux_tree_tapbuf_size2_8_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_9_sram ;
wire [0:1] mux_tree_tapbuf_size2_9_sram_inv ;
wire [0:0] mux_tree_tapbuf_size2_mem_0_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_10_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_11_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_12_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_13_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_14_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_15_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_16_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_1_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_2_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_3_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_4_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_5_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_6_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_7_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_8_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_9_ccff_tail ;
wire [0:1] mux_tree_tapbuf_size3_0_sram ;
wire [0:1] mux_tree_tapbuf_size3_0_sram_inv ;
wire [0:1] mux_tree_tapbuf_size3_1_sram ;
wire [0:1] mux_tree_tapbuf_size3_1_sram_inv ;
wire [0:0] mux_tree_tapbuf_size3_mem_0_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size3_mem_1_ccff_tail ;
wire [0:2] mux_tree_tapbuf_size5_0_sram ;
wire [0:2] mux_tree_tapbuf_size5_0_sram_inv ;
wire [0:2] mux_tree_tapbuf_size5_1_sram ;
wire [0:2] mux_tree_tapbuf_size5_1_sram_inv ;
wire [0:0] mux_tree_tapbuf_size5_mem_0_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size5_mem_1_ccff_tail ;
wire [0:2] mux_tree_tapbuf_size6_0_sram ;
wire [0:2] mux_tree_tapbuf_size6_0_sram_inv ;
wire [0:2] mux_tree_tapbuf_size6_1_sram ;
wire [0:2] mux_tree_tapbuf_size6_1_sram_inv ;
wire [0:0] mux_tree_tapbuf_size6_mem_0_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size6_mem_1_ccff_tail ;
supply1 VDD ;
supply0 VSS ;
//

mux_tree_tapbuf_size6_0 mux_bottom_track_1 (
    .in ( { bottom_right_grid_pin_1_[0] , bottom_left_grid_pin_35_[0] , 
        bottom_left_grid_pin_37_[0] , bottom_left_grid_pin_39_[0] , 
        bottom_left_grid_pin_41_[0] , chanx_left_in[1] } ) ,
    .sram ( mux_tree_tapbuf_size6_0_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size6_0_sram_inv ) , 
    .out ( chany_bottom_out[0] ) , .VDD ( VDD ) , .VSS ( VSS ) , 
    .p0 ( optlc_net_114 ) ) ;
mux_tree_tapbuf_size6 mux_bottom_track_5 (
    .in ( { bottom_right_grid_pin_1_[0] , bottom_left_grid_pin_35_[0] , 
        bottom_left_grid_pin_37_[0] , bottom_left_grid_pin_39_[0] , 
        bottom_left_grid_pin_41_[0] , chanx_left_in[3] } ) ,
    .sram ( mux_tree_tapbuf_size6_1_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size6_1_sram_inv ) , 
    .out ( chany_bottom_out[2] ) , .VDD ( VDD ) , .VSS ( VSS ) , 
    .p0 ( optlc_net_114 ) ) ;
mux_tree_tapbuf_size6_mem_0 mem_bottom_track_1 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( ccff_head ) , 
    .ccff_tail ( mux_tree_tapbuf_size6_mem_0_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size6_0_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size6_0_sram_inv ) , .VDD ( VDD ) , 
    .VSS ( VSS ) ) ;
mux_tree_tapbuf_size6_mem mem_bottom_track_5 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size5_mem_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size6_mem_1_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size6_1_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size6_1_sram_inv ) , .VDD ( VDD ) , 
    .VSS ( VSS ) ) ;
mux_tree_tapbuf_size5_0 mux_bottom_track_3 (
    .in ( { bottom_left_grid_pin_34_[0] , bottom_left_grid_pin_36_[0] , 
        bottom_left_grid_pin_38_[0] , bottom_left_grid_pin_40_[0] , 
        chanx_left_in[2] } ) ,
    .sram ( mux_tree_tapbuf_size5_0_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size5_0_sram_inv ) ,
    .out ( { ropt_net_123 } ) ,
    .VDD ( VDD ) , .VSS ( VSS ) , .p0 ( optlc_net_114 ) ) ;
mux_tree_tapbuf_size5 mux_bottom_track_7 (
    .in ( { bottom_left_grid_pin_34_[0] , bottom_left_grid_pin_36_[0] , 
        bottom_left_grid_pin_38_[0] , bottom_left_grid_pin_40_[0] , 
        chanx_left_in[4] } ) ,
    .sram ( mux_tree_tapbuf_size5_1_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size5_1_sram_inv ) , 
    .out ( chany_bottom_out[3] ) , .VDD ( VDD ) , .VSS ( VSS ) , 
    .p0 ( optlc_net_114 ) ) ;
mux_tree_tapbuf_size5_mem_0 mem_bottom_track_3 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size6_mem_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size5_mem_0_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size5_0_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size5_0_sram_inv ) , .VDD ( VDD ) , 
    .VSS ( VSS ) ) ;
mux_tree_tapbuf_size5_mem mem_bottom_track_7 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size6_mem_1_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size5_mem_1_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size5_1_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size5_1_sram_inv ) , .VDD ( VDD ) , 
    .VSS ( VSS ) ) ;
mux_tree_tapbuf_size3 mux_bottom_track_9 (
    .in ( { bottom_right_grid_pin_1_[0] , bottom_left_grid_pin_41_[0] , 
        chanx_left_in[5] } ) ,
    .sram ( mux_tree_tapbuf_size3_0_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size3_0_sram_inv ) , 
    .out ( chany_bottom_out[4] ) , .VDD ( VDD ) , .VSS ( VSS ) , 
    .p0 ( optlc_net_114 ) ) ;
mux_tree_tapbuf_size3_0 mux_bottom_track_25 (
    .in ( { bottom_right_grid_pin_1_[0] , bottom_left_grid_pin_41_[0] , 
        chanx_left_in[13] } ) ,
    .sram ( mux_tree_tapbuf_size3_1_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size3_1_sram_inv ) ,
    .out ( { ropt_net_130 } ) ,
    .VDD ( VDD ) , .VSS ( VSS ) , .p0 ( optlc_net_115 ) ) ;
mux_tree_tapbuf_size3_mem mem_bottom_track_9 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size5_mem_1_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size3_mem_0_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size3_0_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size3_0_sram_inv ) , .VDD ( VDD ) , 
    .VSS ( VSS ) ) ;
mux_tree_tapbuf_size3_mem_0 mem_bottom_track_25 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_6_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size3_mem_1_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size3_1_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size3_1_sram_inv ) , .VDD ( VDD ) , 
    .VSS ( VSS ) ) ;
mux_tree_tapbuf_size2_0 mux_bottom_track_11 (
    .in ( { bottom_left_grid_pin_34_[0] , chanx_left_in[6] } ) ,
    .sram ( mux_tree_tapbuf_size2_0_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_0_sram_inv ) , 
    .out ( chany_bottom_out[5] ) , .VDD ( VDD ) , .VSS ( VSS ) , 
    .p0 ( optlc_net_114 ) ) ;
mux_tree_tapbuf_size2_1 mux_bottom_track_13 (
    .in ( { bottom_left_grid_pin_35_[0] , chanx_left_in[7] } ) ,
    .sram ( mux_tree_tapbuf_size2_1_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_1_sram_inv ) , 
    .out ( chany_bottom_out[6] ) , .VDD ( VDD ) , .VSS ( VSS ) , 
    .p0 ( optlc_net_115 ) ) ;
mux_tree_tapbuf_size2_2 mux_bottom_track_15 (
    .in ( { bottom_left_grid_pin_36_[0] , chanx_left_in[8] } ) ,
    .sram ( mux_tree_tapbuf_size2_2_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_2_sram_inv ) , 
    .out ( chany_bottom_out[7] ) , .VDD ( VDD ) , .VSS ( VSS ) , 
    .p0 ( optlc_net_115 ) ) ;
mux_tree_tapbuf_size2_3 mux_bottom_track_17 (
    .in ( { bottom_left_grid_pin_37_[0] , chanx_left_in[9] } ) ,
    .sram ( mux_tree_tapbuf_size2_3_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_3_sram_inv ) , 
    .out ( chany_bottom_out[8] ) , .VDD ( VDD ) , .VSS ( VSS ) , 
    .p0 ( optlc_net_112 ) ) ;
mux_tree_tapbuf_size2_4 mux_bottom_track_19 (
    .in ( { bottom_left_grid_pin_38_[0] , chanx_left_in[10] } ) ,
    .sram ( mux_tree_tapbuf_size2_4_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_4_sram_inv ) , 
    .out ( chany_bottom_out[9] ) , .VDD ( VDD ) , .VSS ( VSS ) , 
    .p0 ( optlc_net_114 ) ) ;
mux_tree_tapbuf_size2_5 mux_bottom_track_21 (
    .in ( { bottom_left_grid_pin_39_[0] , chanx_left_in[11] } ) ,
    .sram ( mux_tree_tapbuf_size2_5_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_5_sram_inv ) , 
    .out ( chany_bottom_out[10] ) , .VDD ( VDD ) , .VSS ( VSS ) , 
    .p0 ( optlc_net_115 ) ) ;
mux_tree_tapbuf_size2_6 mux_bottom_track_23 (
    .in ( { bottom_left_grid_pin_40_[0] , chanx_left_in[12] } ) ,
    .sram ( mux_tree_tapbuf_size2_6_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_6_sram_inv ) , 
    .out ( chany_bottom_out[11] ) , .VDD ( VDD ) , .VSS ( VSS ) , 
    .p0 ( optlc_net_113 ) ) ;
mux_tree_tapbuf_size2_7 mux_bottom_track_27 (
    .in ( { bottom_left_grid_pin_34_[0] , chanx_left_in[14] } ) ,
    .sram ( mux_tree_tapbuf_size2_7_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_7_sram_inv ) , 
    .out ( chany_bottom_out[13] ) , .VDD ( VDD ) , .VSS ( VSS ) , 
    .p0 ( optlc_net_114 ) ) ;
mux_tree_tapbuf_size2_8 mux_bottom_track_29 (
    .in ( { bottom_left_grid_pin_35_[0] , chanx_left_in[15] } ) ,
    .sram ( mux_tree_tapbuf_size2_8_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_8_sram_inv ) , 
    .out ( chany_bottom_out[14] ) , .VDD ( VDD ) , .VSS ( VSS ) , 
    .p0 ( optlc_net_115 ) ) ;
mux_tree_tapbuf_size2_9 mux_bottom_track_31 (
    .in ( { bottom_left_grid_pin_36_[0] , chanx_left_in[16] } ) ,
    .sram ( mux_tree_tapbuf_size2_9_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_9_sram_inv ) ,
    .out ( { ropt_net_120 } ) ,
    .VDD ( VDD ) , .VSS ( VSS ) , .p0 ( optlc_net_115 ) ) ;
mux_tree_tapbuf_size2_10 mux_bottom_track_33 (
    .in ( { bottom_left_grid_pin_37_[0] , chanx_left_in[17] } ) ,
    .sram ( mux_tree_tapbuf_size2_10_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_10_sram_inv ) , 
    .out ( chany_bottom_out[16] ) , .VDD ( VDD ) , .VSS ( VSS ) , 
    .p0 ( optlc_net_112 ) ) ;
mux_tree_tapbuf_size2_11 mux_bottom_track_35 (
    .in ( { bottom_left_grid_pin_38_[0] , chanx_left_in[18] } ) ,
    .sram ( mux_tree_tapbuf_size2_11_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_11_sram_inv ) , 
    .out ( chany_bottom_out[17] ) , .VDD ( VDD ) , .VSS ( VSS ) , 
    .p0 ( optlc_net_112 ) ) ;
mux_tree_tapbuf_size2_12 mux_bottom_track_37 (
    .in ( { bottom_left_grid_pin_39_[0] , chanx_left_in[19] } ) ,
    .sram ( mux_tree_tapbuf_size2_12_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_12_sram_inv ) , 
    .out ( chany_bottom_out[18] ) , .VDD ( VDD ) , .VSS ( VSS ) , 
    .p0 ( optlc_net_115 ) ) ;
mux_tree_tapbuf_size2_13 mux_bottom_track_39 (
    .in ( { bottom_left_grid_pin_40_[0] , chanx_left_in[0] } ) ,
    .sram ( mux_tree_tapbuf_size2_13_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_13_sram_inv ) , 
    .out ( chany_bottom_out[19] ) , .VDD ( VDD ) , .VSS ( VSS ) , 
    .p0 ( optlc_net_114 ) ) ;
mux_tree_tapbuf_size2_14 mux_left_track_1 (
    .in ( { chany_bottom_in[19] , left_top_grid_pin_1_[0] } ) ,
    .sram ( mux_tree_tapbuf_size2_14_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_14_sram_inv ) , 
    .out ( chanx_left_out[0] ) , .VDD ( VDD ) , .VSS ( VSS ) , 
    .p0 ( optlc_net_113 ) ) ;
mux_tree_tapbuf_size2_16 mux_left_track_5 (
    .in ( { chany_bottom_in[1] , left_top_grid_pin_1_[0] } ) ,
    .sram ( mux_tree_tapbuf_size2_15_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_15_sram_inv ) , 
    .out ( chanx_left_out[2] ) , .VDD ( VDD ) , .VSS ( VSS ) , 
    .p0 ( optlc_net_113 ) ) ;
mux_tree_tapbuf_size2 mux_left_track_9 (
    .in ( { chany_bottom_in[3] , left_top_grid_pin_1_[0] } ) ,
    .sram ( mux_tree_tapbuf_size2_16_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_16_sram_inv ) , 
    .out ( chanx_left_out[4] ) , .VDD ( VDD ) , .VSS ( VSS ) , 
    .p0 ( optlc_net_113 ) ) ;
mux_tree_tapbuf_size2_15 mux_left_track_25 (
    .in ( { chany_bottom_in[11] , left_top_grid_pin_1_[0] } ) ,
    .sram ( mux_tree_tapbuf_size2_17_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_17_sram_inv ) , 
    .out ( chanx_left_out[12] ) , .VDD ( VDD ) , .VSS ( VSS ) , 
    .p0 ( optlc_net_113 ) ) ;
mux_tree_tapbuf_size2_mem_0 mem_bottom_track_11 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size3_mem_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_0_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_0_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_0_sram_inv ) , .VDD ( VDD ) , 
    .VSS ( VSS ) ) ;
mux_tree_tapbuf_size2_mem_1 mem_bottom_track_13 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_1_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_1_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_1_sram_inv ) , .VDD ( VDD ) , 
    .VSS ( VSS ) ) ;
mux_tree_tapbuf_size2_mem_2 mem_bottom_track_15 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_1_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_2_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_2_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_2_sram_inv ) , .VDD ( VDD ) , 
    .VSS ( VSS ) ) ;
mux_tree_tapbuf_size2_mem_3 mem_bottom_track_17 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_2_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_3_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_3_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_3_sram_inv ) , .VDD ( VDD ) , 
    .VSS ( VSS ) ) ;
mux_tree_tapbuf_size2_mem_4 mem_bottom_track_19 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_3_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_4_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_4_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_4_sram_inv ) , .VDD ( VDD ) , 
    .VSS ( VSS ) ) ;
mux_tree_tapbuf_size2_mem_5 mem_bottom_track_21 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_4_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_5_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_5_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_5_sram_inv ) , .VDD ( VDD ) , 
    .VSS ( VSS ) ) ;
mux_tree_tapbuf_size2_mem_6 mem_bottom_track_23 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_5_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_6_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_6_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_6_sram_inv ) , .VDD ( VDD ) , 
    .VSS ( VSS ) ) ;
mux_tree_tapbuf_size2_mem_7 mem_bottom_track_27 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size3_mem_1_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_7_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_7_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_7_sram_inv ) , .VDD ( VDD ) , 
    .VSS ( VSS ) ) ;
mux_tree_tapbuf_size2_mem_8 mem_bottom_track_29 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_7_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_8_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_8_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_8_sram_inv ) , .VDD ( VDD ) , 
    .VSS ( VSS ) ) ;
mux_tree_tapbuf_size2_mem_9 mem_bottom_track_31 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_8_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_9_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_9_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_9_sram_inv ) , .VDD ( VDD ) , 
    .VSS ( VSS ) ) ;
mux_tree_tapbuf_size2_mem_10 mem_bottom_track_33 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_9_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_10_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_10_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_10_sram_inv ) , .VDD ( VDD ) , 
    .VSS ( VSS ) ) ;
mux_tree_tapbuf_size2_mem_11 mem_bottom_track_35 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_10_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_11_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_11_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_11_sram_inv ) , .VDD ( VDD ) , 
    .VSS ( VSS ) ) ;
mux_tree_tapbuf_size2_mem_12 mem_bottom_track_37 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_11_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_12_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_12_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_12_sram_inv ) , .VDD ( VDD ) , 
    .VSS ( VSS ) ) ;
mux_tree_tapbuf_size2_mem_13 mem_bottom_track_39 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_12_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_13_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_13_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_13_sram_inv ) , .VDD ( VDD ) , 
    .VSS ( VSS ) ) ;
mux_tree_tapbuf_size2_mem_14 mem_left_track_1 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_13_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_14_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_14_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_14_sram_inv ) , .VDD ( VDD ) , 
    .VSS ( VSS ) ) ;
mux_tree_tapbuf_size2_mem_16 mem_left_track_5 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_14_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_15_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_15_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_15_sram_inv ) , .VDD ( VDD ) , 
    .VSS ( VSS ) ) ;
mux_tree_tapbuf_size2_mem mem_left_track_9 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_15_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_16_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_16_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_16_sram_inv ) , .VDD ( VDD ) , 
    .VSS ( VSS ) ) ;
mux_tree_tapbuf_size2_mem_15 mem_left_track_25 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_16_ccff_tail ) ,
    .ccff_tail ( { ropt_net_128 } ) ,
    .mem_out ( mux_tree_tapbuf_size2_17_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_17_sram_inv ) , .VDD ( VDD ) , 
    .VSS ( VSS ) ) ;
sky130_fd_sc_hd__tap_2 tapfiller_sky130_fd_sc_hd__tap_2_2401 ( .VNB ( VSS ) , 
    .VPB ( VDD ) , .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__tap_2 tapfiller_sky130_fd_sc_hd__tap_2_2402 ( .VNB ( VSS ) , 
    .VPB ( VDD ) , .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__tap_2 tapfiller_sky130_fd_sc_hd__tap_2_2403 ( .VNB ( VSS ) , 
    .VPB ( VDD ) , .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__tap_2 tapfiller_sky130_fd_sc_hd__tap_2_2404 ( .VNB ( VSS ) , 
    .VPB ( VDD ) , .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__tap_2 tapfiller_sky130_fd_sc_hd__tap_2_2405 ( .VNB ( VSS ) , 
    .VPB ( VDD ) , .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__tap_2 tapfiller_sky130_fd_sc_hd__tap_2_2406 ( .VNB ( VSS ) , 
    .VPB ( VDD ) , .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__tap_2 tapfiller_sky130_fd_sc_hd__tap_2_2407 ( .VNB ( VSS ) , 
    .VPB ( VDD ) , .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__tap_2 tapfiller_sky130_fd_sc_hd__tap_2_2408 ( .VNB ( VSS ) , 
    .VPB ( VDD ) , .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__tap_2 tapfiller_sky130_fd_sc_hd__tap_2_2409 ( .VNB ( VSS ) , 
    .VPB ( VDD ) , .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__tap_2 tapfiller_sky130_fd_sc_hd__tap_2_2410 ( .VNB ( VSS ) , 
    .VPB ( VDD ) , .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__tap_2 tapfiller_sky130_fd_sc_hd__tap_2_2411 ( .VNB ( VSS ) , 
    .VPB ( VDD ) , .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__tap_2 tapfiller_sky130_fd_sc_hd__tap_2_2412 ( .VNB ( VSS ) , 
    .VPB ( VDD ) , .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__tap_2 tapfiller_sky130_fd_sc_hd__tap_2_2413 ( .VNB ( VSS ) , 
    .VPB ( VDD ) , .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__tap_2 tapfiller_sky130_fd_sc_hd__tap_2_2414 ( .VNB ( VSS ) , 
    .VPB ( VDD ) , .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__tap_2 tapfiller_sky130_fd_sc_hd__tap_2_2415 ( .VNB ( VSS ) , 
    .VPB ( VDD ) , .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__tap_2 tapfiller_sky130_fd_sc_hd__tap_2_2416 ( .VNB ( VSS ) , 
    .VPB ( VDD ) , .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__conb_1 optlc_107 ( .LO ( SYNOPSYS_UNCONNECTED_1 ) , 
    .HI ( optlc_net_112 ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__conb_1 optlc_109 ( .LO ( SYNOPSYS_UNCONNECTED_2 ) , 
    .HI ( optlc_net_113 ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__conb_1 optlc_111 ( .LO ( SYNOPSYS_UNCONNECTED_3 ) , 
    .HI ( optlc_net_114 ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__conb_1 optlc_113 ( .LO ( SYNOPSYS_UNCONNECTED_4 ) , 
    .HI ( optlc_net_115 ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_703 ( .A ( chany_bottom_in[2] ) , 
    .X ( chanx_left_out[3] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_704 ( .A ( chany_bottom_in[7] ) , 
    .X ( ropt_net_138 ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_705 ( 
    .A ( chany_bottom_in[16] ) , .X ( chanx_left_out[17] ) , .VPWR ( VDD ) , 
    .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_706 ( .A ( ropt_net_120 ) , 
    .X ( ropt_net_137 ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_707 ( 
    .A ( chany_bottom_in[17] ) , .X ( chanx_left_out[18] ) , .VPWR ( VDD ) , 
    .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_708 ( .A ( chany_bottom_in[8] ) , 
    .X ( chanx_left_out[9] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_709 ( .A ( ropt_net_123 ) , 
    .X ( ropt_net_141 ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_710 ( 
    .A ( chany_bottom_in[15] ) , .X ( ropt_net_135 ) , .VPWR ( VDD ) , 
    .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_711 ( .A ( chany_bottom_in[0] ) , 
    .X ( chanx_left_out[1] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_712 ( 
    .A ( chany_bottom_in[12] ) , .X ( ropt_net_134 ) , .VPWR ( VDD ) , 
    .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_719 ( .A ( ropt_net_133 ) , 
    .X ( chanx_left_out[6] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_713 ( 
    .A ( chany_bottom_in[18] ) , .X ( chanx_left_out[19] ) , .VPWR ( VDD ) , 
    .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_714 ( .A ( ropt_net_128 ) , 
    .X ( ropt_net_140 ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_715 ( .A ( ropt_net_129 ) , 
    .X ( ropt_net_136 ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_46 ( .A ( chany_bottom_in[4] ) , 
    .X ( BUF_net_46 ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_47 ( .A ( chany_bottom_in[5] ) , 
    .X ( ropt_net_131 ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_716 ( .A ( ropt_net_130 ) , 
    .X ( chany_bottom_out[12] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_720 ( .A ( ropt_net_134 ) , 
    .X ( chanx_left_out[13] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_721 ( .A ( ropt_net_135 ) , 
    .X ( chanx_left_out[16] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_51 ( .A ( chany_bottom_in[9] ) , 
    .X ( BUF_net_51 ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_52 ( .A ( chany_bottom_in[10] ) , 
    .X ( BUF_net_52 ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_722 ( .A ( ropt_net_136 ) , 
    .X ( chanx_left_out[7] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_54 ( .A ( chany_bottom_in[13] ) , 
    .X ( BUF_net_54 ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_55 ( .A ( chany_bottom_in[14] ) , 
    .X ( BUF_net_55 ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_718 ( .A ( ropt_net_131 ) , 
    .X ( ropt_net_133 ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_723 ( .A ( ropt_net_137 ) , 
    .X ( chany_bottom_out[15] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_724 ( .A ( ropt_net_138 ) , 
    .X ( chanx_left_out[8] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_725 ( .A ( ropt_net_139 ) , 
    .X ( chanx_left_out[5] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_726 ( .A ( ropt_net_140 ) , 
    .X ( ccff_tail[0] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_727 ( .A ( ropt_net_141 ) , 
    .X ( chany_bottom_out[1] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x184000y0 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x220800y0 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x257600y0 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x294400y0 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x331200y0 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x368000y0 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x404800y0 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x441600y0 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x460000y0 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x469200y0 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x483000y0 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 BUFT_P_93 ( .A ( BUF_net_46 ) , 
    .X ( ropt_net_139 ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x519800y0 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_P_95 ( .A ( chany_bottom_in[6] ) , 
    .X ( ropt_net_129 ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x556600y0 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x593400y0 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 BUFT_P_98 ( .A ( BUF_net_51 ) , 
    .X ( chanx_left_out[10] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 BUFT_P_99 ( .A ( BUF_net_52 ) , 
    .X ( chanx_left_out[11] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x630200y0 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 BUFT_P_101 ( .A ( BUF_net_54 ) , 
    .X ( chanx_left_out[14] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 BUFT_P_102 ( .A ( BUF_net_55 ) , 
    .X ( chanx_left_out[15] ) , .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x667000y0 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x703800y0 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x740600y0 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x777400y0 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x814200y0 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x832600y0 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x841800y0 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x184000y27200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x220800y27200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x239200y27200 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x285200y27200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x414000y27200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x423200y27200 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x680800y27200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x690000y27200 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x722200y27200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x759000y27200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x795800y27200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x832600y27200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x841800y27200 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x184000y54400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x220800y54400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x257600y54400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x312800y54400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x349600y54400 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x395600y54400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x414000y54400 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x657800y54400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x694600y54400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x759000y54400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x795800y54400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x832600y54400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x841800y54400 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x184000y81600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x202400y81600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x340400y81600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x358800y81600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x368000y81600 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x469200y81600 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x510600y81600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x519800y81600 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x552000y81600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x588800y81600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x625600y81600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x662400y81600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x726800y81600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x763600y81600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x800400y81600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x837200y81600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x184000y108800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x220800y108800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x239200y108800 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x285200y108800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x322000y108800 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x368000y108800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x492200y108800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x529000y108800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x547400y108800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x598000y108800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x607200y108800 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x639400y108800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x676200y108800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x713000y108800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x749800y108800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x795800y108800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x832600y108800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x841800y108800 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x184000y136000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x202400y136000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x253000y136000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x289800y136000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x386400y136000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x423200y136000 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x464600y136000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x483000y136000 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x529000y136000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x565800y136000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x575000y136000 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x667000y136000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x703800y136000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x800400y136000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x837200y136000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x0y163200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x36800y163200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x73600y163200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x110400y163200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x147200y163200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x184000y163200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x220800y163200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x239200y163200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x289800y163200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x308200y163200 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x400200y163200 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x492200y163200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x529000y163200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x565800y163200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x575000y163200 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x616400y163200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x634800y163200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x644000y163200 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x690000y163200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x726800y163200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x745200y163200 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x791200y163200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x828000y163200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x0y190400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x18400y190400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x197800y190400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x234600y190400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x271400y190400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x289800y190400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x340400y190400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x377200y190400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x483000y190400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x519800y190400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x529000y190400 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x621000y190400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x657800y190400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x694600y190400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x731400y190400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x768200y190400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x805000y190400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x841800y190400 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x0y217600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x18400y217600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x239200y217600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x299000y217600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x317400y217600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x326600y217600 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x414000y217600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x450800y217600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x487600y217600 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x529000y217600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x565800y217600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x602600y217600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x639400y217600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x676200y217600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x685400y217600 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x731400y217600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x768200y217600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x805000y217600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x841800y217600 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x0y244800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x18400y244800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x156400y244800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x193200y244800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x211600y244800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x220800y244800 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x266800y244800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x285200y244800 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x331200y244800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x368000y244800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x404800y244800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x464600y244800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x483000y244800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x519800y244800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x538200y244800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x634800y244800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x671600y244800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x690000y244800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x699200y244800 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x791200y244800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x828000y244800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x0y272000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x18400y272000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x161000y272000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x197800y272000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x331200y272000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x381800y272000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x400200y272000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x450800y272000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x469200y272000 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x515200y272000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x533600y272000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x542800y272000 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x584200y272000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x621000y272000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x657800y272000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x676200y272000 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x768200y272000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x805000y272000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x841800y272000 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x0y299200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x18400y299200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x82800y299200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x119600y299200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x128800y299200 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x174800y299200 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x220800y299200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x230000y299200 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x271400y299200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x308200y299200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x340400y299200 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x432400y299200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x469200y299200 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x483000y299200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x519800y299200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x538200y299200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x584200y299200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x621000y299200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x657800y299200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x694600y299200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x731400y299200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x768200y299200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x805000y299200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x841800y299200 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x0y326400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x18400y326400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x368000y326400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x386400y326400 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x478400y326400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x515200y326400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x621000y326400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x657800y326400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x782000y326400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x818800y326400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x837200y326400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x0y353600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x18400y353600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x73600y353600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x82800y353600 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x165600y353600 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x202400y353600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x239200y353600 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x285200y353600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x335800y353600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x395600y353600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x414000y353600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x460000y353600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x469200y353600 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x483000y353600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x501400y353600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x607200y353600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x644000y353600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x653200y353600 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x745200y353600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x782000y353600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x818800y353600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x837200y353600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x0y380800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x18400y380800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x73600y380800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x82800y380800 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x151800y380800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x170200y380800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x253000y380800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x289800y380800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x326600y380800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x363400y380800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x460000y380800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x496800y380800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x533600y380800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x570400y380800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x607200y380800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x644000y380800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x680800y380800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x717600y380800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x754400y380800 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x795800y380800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x832600y380800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x841800y380800 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x0y408000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x18400y408000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x193200y408000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x211600y408000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x220800y408000 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x266800y408000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x276000y408000 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x322000y408000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x358800y408000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x395600y408000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x432400y408000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x469200y408000 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x483000y408000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x561200y408000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x598000y408000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x634800y408000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x671600y408000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x680800y408000 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x772800y408000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x809600y408000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x0y435200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x18400y435200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x248400y435200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x285200y435200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x322000y435200 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x414000y435200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x450800y435200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x575000y435200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x611800y435200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x648600y435200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x667000y435200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x676200y435200 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x768200y435200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x805000y435200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x841800y435200 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x0y462400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x18400y462400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x161000y462400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x197800y462400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x216200y462400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x312800y462400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x349600y462400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x386400y462400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x464600y462400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x483000y462400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x533600y462400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x570400y462400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x607200y462400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x644000y462400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x680800y462400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x717600y462400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x754400y462400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x791200y462400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x828000y462400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x0y489600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x18400y489600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x110400y489600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x128800y489600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x216200y489600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x234600y489600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x280600y489600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x317400y489600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x368000y489600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x404800y489600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x441600y489600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x478400y489600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x515200y489600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x593400y489600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x630200y489600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x667000y489600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x703800y489600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x777400y489600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x814200y489600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x832600y489600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x841800y489600 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x0y516800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x18400y516800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x73600y516800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x193200y516800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x299000y516800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x400200y516800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x437000y516800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x483000y516800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x542800y516800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x579600y516800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x616400y516800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x653200y516800 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x699200y516800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x736000y516800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x772800y516800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x809600y516800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x0y544000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x18400y544000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x55200y544000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x161000y544000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x197800y544000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x234600y544000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x271400y544000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x308200y544000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x317400y544000 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x409400y544000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x446200y544000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x542800y544000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x579600y544000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x616400y544000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x653200y544000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x662400y544000 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x708400y544000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x745200y544000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x782000y544000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x818800y544000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x837200y544000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x0y571200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x18400y571200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x202400y571200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x308200y571200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x326600y571200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x335800y571200 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x377200y571200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x414000y571200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x450800y571200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x469200y571200 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x483000y571200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x519800y571200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x556600y571200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x653200y571200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x699200y571200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x736000y571200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x772800y571200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x809600y571200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x0y598400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x18400y598400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x161000y598400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x197800y598400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x234600y598400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x253000y598400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x262200y598400 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x345000y598400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x381800y598400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x400200y598400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x409400y598400 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x501400y598400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x519800y598400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x529000y598400 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x575000y598400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x680800y598400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x717600y598400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x754400y598400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x791200y598400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x828000y598400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x0y625600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x18400y625600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x151800y625600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x188600y625600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x225400y625600 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x271400y625600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x395600y625600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x469200y625600 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x483000y625600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x519800y625600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x556600y625600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x593400y625600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x630200y625600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x648600y625600 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x690000y625600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x726800y625600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x763600y625600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x800400y625600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x837200y625600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x0y652800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x18400y652800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x119600y652800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x128800y652800 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x174800y652800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x211600y652800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x230000y652800 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x322000y652800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x427800y652800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x464600y652800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x501400y652800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x579600y652800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x616400y652800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x713000y652800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x749800y652800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x786600y652800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x823400y652800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x841800y652800 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x0y680000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x18400y680000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x161000y680000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x197800y680000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x234600y680000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x253000y680000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x299000y680000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x335800y680000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x372600y680000 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x418600y680000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x455400y680000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x483000y680000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x501400y680000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x598000y680000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x634800y680000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x671600y680000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x708400y680000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x745200y680000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x782000y680000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x818800y680000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x837200y680000 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x0y707200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x18400y707200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x161000y707200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x197800y707200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x234600y707200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x340400y707200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x358800y707200 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x450800y707200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x487600y707200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x584200y707200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x621000y707200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x657800y707200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x694600y707200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x731400y707200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x768200y707200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x805000y707200 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x841800y707200 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x0y734400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x18400y734400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x73600y734400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x207000y734400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x243800y734400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x280600y734400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x317400y734400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x354200y734400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x391000y734400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x427800y734400 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x483000y734400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x519800y734400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x556600y734400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x593400y734400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x630200y734400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x667000y734400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x703800y734400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x740600y734400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x777400y734400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x814200y734400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x832600y734400 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x841800y734400 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x0y761600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x18400y761600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x105800y761600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x142600y761600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x179400y761600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x216200y761600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x253000y761600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x289800y761600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x326600y761600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x363400y761600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x400200y761600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x437000y761600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x510600y761600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x547400y761600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x584200y761600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x621000y761600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x657800y761600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x694600y761600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x731400y761600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x768200y761600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x805000y761600 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x841800y761600 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x0y788800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x36800y788800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x73600y788800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x110400y788800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x147200y788800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x184000y788800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x220800y788800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x257600y788800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x294400y788800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x331200y788800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x368000y788800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x404800y788800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x441600y788800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x460000y788800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x469200y788800 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x483000y788800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x519800y788800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x556600y788800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x593400y788800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x630200y788800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x667000y788800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x703800y788800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x740600y788800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_8 xofiller_sky130_fd_sc_hd__fill_8_x777400y788800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_4 xofiller_sky130_fd_sc_hd__fill_4_x814200y788800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_2 xofiller_sky130_fd_sc_hd__fill_2_x832600y788800 ( 
    .VGND ( VSS ) , .VPWR ( VDD ) ) ;
sky130_fd_sc_hd__fill_1 xofiller_sky130_fd_sc_hd__fill_1_x841800y788800 ( 
    .VPWR ( VDD ) , .VGND ( VSS ) ) ;
endmodule


