VERSION 5.7 ;
BUSBITCHARS "[]" ;

UNITS
  DATABASE MICRONS 1000 ;
END UNITS

MANUFACTURINGGRID 0.005 ;

LAYER li1
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.46 ;
  WIDTH 0.17 ;
END li1

LAYER mcon
  TYPE CUT ;
END mcon

LAYER met1
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.34 ;
  WIDTH 0.14 ;
END met1

LAYER via
  TYPE CUT ;
END via

LAYER met2
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.46 ;
  WIDTH 0.14 ;
END met2

LAYER via2
  TYPE CUT ;
END via2

LAYER met3
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.68 ;
  WIDTH 0.3 ;
END met3

LAYER via3
  TYPE CUT ;
END via3

LAYER met4
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.92 ;
  WIDTH 0.3 ;
END met4

LAYER via4
  TYPE CUT ;
END via4

LAYER met5
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 3.4 ;
  WIDTH 1.6 ;
END met5

LAYER nwell
  TYPE MASTERSLICE ;
END nwell

LAYER pwell
  TYPE MASTERSLICE ;
END pwell

LAYER OVERLAP
  TYPE OVERLAP ;
END OVERLAP

VIA L1M1_PR
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.145 -0.115 0.145 0.115 ;
END L1M1_PR

VIA L1M1_PR_R
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.115 -0.145 0.115 0.145 ;
END L1M1_PR_R

VIA L1M1_PR_M
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.115 -0.145 0.115 0.145 ;
END L1M1_PR_M

VIA L1M1_PR_MR
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.145 -0.115 0.145 0.115 ;
END L1M1_PR_MR

VIA L1M1_PR_C
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.145 -0.145 0.145 0.145 ;
END L1M1_PR_C

VIA M1M2_PR
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR

VIA M1M2_PR_Enc
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_Enc

VIA M1M2_PR_R
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_R

VIA M1M2_PR_R_Enc
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR_R_Enc

VIA M1M2_PR_M
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_M

VIA M1M2_PR_M_Enc
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR_M_Enc

VIA M1M2_PR_MR
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR_MR

VIA M1M2_PR_MR_Enc
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_MR_Enc

VIA M1M2_PR_C
  LAYER met1 ;
    RECT -0.16 -0.16 0.16 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.16 0.16 0.16 ;
END M1M2_PR_C

VIA M2M3_PR
  LAYER met2 ;
    RECT -0.14 -0.185 0.14 0.185 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR

VIA M2M3_PR_R
  LAYER met2 ;
    RECT -0.185 -0.14 0.185 0.14 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_R

VIA M2M3_PR_M
  LAYER met2 ;
    RECT -0.14 -0.185 0.14 0.185 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_M

VIA M2M3_PR_MR
  LAYER met2 ;
    RECT -0.185 -0.14 0.185 0.14 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_MR

VIA M2M3_PR_C
  LAYER met2 ;
    RECT -0.185 -0.185 0.185 0.185 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_C

VIA M3M4_PR
  LAYER met3 ;
    RECT -0.19 -0.16 0.19 0.16 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR

VIA M3M4_PR_R
  LAYER met3 ;
    RECT -0.16 -0.19 0.16 0.19 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_R

VIA M3M4_PR_M
  LAYER met3 ;
    RECT -0.19 -0.16 0.19 0.16 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_M

VIA M3M4_PR_MR
  LAYER met3 ;
    RECT -0.16 -0.19 0.16 0.19 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_MR

VIA M3M4_PR_C
  LAYER met3 ;
    RECT -0.19 -0.19 0.19 0.19 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_C

VIA M4M5_PR
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR

VIA M4M5_PR_R
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_R

VIA M4M5_PR_M
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_M

VIA M4M5_PR_MR
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_MR

VIA M4M5_PR_C
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_C

SITE unit
  CLASS CORE ;
  SYMMETRY Y ;
  SIZE 0.46 BY 2.72 ;
END unit

SITE unithddbl
  CLASS CORE ;
  SIZE 0.46 BY 5.44 ;
END unithddbl

MACRO cbx_1__2_
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  SIZE 75.44 BY 76.16 ;
  SYMMETRY X Y ;
  PIN pReset[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 47.11 0.8 47.41 ;
    END
  END pReset[0]
  PIN chanx_left_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 36.23 0.8 36.53 ;
    END
  END chanx_left_in[0]
  PIN chanx_left_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 34.1 0.595 34.24 ;
    END
  END chanx_left_in[1]
  PIN chanx_left_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 36.82 0.595 36.96 ;
    END
  END chanx_left_in[2]
  PIN chanx_left_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 37.59 0.8 37.89 ;
    END
  END chanx_left_in[3]
  PIN chanx_left_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 13.11 0.8 13.41 ;
    END
  END chanx_left_in[4]
  PIN chanx_left_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 28.07 0.8 28.37 ;
    END
  END chanx_left_in[5]
  PIN chanx_left_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 14.47 0.8 14.77 ;
    END
  END chanx_left_in[6]
  PIN chanx_left_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 5.63 0.8 5.93 ;
    END
  END chanx_left_in[7]
  PIN chanx_left_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 19.82 0.595 19.96 ;
    END
  END chanx_left_in[8]
  PIN chanx_left_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 27.98 0.595 28.12 ;
    END
  END chanx_left_in[9]
  PIN chanx_left_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 15.83 0.8 16.13 ;
    END
  END chanx_left_in[10]
  PIN chanx_left_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 15.06 0.595 15.2 ;
    END
  END chanx_left_in[11]
  PIN chanx_left_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 18.12 0.595 18.26 ;
    END
  END chanx_left_in[12]
  PIN chanx_left_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 11.75 0.8 12.05 ;
    END
  END chanx_left_in[13]
  PIN chanx_left_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 30.79 0.8 31.09 ;
    END
  END chanx_left_in[14]
  PIN chanx_left_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 29.43 0.8 29.73 ;
    END
  END chanx_left_in[15]
  PIN chanx_left_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 6.99 0.8 7.29 ;
    END
  END chanx_left_in[16]
  PIN chanx_left_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 17.44 0.595 17.58 ;
    END
  END chanx_left_in[17]
  PIN chanx_left_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 33.51 0.8 33.81 ;
    END
  END chanx_left_in[18]
  PIN chanx_left_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 9.71 0.8 10.01 ;
    END
  END chanx_left_in[19]
  PIN chanx_left_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 17.19 0.8 17.49 ;
    END
  END chanx_left_in[20]
  PIN chanx_left_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 26.71 0.8 27.01 ;
    END
  END chanx_left_in[21]
  PIN chanx_left_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 33.42 0.595 33.56 ;
    END
  END chanx_left_in[22]
  PIN chanx_left_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 19.91 0.8 20.21 ;
    END
  END chanx_left_in[23]
  PIN chanx_left_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 40.31 0.8 40.61 ;
    END
  END chanx_left_in[24]
  PIN chanx_left_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 38.95 0.8 39.25 ;
    END
  END chanx_left_in[25]
  PIN chanx_left_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 47.7 0.595 47.84 ;
    END
  END chanx_left_in[26]
  PIN chanx_left_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 44.3 0.595 44.44 ;
    END
  END chanx_left_in[27]
  PIN chanx_left_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 8.35 0.8 8.65 ;
    END
  END chanx_left_in[28]
  PIN chanx_left_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 18.55 0.8 18.85 ;
    END
  END chanx_left_in[29]
  PIN chanx_right_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 74.845 42.6 75.44 42.74 ;
    END
  END chanx_right_in[0]
  PIN chanx_right_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 74.845 37.16 75.44 37.3 ;
    END
  END chanx_right_in[1]
  PIN chanx_right_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 74.845 45.32 75.44 45.46 ;
    END
  END chanx_right_in[2]
  PIN chanx_right_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 74.64 36.91 75.44 37.21 ;
    END
  END chanx_right_in[3]
  PIN chanx_right_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 74.64 39.63 75.44 39.93 ;
    END
  END chanx_right_in[4]
  PIN chanx_right_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 74.64 38.27 75.44 38.57 ;
    END
  END chanx_right_in[5]
  PIN chanx_right_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 74.64 26.03 75.44 26.33 ;
    END
  END chanx_right_in[6]
  PIN chanx_right_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 74.845 7.24 75.44 7.38 ;
    END
  END chanx_right_in[7]
  PIN chanx_right_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 74.64 19.23 75.44 19.53 ;
    END
  END chanx_right_in[8]
  PIN chanx_right_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 74.64 17.87 75.44 18.17 ;
    END
  END chanx_right_in[9]
  PIN chanx_right_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 74.64 27.39 75.44 27.69 ;
    END
  END chanx_right_in[10]
  PIN chanx_right_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 74.64 21.95 75.44 22.25 ;
    END
  END chanx_right_in[11]
  PIN chanx_right_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 74.845 14.72 75.44 14.86 ;
    END
  END chanx_right_in[12]
  PIN chanx_right_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 74.845 4.52 75.44 4.66 ;
    END
  END chanx_right_in[13]
  PIN chanx_right_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 74.64 35.55 75.44 35.85 ;
    END
  END chanx_right_in[14]
  PIN chanx_right_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 74.64 34.19 75.44 34.49 ;
    END
  END chanx_right_in[15]
  PIN chanx_right_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 74.845 3.84 75.44 3.98 ;
    END
  END chanx_right_in[16]
  PIN chanx_right_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 74.845 15.4 75.44 15.54 ;
    END
  END chanx_right_in[17]
  PIN chanx_right_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 74.845 53.14 75.44 53.28 ;
    END
  END chanx_right_in[18]
  PIN chanx_right_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 74.64 7.67 75.44 7.97 ;
    END
  END chanx_right_in[19]
  PIN chanx_right_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 74.845 30.7 75.44 30.84 ;
    END
  END chanx_right_in[20]
  PIN chanx_right_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 74.845 28.66 75.44 28.8 ;
    END
  END chanx_right_in[21]
  PIN chanx_right_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 74.64 12.43 75.44 12.73 ;
    END
  END chanx_right_in[22]
  PIN chanx_right_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 74.845 20.16 75.44 20.3 ;
    END
  END chanx_right_in[23]
  PIN chanx_right_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 74.64 31.47 75.44 31.77 ;
    END
  END chanx_right_in[24]
  PIN chanx_right_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 74.845 34.1 75.44 34.24 ;
    END
  END chanx_right_in[25]
  PIN chanx_right_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 74.64 28.75 75.44 29.05 ;
    END
  END chanx_right_in[26]
  PIN chanx_right_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 74.845 38.86 75.44 39 ;
    END
  END chanx_right_in[27]
  PIN chanx_right_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 74.64 6.31 75.44 6.61 ;
    END
  END chanx_right_in[28]
  PIN chanx_right_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 74.845 18.12 75.44 18.26 ;
    END
  END chanx_right_in[29]
  PIN ccff_head[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 74.64 11.07 75.44 11.37 ;
    END
  END ccff_head[0]
  PIN chanx_left_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 32.15 0.8 32.45 ;
    END
  END chanx_left_out[0]
  PIN chanx_left_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 66.4 0.595 66.54 ;
    END
  END chanx_left_out[1]
  PIN chanx_left_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 50.42 0.595 50.56 ;
    END
  END chanx_left_out[2]
  PIN chanx_left_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 39.54 0.595 39.68 ;
    END
  END chanx_left_out[3]
  PIN chanx_left_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 44.39 0.8 44.69 ;
    END
  END chanx_left_out[4]
  PIN chanx_left_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 42.6 0.595 42.74 ;
    END
  END chanx_left_out[5]
  PIN chanx_left_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 45.75 0.8 46.05 ;
    END
  END chanx_left_out[6]
  PIN chanx_left_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 7.24 0.595 7.38 ;
    END
  END chanx_left_out[7]
  PIN chanx_left_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 25.35 0.8 25.65 ;
    END
  END chanx_left_out[8]
  PIN chanx_left_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 41.58 0.595 41.72 ;
    END
  END chanx_left_out[9]
  PIN chanx_left_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 21.27 0.8 21.57 ;
    END
  END chanx_left_out[10]
  PIN chanx_left_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 23.99 0.8 24.29 ;
    END
  END chanx_left_out[11]
  PIN chanx_left_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 25.26 0.595 25.4 ;
    END
  END chanx_left_out[12]
  PIN chanx_left_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 38.86 0.595 39 ;
    END
  END chanx_left_out[13]
  PIN chanx_left_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 49.74 0.595 49.88 ;
    END
  END chanx_left_out[14]
  PIN chanx_left_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 22.63 0.8 22.93 ;
    END
  END chanx_left_out[15]
  PIN chanx_left_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 43.03 0.8 43.33 ;
    END
  END chanx_left_out[16]
  PIN chanx_left_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 12.68 0.595 12.82 ;
    END
  END chanx_left_out[17]
  PIN chanx_left_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 20.84 0.595 20.98 ;
    END
  END chanx_left_out[18]
  PIN chanx_left_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 44.98 0.595 45.12 ;
    END
  END chanx_left_out[19]
  PIN chanx_left_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 57.9 0.595 58.04 ;
    END
  END chanx_left_out[20]
  PIN chanx_left_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 26.28 0.595 26.42 ;
    END
  END chanx_left_out[21]
  PIN chanx_left_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 41.67 0.8 41.97 ;
    END
  END chanx_left_out[22]
  PIN chanx_left_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 22.88 0.595 23.02 ;
    END
  END chanx_left_out[23]
  PIN chanx_left_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 47.02 0.595 47.16 ;
    END
  END chanx_left_out[24]
  PIN chanx_left_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 34.87 0.8 35.17 ;
    END
  END chanx_left_out[25]
  PIN chanx_left_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 23.56 0.595 23.7 ;
    END
  END chanx_left_out[26]
  PIN chanx_left_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 60.62 0.595 60.76 ;
    END
  END chanx_left_out[27]
  PIN chanx_left_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 30.7 0.595 30.84 ;
    END
  END chanx_left_out[28]
  PIN chanx_left_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 58.58 0.595 58.72 ;
    END
  END chanx_left_out[29]
  PIN chanx_right_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 74.845 27.98 75.44 28.12 ;
    END
  END chanx_right_out[0]
  PIN chanx_right_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 74.64 13.79 75.44 14.09 ;
    END
  END chanx_right_out[1]
  PIN chanx_right_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 74.64 32.83 75.44 33.13 ;
    END
  END chanx_right_out[2]
  PIN chanx_right_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 74.845 9.96 75.44 10.1 ;
    END
  END chanx_right_out[3]
  PIN chanx_right_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 74.64 16.51 75.44 16.81 ;
    END
  END chanx_right_out[4]
  PIN chanx_right_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 74.845 12.68 75.44 12.82 ;
    END
  END chanx_right_out[5]
  PIN chanx_right_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 74.845 23.56 75.44 23.7 ;
    END
  END chanx_right_out[6]
  PIN chanx_right_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 74.64 15.15 75.44 15.45 ;
    END
  END chanx_right_out[7]
  PIN chanx_right_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 74.845 12 75.44 12.14 ;
    END
  END chanx_right_out[8]
  PIN chanx_right_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 74.845 52.46 75.44 52.6 ;
    END
  END chanx_right_out[9]
  PIN chanx_right_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 74.845 47.02 75.44 47.16 ;
    END
  END chanx_right_out[10]
  PIN chanx_right_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 74.845 33.42 75.44 33.56 ;
    END
  END chanx_right_out[11]
  PIN chanx_right_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 74.64 24.67 75.44 24.97 ;
    END
  END chanx_right_out[12]
  PIN chanx_right_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 74.845 31.38 75.44 31.52 ;
    END
  END chanx_right_out[13]
  PIN chanx_right_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 74.845 44.3 75.44 44.44 ;
    END
  END chanx_right_out[14]
  PIN chanx_right_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 74.845 39.54 75.44 39.68 ;
    END
  END chanx_right_out[15]
  PIN chanx_right_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 74.845 50.42 75.44 50.56 ;
    END
  END chanx_right_out[16]
  PIN chanx_right_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 74.845 20.84 75.44 20.98 ;
    END
  END chanx_right_out[17]
  PIN chanx_right_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 74.845 36.14 75.44 36.28 ;
    END
  END chanx_right_out[18]
  PIN chanx_right_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 74.64 20.59 75.44 20.89 ;
    END
  END chanx_right_out[19]
  PIN chanx_right_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 74.64 30.11 75.44 30.41 ;
    END
  END chanx_right_out[20]
  PIN chanx_right_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 74.64 23.31 75.44 23.61 ;
    END
  END chanx_right_out[21]
  PIN chanx_right_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 74.845 17.44 75.44 17.58 ;
    END
  END chanx_right_out[22]
  PIN chanx_right_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 74.845 25.94 75.44 26.08 ;
    END
  END chanx_right_out[23]
  PIN chanx_right_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 74.845 22.88 75.44 23.02 ;
    END
  END chanx_right_out[24]
  PIN chanx_right_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 74.845 41.58 75.44 41.72 ;
    END
  END chanx_right_out[25]
  PIN chanx_right_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 74.845 47.7 75.44 47.84 ;
    END
  END chanx_right_out[26]
  PIN chanx_right_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 74.845 49.74 75.44 49.88 ;
    END
  END chanx_right_out[27]
  PIN chanx_right_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 74.64 42.35 75.44 42.65 ;
    END
  END chanx_right_out[28]
  PIN chanx_right_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 74.845 25.26 75.44 25.4 ;
    END
  END chanx_right_out[29]
  PIN top_grid_pin_0_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.8 0 38.94 0.485 ;
    END
  END top_grid_pin_0_[0]
  PIN bottom_grid_pin_0_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.38 0 3.52 0.485 ;
    END
  END bottom_grid_pin_0_[0]
  PIN bottom_grid_pin_1_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 1.8 0.595 1.94 ;
    END
  END bottom_grid_pin_1_[0]
  PIN bottom_grid_pin_2_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.46 0 2.6 0.485 ;
    END
  END bottom_grid_pin_2_[0]
  PIN bottom_grid_pin_3_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.3 0 4.44 0.485 ;
    END
  END bottom_grid_pin_3_[0]
  PIN bottom_grid_pin_4_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.34 0 15.48 0.485 ;
    END
  END bottom_grid_pin_4_[0]
  PIN bottom_grid_pin_5_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.06 0 30.2 0.485 ;
    END
  END bottom_grid_pin_5_[0]
  PIN bottom_grid_pin_6_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.76 0 27.9 0.485 ;
    END
  END bottom_grid_pin_6_[0]
  PIN bottom_grid_pin_7_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.96 0 37.1 0.485 ;
    END
  END bottom_grid_pin_7_[0]
  PIN bottom_grid_pin_8_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.9 0 9.04 0.485 ;
    END
  END bottom_grid_pin_8_[0]
  PIN bottom_grid_pin_9_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.98 0 8.12 0.485 ;
    END
  END bottom_grid_pin_9_[0]
  PIN bottom_grid_pin_10_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.22 0 5.36 0.485 ;
    END
  END bottom_grid_pin_10_[0]
  PIN bottom_grid_pin_11_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.14 0 6.28 0.485 ;
    END
  END bottom_grid_pin_11_[0]
  PIN bottom_grid_pin_12_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.24 0 22.38 0.485 ;
    END
  END bottom_grid_pin_12_[0]
  PIN bottom_grid_pin_13_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.42 0 14.56 0.485 ;
    END
  END bottom_grid_pin_13_[0]
  PIN bottom_grid_pin_14_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.36 0 32.5 0.485 ;
    END
  END bottom_grid_pin_14_[0]
  PIN bottom_grid_pin_15_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.26 0 16.4 0.485 ;
    END
  END bottom_grid_pin_15_[0]
  PIN ccff_tail[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 6.56 0.595 6.7 ;
    END
  END ccff_tail[0]
  PIN IO_ISOL_N[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 3.5 0.595 3.64 ;
    END
  END IO_ISOL_N[0]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.06 75.675 7.2 76.16 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[0]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.68 75.675 5.82 76.16 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[0]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.92 75.675 3.06 76.16 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[0]
  PIN bottom_width_0_height_0__pin_0_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.88 0 38.02 0.485 ;
    END
  END bottom_width_0_height_0__pin_0_[0]
  PIN bottom_width_0_height_0__pin_1_upper[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 31.38 0.595 31.52 ;
    END
  END bottom_width_0_height_0__pin_1_upper[0]
  PIN bottom_width_0_height_0__pin_1_lower[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 74.64 40.99 75.44 41.29 ;
    END
  END bottom_width_0_height_0__pin_1_lower[0]
  PIN SC_IN_TOP
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 11.66 0.595 11.8 ;
    END
  END SC_IN_TOP
  PIN SC_OUT_BOT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.92 0 26.06 0.485 ;
    END
  END SC_OUT_BOT
  PIN SC_IN_BOT
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.56 0 64.7 0.485 ;
    END
  END SC_IN_BOT
  PIN SC_OUT_TOP
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 74.64 9.03 75.44 9.33 ;
    END
  END SC_OUT_TOP
  PIN pReset_E_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 74.64 4.27 75.44 4.57 ;
    END
  END pReset_E_in
  PIN pReset_W_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 36.14 0.595 36.28 ;
    END
  END pReset_W_in
  PIN pReset_W_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 29 0.595 29.14 ;
    END
  END pReset_W_out
  PIN pReset_S_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.72 0 62.86 0.485 ;
    END
  END pReset_S_out
  PIN pReset_E_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 74.845 6.56 75.44 6.7 ;
    END
  END pReset_E_out
  PIN prog_clk_0_S_in
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER met2 ;
        RECT 26.84 0 26.98 0.485 ;
    END
  END prog_clk_0_S_in
  PIN prog_clk_0_W_out
    DIRECTION OUTPUT ;
    USE CLOCK ;
    PORT
      LAYER met1 ;
        RECT 0 14.38 0.595 14.52 ;
    END
  END prog_clk_0_W_out
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0 16.08 3.2 19.28 ;
        RECT 72.24 16.08 75.44 19.28 ;
        RECT 0 56.88 3.2 60.08 ;
        RECT 72.24 56.88 75.44 60.08 ;
      LAYER met4 ;
        RECT 7.98 0 8.58 0.6 ;
        RECT 37.42 0 38.02 0.6 ;
        RECT 66.86 0 67.46 0.6 ;
        RECT 7.98 75.56 8.58 76.16 ;
        RECT 37.42 75.56 38.02 76.16 ;
        RECT 66.86 75.56 67.46 76.16 ;
      LAYER met1 ;
        RECT 0 2.48 0.48 2.96 ;
        RECT 74.96 2.48 75.44 2.96 ;
        RECT 0 7.92 0.48 8.4 ;
        RECT 74.96 7.92 75.44 8.4 ;
        RECT 0 13.36 0.48 13.84 ;
        RECT 74.96 13.36 75.44 13.84 ;
        RECT 0 18.8 0.48 19.28 ;
        RECT 74.96 18.8 75.44 19.28 ;
        RECT 0 24.24 0.48 24.72 ;
        RECT 74.96 24.24 75.44 24.72 ;
        RECT 0 29.68 0.48 30.16 ;
        RECT 74.96 29.68 75.44 30.16 ;
        RECT 0 35.12 0.48 35.6 ;
        RECT 74.96 35.12 75.44 35.6 ;
        RECT 0 40.56 0.48 41.04 ;
        RECT 74.96 40.56 75.44 41.04 ;
        RECT 0 46 0.48 46.48 ;
        RECT 74.96 46 75.44 46.48 ;
        RECT 0 51.44 0.48 51.92 ;
        RECT 74.96 51.44 75.44 51.92 ;
        RECT 0 56.88 0.48 57.36 ;
        RECT 74.96 56.88 75.44 57.36 ;
        RECT 0 62.32 0.48 62.8 ;
        RECT 74.96 62.32 75.44 62.8 ;
        RECT 0 67.76 0.48 68.24 ;
        RECT 74.96 67.76 75.44 68.24 ;
        RECT 0 73.2 0.48 73.68 ;
        RECT 74.96 73.2 75.44 73.68 ;
    END
  END VDD
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0 36.48 3.2 39.68 ;
        RECT 72.24 36.48 75.44 39.68 ;
      LAYER met4 ;
        RECT 22.7 0 23.3 0.6 ;
        RECT 52.14 0 52.74 0.6 ;
        RECT 22.7 75.56 23.3 76.16 ;
        RECT 52.14 75.56 52.74 76.16 ;
      LAYER met1 ;
        RECT 0 -0.24 0.48 0.24 ;
        RECT 74.96 -0.24 75.44 0.24 ;
        RECT 0 5.2 0.48 5.68 ;
        RECT 74.96 5.2 75.44 5.68 ;
        RECT 0 10.64 0.48 11.12 ;
        RECT 74.96 10.64 75.44 11.12 ;
        RECT 0 16.08 0.48 16.56 ;
        RECT 74.96 16.08 75.44 16.56 ;
        RECT 0 21.52 0.48 22 ;
        RECT 74.96 21.52 75.44 22 ;
        RECT 0 26.96 0.48 27.44 ;
        RECT 74.96 26.96 75.44 27.44 ;
        RECT 0 32.4 0.48 32.88 ;
        RECT 74.96 32.4 75.44 32.88 ;
        RECT 0 37.84 0.48 38.32 ;
        RECT 74.96 37.84 75.44 38.32 ;
        RECT 0 43.28 0.48 43.76 ;
        RECT 74.96 43.28 75.44 43.76 ;
        RECT 0 48.72 0.48 49.2 ;
        RECT 74.96 48.72 75.44 49.2 ;
        RECT 0 54.16 0.48 54.64 ;
        RECT 74.96 54.16 75.44 54.64 ;
        RECT 0 59.6 0.48 60.08 ;
        RECT 74.96 59.6 75.44 60.08 ;
        RECT 0 65.04 0.48 65.52 ;
        RECT 74.96 65.04 75.44 65.52 ;
        RECT 0 70.48 0.48 70.96 ;
        RECT 74.96 70.48 75.44 70.96 ;
        RECT 0 75.92 0.48 76.4 ;
        RECT 74.96 75.92 75.44 76.4 ;
    END
  END VSS
  OBS
    LAYER met3 ;
      POLYGON 52.605 76.205 52.605 76.2 52.82 76.2 52.82 75.88 52.605 75.88 52.605 75.875 52.275 75.875 52.275 75.88 52.06 75.88 52.06 76.2 52.275 76.2 52.275 76.205 ;
      POLYGON 23.165 76.205 23.165 76.2 23.38 76.2 23.38 75.88 23.165 75.88 23.165 75.875 22.835 75.875 22.835 75.88 22.62 75.88 22.62 76.2 22.835 76.2 22.835 76.205 ;
      POLYGON 4.98 41.29 4.98 40.99 0.65 40.99 0.65 41.27 1.2 41.27 1.2 41.29 ;
      POLYGON 1.76 14.09 1.76 13.79 1.2 13.79 1.2 13.81 0 13.81 0 14.09 ;
      POLYGON 52.605 0.285 52.605 0.28 52.82 0.28 52.82 -0.04 52.605 -0.04 52.605 -0.045 52.275 -0.045 52.275 -0.04 52.06 -0.04 52.06 0.28 52.275 0.28 52.275 0.285 ;
      POLYGON 23.165 0.285 23.165 0.28 23.38 0.28 23.38 -0.04 23.165 -0.04 23.165 -0.045 22.835 -0.045 22.835 -0.04 22.62 -0.04 22.62 0.28 22.835 0.28 22.835 0.285 ;
      POLYGON 75.04 75.76 75.04 43.05 74.24 43.05 74.24 41.95 75.04 41.95 75.04 41.69 74.24 41.69 74.24 40.59 75.04 40.59 75.04 40.33 74.24 40.33 74.24 39.23 75.04 39.23 75.04 38.97 74.24 38.97 74.24 37.87 75.04 37.87 75.04 37.61 74.24 37.61 74.24 36.51 75.04 36.51 75.04 36.25 74.24 36.25 74.24 35.15 75.04 35.15 75.04 34.89 74.24 34.89 74.24 33.79 75.04 33.79 75.04 33.53 74.24 33.53 74.24 32.43 75.04 32.43 75.04 32.17 74.24 32.17 74.24 31.07 75.04 31.07 75.04 30.81 74.24 30.81 74.24 29.71 75.04 29.71 75.04 29.45 74.24 29.45 74.24 28.35 75.04 28.35 75.04 28.09 74.24 28.09 74.24 26.99 75.04 26.99 75.04 26.73 74.24 26.73 74.24 25.63 75.04 25.63 75.04 25.37 74.24 25.37 74.24 24.27 75.04 24.27 75.04 24.01 74.24 24.01 74.24 22.91 75.04 22.91 75.04 22.65 74.24 22.65 74.24 21.55 75.04 21.55 75.04 21.29 74.24 21.29 74.24 20.19 75.04 20.19 75.04 19.93 74.24 19.93 74.24 18.83 75.04 18.83 75.04 18.57 74.24 18.57 74.24 17.47 75.04 17.47 75.04 17.21 74.24 17.21 74.24 16.11 75.04 16.11 75.04 15.85 74.24 15.85 74.24 14.75 75.04 14.75 75.04 14.49 74.24 14.49 74.24 13.39 75.04 13.39 75.04 13.13 74.24 13.13 74.24 12.03 75.04 12.03 75.04 11.77 74.24 11.77 74.24 10.67 75.04 10.67 75.04 9.73 74.24 9.73 74.24 8.63 75.04 8.63 75.04 8.37 74.24 8.37 74.24 7.27 75.04 7.27 75.04 7.01 74.24 7.01 74.24 5.91 75.04 5.91 75.04 4.97 74.24 4.97 74.24 3.87 75.04 3.87 75.04 0.4 0.4 0.4 0.4 5.23 1.2 5.23 1.2 6.33 0.4 6.33 0.4 6.59 1.2 6.59 1.2 7.69 0.4 7.69 0.4 7.95 1.2 7.95 1.2 9.05 0.4 9.05 0.4 9.31 1.2 9.31 1.2 10.41 0.4 10.41 0.4 11.35 1.2 11.35 1.2 12.45 0.4 12.45 0.4 12.71 1.2 12.71 1.2 13.81 0.4 13.81 0.4 14.07 1.2 14.07 1.2 15.17 0.4 15.17 0.4 15.43 1.2 15.43 1.2 16.53 0.4 16.53 0.4 16.79 1.2 16.79 1.2 17.89 0.4 17.89 0.4 18.15 1.2 18.15 1.2 19.25 0.4 19.25 0.4 19.51 1.2 19.51 1.2 20.61 0.4 20.61 0.4 20.87 1.2 20.87 1.2 21.97 0.4 21.97 0.4 22.23 1.2 22.23 1.2 23.33 0.4 23.33 0.4 23.59 1.2 23.59 1.2 24.69 0.4 24.69 0.4 24.95 1.2 24.95 1.2 26.05 0.4 26.05 0.4 26.31 1.2 26.31 1.2 27.41 0.4 27.41 0.4 27.67 1.2 27.67 1.2 28.77 0.4 28.77 0.4 29.03 1.2 29.03 1.2 30.13 0.4 30.13 0.4 30.39 1.2 30.39 1.2 31.49 0.4 31.49 0.4 31.75 1.2 31.75 1.2 32.85 0.4 32.85 0.4 33.11 1.2 33.11 1.2 34.21 0.4 34.21 0.4 34.47 1.2 34.47 1.2 35.57 0.4 35.57 0.4 35.83 1.2 35.83 1.2 36.93 0.4 36.93 0.4 37.19 1.2 37.19 1.2 38.29 0.4 38.29 0.4 38.55 1.2 38.55 1.2 39.65 0.4 39.65 0.4 39.91 1.2 39.91 1.2 41.01 0.4 41.01 0.4 41.27 1.2 41.27 1.2 42.37 0.4 42.37 0.4 42.63 1.2 42.63 1.2 43.73 0.4 43.73 0.4 43.99 1.2 43.99 1.2 45.09 0.4 45.09 0.4 45.35 1.2 45.35 1.2 46.45 0.4 46.45 0.4 46.71 1.2 46.71 1.2 47.81 0.4 47.81 0.4 75.76 ;
    LAYER met1 ;
      POLYGON 74.68 76.4 74.68 75.92 52.6 75.92 52.6 75.91 52.28 75.91 52.28 75.92 23.16 75.92 23.16 75.91 22.84 75.91 22.84 75.92 0.76 75.92 0.76 76.4 ;
      POLYGON 74.82 32.2 74.82 31.8 74.68 31.8 74.68 32.06 68.24 32.06 68.24 32.2 ;
      POLYGON 1.68 11.46 1.68 11.32 0.525 11.32 0.525 11.38 0.875 11.38 0.875 11.46 ;
      POLYGON 52.6 0.25 52.6 0.24 74.68 0.24 74.68 -0.24 0.76 -0.24 0.76 0.24 22.84 0.24 22.84 0.25 23.16 0.25 23.16 0.24 52.28 0.24 52.28 0.25 ;
      POLYGON 74.68 75.88 74.68 75.64 75.16 75.64 75.16 73.96 74.68 73.96 74.68 72.92 75.16 72.92 75.16 71.24 74.68 71.24 74.68 70.2 75.16 70.2 75.16 68.52 74.68 68.52 74.68 67.48 75.16 67.48 75.16 65.8 74.68 65.8 74.68 64.76 75.16 64.76 75.16 63.08 74.68 63.08 74.68 62.04 75.16 62.04 75.16 60.36 74.68 60.36 74.68 59.32 75.16 59.32 75.16 57.64 74.68 57.64 74.68 56.6 75.16 56.6 75.16 54.92 74.68 54.92 74.68 53.88 75.16 53.88 75.16 53.56 74.565 53.56 74.565 52.18 74.68 52.18 74.68 51.16 75.16 51.16 75.16 50.84 74.565 50.84 74.565 49.46 74.68 49.46 74.68 48.44 75.16 48.44 75.16 48.12 74.565 48.12 74.565 46.74 74.68 46.74 74.68 45.74 74.565 45.74 74.565 45.04 75.16 45.04 75.16 44.72 74.565 44.72 74.565 44.02 74.68 44.02 74.68 43.02 74.565 43.02 74.565 42.32 75.16 42.32 75.16 42 74.565 42 74.565 41.3 74.68 41.3 74.68 40.28 75.16 40.28 75.16 39.96 74.565 39.96 74.565 38.58 74.68 38.58 74.68 37.58 74.565 37.58 74.565 36.88 75.16 36.88 75.16 36.56 74.565 36.56 74.565 35.86 74.68 35.86 74.68 34.84 75.16 34.84 75.16 34.52 74.565 34.52 74.565 33.14 74.68 33.14 74.68 32.12 75.16 32.12 75.16 31.8 74.565 31.8 74.565 30.42 74.68 30.42 74.68 29.4 75.16 29.4 75.16 29.08 74.565 29.08 74.565 27.7 74.68 27.7 74.68 26.68 75.16 26.68 75.16 26.36 74.565 26.36 74.565 24.98 74.68 24.98 74.68 23.98 74.565 23.98 74.565 22.6 75.16 22.6 75.16 22.28 74.68 22.28 74.68 21.26 74.565 21.26 74.565 19.88 75.16 19.88 75.16 19.56 74.68 19.56 74.68 18.54 74.565 18.54 74.565 17.16 75.16 17.16 75.16 16.84 74.68 16.84 74.68 15.82 74.565 15.82 74.565 14.44 75.16 14.44 75.16 14.12 74.68 14.12 74.68 13.1 74.565 13.1 74.565 11.72 75.16 11.72 75.16 11.4 74.68 11.4 74.68 10.38 74.565 10.38 74.565 9.68 75.16 9.68 75.16 8.68 74.68 8.68 74.68 7.66 74.565 7.66 74.565 6.28 75.16 6.28 75.16 5.96 74.68 5.96 74.68 4.94 74.565 4.94 74.565 3.56 75.16 3.56 75.16 3.24 74.68 3.24 74.68 2.2 75.16 2.2 75.16 0.52 74.68 0.52 74.68 0.28 0.76 0.28 0.76 0.52 0.28 0.52 0.28 1.52 0.875 1.52 0.875 2.22 0.76 2.22 0.76 3.22 0.875 3.22 0.875 3.92 0.28 3.92 0.28 4.92 0.76 4.92 0.76 5.96 0.28 5.96 0.28 6.28 0.875 6.28 0.875 7.66 0.76 7.66 0.76 8.68 0.28 8.68 0.28 10.36 0.76 10.36 0.76 11.38 0.875 11.38 0.875 12.08 0.28 12.08 0.28 12.4 0.875 12.4 0.875 13.1 0.76 13.1 0.76 14.1 0.875 14.1 0.875 15.48 0.28 15.48 0.28 15.8 0.76 15.8 0.76 16.84 0.28 16.84 0.28 17.16 0.875 17.16 0.875 18.54 0.76 18.54 0.76 19.54 0.875 19.54 0.875 20.24 0.28 20.24 0.28 20.56 0.875 20.56 0.875 21.26 0.76 21.26 0.76 22.28 0.28 22.28 0.28 22.6 0.875 22.6 0.875 23.98 0.76 23.98 0.76 24.98 0.875 24.98 0.875 25.68 0.28 25.68 0.28 26 0.875 26 0.875 26.7 0.76 26.7 0.76 27.7 0.875 27.7 0.875 28.4 0.28 28.4 0.28 28.72 0.875 28.72 0.875 29.42 0.76 29.42 0.76 30.42 0.875 30.42 0.875 31.8 0.28 31.8 0.28 32.12 0.76 32.12 0.76 33.14 0.875 33.14 0.875 34.52 0.28 34.52 0.28 34.84 0.76 34.84 0.76 35.86 0.875 35.86 0.875 37.24 0.28 37.24 0.28 37.56 0.76 37.56 0.76 38.58 0.875 38.58 0.875 39.96 0.28 39.96 0.28 40.28 0.76 40.28 0.76 41.3 0.875 41.3 0.875 42 0.28 42 0.28 42.32 0.875 42.32 0.875 43.02 0.76 43.02 0.76 44.02 0.875 44.02 0.875 45.4 0.28 45.4 0.28 45.72 0.76 45.72 0.76 46.74 0.875 46.74 0.875 48.12 0.28 48.12 0.28 48.44 0.76 48.44 0.76 49.46 0.875 49.46 0.875 50.84 0.28 50.84 0.28 51.16 0.76 51.16 0.76 52.2 0.28 52.2 0.28 53.88 0.76 53.88 0.76 54.92 0.28 54.92 0.28 56.6 0.76 56.6 0.76 57.62 0.875 57.62 0.875 59 0.28 59 0.28 59.32 0.76 59.32 0.76 60.34 0.875 60.34 0.875 61.04 0.28 61.04 0.28 62.04 0.76 62.04 0.76 63.08 0.28 63.08 0.28 64.76 0.76 64.76 0.76 65.8 0.28 65.8 0.28 66.12 0.875 66.12 0.875 66.82 0.28 66.82 0.28 67.48 0.76 67.48 0.76 68.52 0.28 68.52 0.28 70.2 0.76 70.2 0.76 71.24 0.28 71.24 0.28 72.92 0.76 72.92 0.76 73.96 0.28 73.96 0.28 75.64 0.76 75.64 0.76 75.88 ;
    LAYER met2 ;
      RECT 52.3 75.855 52.58 76.225 ;
      RECT 22.86 75.855 23.14 76.225 ;
      RECT 4.7 0.69 4.96 1.01 ;
      RECT 52.3 -0.065 52.58 0.305 ;
      RECT 22.86 -0.065 23.14 0.305 ;
      POLYGON 75.16 75.88 75.16 0.28 64.98 0.28 64.98 0.765 64.28 0.765 64.28 0.28 63.14 0.28 63.14 0.765 62.44 0.765 62.44 0.28 39.22 0.28 39.22 0.765 38.52 0.765 38.52 0.28 38.3 0.28 38.3 0.765 37.6 0.765 37.6 0.28 37.38 0.28 37.38 0.765 36.68 0.765 36.68 0.28 32.78 0.28 32.78 0.765 32.08 0.765 32.08 0.28 30.48 0.28 30.48 0.765 29.78 0.765 29.78 0.28 28.18 0.28 28.18 0.765 27.48 0.765 27.48 0.28 27.26 0.28 27.26 0.765 26.56 0.765 26.56 0.28 26.34 0.28 26.34 0.765 25.64 0.765 25.64 0.28 22.66 0.28 22.66 0.765 21.96 0.765 21.96 0.28 16.68 0.28 16.68 0.765 15.98 0.765 15.98 0.28 15.76 0.28 15.76 0.765 15.06 0.765 15.06 0.28 14.84 0.28 14.84 0.765 14.14 0.765 14.14 0.28 9.32 0.28 9.32 0.765 8.62 0.765 8.62 0.28 8.4 0.28 8.4 0.765 7.7 0.765 7.7 0.28 6.56 0.28 6.56 0.765 5.86 0.765 5.86 0.28 5.64 0.28 5.64 0.765 4.94 0.765 4.94 0.28 4.72 0.28 4.72 0.765 4.02 0.765 4.02 0.28 3.8 0.28 3.8 0.765 3.1 0.765 3.1 0.28 2.88 0.28 2.88 0.765 2.18 0.765 2.18 0.28 0.28 0.28 0.28 75.88 2.64 75.88 2.64 75.395 3.34 75.395 3.34 75.88 5.4 75.88 5.4 75.395 6.1 75.395 6.1 75.88 6.78 75.88 6.78 75.395 7.48 75.395 7.48 75.88 ;
    LAYER met4 ;
      POLYGON 75.04 75.76 75.04 0.4 67.86 0.4 67.86 1 66.46 1 66.46 0.4 53.14 0.4 53.14 1 51.74 1 51.74 0.4 38.42 0.4 38.42 1 37.02 1 37.02 0.4 23.7 0.4 23.7 1 22.3 1 22.3 0.4 8.98 0.4 8.98 1 7.58 1 7.58 0.4 0.4 0.4 0.4 75.76 7.58 75.76 7.58 75.16 8.98 75.16 8.98 75.76 22.3 75.76 22.3 75.16 23.7 75.16 23.7 75.76 37.02 75.76 37.02 75.16 38.42 75.16 38.42 75.76 51.74 75.76 51.74 75.16 53.14 75.16 53.14 75.76 66.46 75.76 66.46 75.16 67.86 75.16 67.86 75.76 ;
    LAYER met5 ;
      POLYGON 73.84 74.56 73.84 61.68 70.64 61.68 70.64 55.28 73.84 55.28 73.84 41.28 70.64 41.28 70.64 34.88 73.84 34.88 73.84 20.88 70.64 20.88 70.64 14.48 73.84 14.48 73.84 1.6 1.6 1.6 1.6 14.48 4.8 14.48 4.8 20.88 1.6 20.88 1.6 34.88 4.8 34.88 4.8 41.28 1.6 41.28 1.6 55.28 4.8 55.28 4.8 61.68 1.6 61.68 1.6 74.56 ;
    LAYER li1 ;
      POLYGON 75.44 76.245 75.44 76.075 71.855 76.075 71.855 75.54 71.345 75.54 71.345 76.075 69.385 76.075 69.385 75.675 69.055 75.675 69.055 76.075 68.025 76.075 68.025 75.615 67.72 75.615 67.72 76.075 66.235 76.075 66.235 75.635 66.045 75.635 66.045 76.075 64.145 76.075 64.145 75.615 63.815 75.615 63.815 76.075 61.215 76.075 61.215 75.715 60.885 75.715 60.885 76.075 60.185 76.075 60.185 75.695 59.855 75.695 59.855 76.075 58.825 76.075 58.825 75.615 58.52 75.615 58.52 76.075 57.035 76.075 57.035 75.635 56.845 75.635 56.845 76.075 54.945 76.075 54.945 75.615 54.615 75.615 54.615 76.075 52.015 76.075 52.015 75.715 51.685 75.715 51.685 76.075 50.985 76.075 50.985 75.695 50.655 75.695 50.655 76.075 49.625 76.075 49.625 75.615 49.32 75.615 49.32 76.075 47.835 76.075 47.835 75.635 47.645 75.635 47.645 76.075 45.745 76.075 45.745 75.615 45.415 75.615 45.415 76.075 42.815 76.075 42.815 75.715 42.485 75.715 42.485 76.075 41.785 76.075 41.785 75.695 41.455 75.695 41.455 76.075 40.425 76.075 40.425 75.615 40.12 75.615 40.12 76.075 38.635 76.075 38.635 75.635 38.445 75.635 38.445 76.075 36.545 76.075 36.545 75.615 36.215 75.615 36.215 76.075 33.615 76.075 33.615 75.715 33.285 75.715 33.285 76.075 32.585 76.075 32.585 75.695 32.255 75.695 32.255 76.075 31.225 76.075 31.225 75.615 30.92 75.615 30.92 76.075 29.435 76.075 29.435 75.635 29.245 75.635 29.245 76.075 27.345 76.075 27.345 75.615 27.015 75.615 27.015 76.075 24.415 76.075 24.415 75.715 24.085 75.715 24.085 76.075 23.385 76.075 23.385 75.695 23.055 75.695 23.055 76.075 22.025 76.075 22.025 75.615 21.72 75.615 21.72 76.075 20.235 76.075 20.235 75.635 20.045 75.635 20.045 76.075 18.145 76.075 18.145 75.615 17.815 75.615 17.815 76.075 15.215 76.075 15.215 75.715 14.885 75.715 14.885 76.075 14.185 76.075 14.185 75.695 13.855 75.695 13.855 76.075 10.875 76.075 10.875 75.675 10.545 75.675 10.545 76.075 10.035 76.075 10.035 75.675 9.705 75.675 9.705 76.075 8.29 76.075 8.29 75.565 7.875 75.565 7.875 76.075 6.765 76.075 6.765 75.615 6.46 75.615 6.46 76.075 5.79 76.075 5.79 75.615 5.62 75.615 5.62 76.075 4.95 76.075 4.95 75.615 4.78 75.615 4.78 76.075 4.11 76.075 4.11 75.615 3.94 75.615 3.94 76.075 3.27 76.075 3.27 75.615 3.015 75.615 3.015 76.075 0 76.075 0 76.245 ;
      RECT 74.52 73.355 75.44 73.525 ;
      RECT 0 73.355 1.84 73.525 ;
      RECT 74.52 70.635 75.44 70.805 ;
      RECT 0 70.635 1.84 70.805 ;
      RECT 74.52 67.915 75.44 68.085 ;
      RECT 0 67.915 1.84 68.085 ;
      RECT 74.52 65.195 75.44 65.365 ;
      RECT 0 65.195 1.84 65.365 ;
      RECT 74.52 62.475 75.44 62.645 ;
      RECT 0 62.475 1.84 62.645 ;
      RECT 74.52 59.755 75.44 59.925 ;
      RECT 0 59.755 1.84 59.925 ;
      RECT 74.52 57.035 75.44 57.205 ;
      RECT 0 57.035 1.84 57.205 ;
      RECT 74.52 54.315 75.44 54.485 ;
      RECT 0 54.315 1.84 54.485 ;
      RECT 74.52 51.595 75.44 51.765 ;
      RECT 0 51.595 1.84 51.765 ;
      RECT 74.52 48.875 75.44 49.045 ;
      RECT 0 48.875 1.84 49.045 ;
      RECT 74.52 46.155 75.44 46.325 ;
      RECT 0 46.155 3.68 46.325 ;
      RECT 74.52 43.435 75.44 43.605 ;
      RECT 0 43.435 3.68 43.605 ;
      RECT 74.52 40.715 75.44 40.885 ;
      RECT 0 40.715 1.84 40.885 ;
      RECT 74.52 37.995 75.44 38.165 ;
      RECT 0 37.995 1.84 38.165 ;
      RECT 74.52 35.275 75.44 35.445 ;
      RECT 0 35.275 1.84 35.445 ;
      RECT 74.52 32.555 75.44 32.725 ;
      RECT 0 32.555 1.84 32.725 ;
      RECT 71.76 29.835 75.44 30.005 ;
      RECT 0 29.835 1.84 30.005 ;
      RECT 71.76 27.115 75.44 27.285 ;
      RECT 0 27.115 1.84 27.285 ;
      RECT 74.52 24.395 75.44 24.565 ;
      RECT 0 24.395 1.84 24.565 ;
      RECT 74.52 21.675 75.44 21.845 ;
      RECT 0 21.675 1.84 21.845 ;
      RECT 74.52 18.955 75.44 19.125 ;
      RECT 0 18.955 1.84 19.125 ;
      RECT 74.52 16.235 75.44 16.405 ;
      RECT 0 16.235 1.84 16.405 ;
      RECT 74.52 13.515 75.44 13.685 ;
      RECT 0 13.515 1.84 13.685 ;
      RECT 74.52 10.795 75.44 10.965 ;
      RECT 0 10.795 1.84 10.965 ;
      RECT 74.52 8.075 75.44 8.245 ;
      RECT 0 8.075 3.68 8.245 ;
      RECT 74.52 5.355 75.44 5.525 ;
      RECT 0 5.355 3.68 5.525 ;
      RECT 74.52 2.635 75.44 2.805 ;
      RECT 0 2.635 1.84 2.805 ;
      POLYGON 49.555 0.905 49.555 0.085 50.195 0.085 50.195 0.465 50.525 0.465 50.525 0.085 51.225 0.085 51.225 0.445 51.555 0.445 51.555 0.085 54.155 0.085 54.155 0.545 54.485 0.545 54.485 0.085 56.385 0.085 56.385 0.525 56.575 0.525 56.575 0.085 58.06 0.085 58.06 0.545 58.365 0.545 58.365 0.085 59.355 0.085 59.355 0.885 59.685 0.885 59.685 0.085 60.195 0.085 60.195 0.565 60.525 0.565 60.525 0.085 61.035 0.085 61.035 0.565 61.365 0.565 61.365 0.085 61.875 0.085 61.875 0.565 62.205 0.565 62.205 0.085 62.715 0.085 62.715 0.565 63.045 0.565 63.045 0.085 63.555 0.085 63.555 0.565 63.885 0.565 63.885 0.085 64.835 0.085 64.835 0.565 65.005 0.565 65.005 0.085 65.675 0.085 65.675 0.565 65.845 0.565 65.845 0.085 66.435 0.085 66.435 0.565 66.765 0.565 66.765 0.085 67.275 0.085 67.275 0.565 67.605 0.565 67.605 0.085 68.115 0.085 68.115 0.885 68.445 0.885 68.445 0.085 70.445 0.085 70.445 0.565 70.685 0.565 70.685 0.085 71.275 0.085 71.275 0.565 71.605 0.565 71.605 0.085 72.115 0.085 72.115 0.885 72.445 0.885 72.445 0.085 75.44 0.085 75.44 -0.085 0 -0.085 0 0.085 3.195 0.085 3.195 0.565 3.365 0.565 3.365 0.085 4.035 0.085 4.035 0.565 4.205 0.565 4.205 0.085 4.795 0.085 4.795 0.565 5.125 0.565 5.125 0.085 5.635 0.085 5.635 0.565 5.965 0.565 5.965 0.085 6.475 0.085 6.475 0.885 6.805 0.885 6.805 0.085 8.375 0.085 8.375 0.885 8.705 0.885 8.705 0.085 9.215 0.085 9.215 0.565 9.545 0.565 9.545 0.085 10.055 0.085 10.055 0.565 10.385 0.565 10.385 0.085 10.975 0.085 10.975 0.565 11.145 0.565 11.145 0.085 11.815 0.085 11.815 0.565 11.985 0.565 11.985 0.085 14.885 0.085 14.885 0.485 15.215 0.485 15.215 0.085 15.725 0.085 15.725 0.485 16.055 0.485 16.055 0.085 17.47 0.085 17.47 0.595 17.885 0.595 17.885 0.085 18.495 0.085 18.495 0.885 18.825 0.885 18.825 0.085 19.335 0.085 19.335 0.565 19.665 0.565 19.665 0.085 20.175 0.085 20.175 0.565 20.505 0.565 20.505 0.085 21.095 0.085 21.095 0.565 21.265 0.565 21.265 0.085 21.935 0.085 21.935 0.565 22.105 0.565 22.105 0.085 22.725 0.085 22.725 0.55 22.975 0.55 22.975 0.085 23.565 0.085 23.565 0.545 23.735 0.545 23.735 0.085 24.405 0.085 24.405 0.545 24.575 0.545 24.575 0.085 25.365 0.085 25.365 0.545 25.63 0.545 25.63 0.085 25.855 0.085 25.855 0.885 26.185 0.885 26.185 0.085 26.695 0.085 26.695 0.565 27.025 0.565 27.025 0.085 27.535 0.085 27.535 0.565 27.865 0.565 27.865 0.085 28.455 0.085 28.455 0.565 28.625 0.565 28.625 0.085 29.295 0.085 29.295 0.565 29.465 0.565 29.465 0.085 30.915 0.085 30.915 0.885 31.245 0.885 31.245 0.085 31.755 0.085 31.755 0.565 32.085 0.565 32.085 0.085 32.595 0.085 32.595 0.565 32.925 0.565 32.925 0.085 33.515 0.085 33.515 0.565 33.685 0.565 33.685 0.085 34.355 0.085 34.355 0.565 34.525 0.565 34.525 0.085 35.215 0.085 35.215 0.545 35.47 0.545 35.47 0.085 36.14 0.085 36.14 0.545 36.31 0.545 36.31 0.085 36.98 0.085 36.98 0.545 37.15 0.545 37.15 0.085 37.82 0.085 37.82 0.545 37.99 0.545 37.99 0.085 38.66 0.085 38.66 0.545 38.965 0.545 38.965 0.085 39.615 0.085 39.615 0.465 39.945 0.465 39.945 0.085 40.645 0.085 40.645 0.445 40.975 0.445 40.975 0.085 43.575 0.085 43.575 0.545 43.905 0.545 43.905 0.085 45.805 0.085 45.805 0.525 45.995 0.525 45.995 0.085 47.48 0.085 47.48 0.545 47.785 0.545 47.785 0.085 48.445 0.085 48.445 0.905 48.655 0.905 48.655 0.085 49.325 0.085 49.325 0.905 ;
      RECT 0.17 0.17 75.27 75.99 ;
    LAYER via ;
      RECT 52.365 75.965 52.515 76.115 ;
      RECT 22.925 75.965 23.075 76.115 ;
      RECT 32.355 0.435 32.505 0.585 ;
      RECT 16.255 0.435 16.405 0.585 ;
      RECT 2.455 0.435 2.605 0.585 ;
      RECT 52.365 0.045 52.515 0.195 ;
      RECT 22.925 0.045 23.075 0.195 ;
    LAYER via2 ;
      RECT 52.34 75.94 52.54 76.14 ;
      RECT 22.9 75.94 23.1 76.14 ;
      RECT 74.19 13.84 74.39 14.04 ;
      RECT 52.34 0.02 52.54 0.22 ;
      RECT 22.9 0.02 23.1 0.22 ;
    LAYER via3 ;
      RECT 52.34 75.94 52.54 76.14 ;
      RECT 22.9 75.94 23.1 76.14 ;
      RECT 52.34 0.02 52.54 0.22 ;
      RECT 22.9 0.02 23.1 0.22 ;
    LAYER OVERLAP ;
      POLYGON 0 0 0 76.16 75.44 76.16 75.44 0 ;
  END
END cbx_1__2_

END LIBRARY
