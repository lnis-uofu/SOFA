VERSION 5.7 ;
BUSBITCHARS "[]" ;

UNITS
  DATABASE MICRONS 1000 ;
END UNITS

MANUFACTURINGGRID 0.005 ;

LAYER li1
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.46 ;
  WIDTH 0.17 ;
END li1

LAYER mcon
  TYPE CUT ;
END mcon

LAYER met1
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.34 ;
  WIDTH 0.14 ;
END met1

LAYER via
  TYPE CUT ;
END via

LAYER met2
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.46 ;
  WIDTH 0.14 ;
END met2

LAYER via2
  TYPE CUT ;
END via2

LAYER met3
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.68 ;
  WIDTH 0.3 ;
END met3

LAYER via3
  TYPE CUT ;
END via3

LAYER met4
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.92 ;
  WIDTH 0.3 ;
END met4

LAYER via4
  TYPE CUT ;
END via4

LAYER met5
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 3.4 ;
  WIDTH 1.6 ;
END met5

LAYER nwell
  TYPE MASTERSLICE ;
END nwell

LAYER pwell
  TYPE MASTERSLICE ;
END pwell

LAYER OVERLAP
  TYPE OVERLAP ;
END OVERLAP

VIA L1M1_PR
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.145 -0.115 0.145 0.115 ;
END L1M1_PR

VIA L1M1_PR_R
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.115 -0.145 0.115 0.145 ;
END L1M1_PR_R

VIA L1M1_PR_M
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.115 -0.145 0.115 0.145 ;
END L1M1_PR_M

VIA L1M1_PR_MR
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.145 -0.115 0.145 0.115 ;
END L1M1_PR_MR

VIA L1M1_PR_C
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.145 -0.145 0.145 0.145 ;
END L1M1_PR_C

VIA M1M2_PR
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR

VIA M1M2_PR_Enc
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_Enc

VIA M1M2_PR_R
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_R

VIA M1M2_PR_R_Enc
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR_R_Enc

VIA M1M2_PR_M
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_M

VIA M1M2_PR_M_Enc
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR_M_Enc

VIA M1M2_PR_MR
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR_MR

VIA M1M2_PR_MR_Enc
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_MR_Enc

VIA M1M2_PR_C
  LAYER met1 ;
    RECT -0.16 -0.16 0.16 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.16 0.16 0.16 ;
END M1M2_PR_C

VIA M2M3_PR
  LAYER met2 ;
    RECT -0.14 -0.185 0.14 0.185 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR

VIA M2M3_PR_R
  LAYER met2 ;
    RECT -0.185 -0.14 0.185 0.14 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_R

VIA M2M3_PR_M
  LAYER met2 ;
    RECT -0.14 -0.185 0.14 0.185 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_M

VIA M2M3_PR_MR
  LAYER met2 ;
    RECT -0.185 -0.14 0.185 0.14 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_MR

VIA M2M3_PR_C
  LAYER met2 ;
    RECT -0.185 -0.185 0.185 0.185 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_C

VIA M3M4_PR
  LAYER met3 ;
    RECT -0.19 -0.16 0.19 0.16 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR

VIA M3M4_PR_R
  LAYER met3 ;
    RECT -0.16 -0.19 0.16 0.19 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_R

VIA M3M4_PR_M
  LAYER met3 ;
    RECT -0.19 -0.16 0.19 0.16 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_M

VIA M3M4_PR_MR
  LAYER met3 ;
    RECT -0.16 -0.19 0.16 0.19 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_MR

VIA M3M4_PR_C
  LAYER met3 ;
    RECT -0.19 -0.19 0.19 0.19 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_C

VIA M4M5_PR
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR

VIA M4M5_PR_R
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_R

VIA M4M5_PR_M
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_M

VIA M4M5_PR_MR
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_MR

VIA M4M5_PR_C
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_C

SITE unit
  CLASS CORE ;
  SYMMETRY Y ;
  SIZE 0.46 BY 2.72 ;
END unit

SITE unithddbl
  CLASS CORE ;
  SIZE 0.46 BY 5.44 ;
END unithddbl

MACRO sb_2__0_
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  SIZE 92 BY 97.92 ;
  SYMMETRY X Y ;
  PIN chany_top_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.74 97.435 56.88 97.92 ;
    END
  END chany_top_in[0]
  PIN chany_top_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.04 97.435 59.18 97.92 ;
    END
  END chany_top_in[1]
  PIN chany_top_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.02 97.435 65.16 97.92 ;
    END
  END chany_top_in[2]
  PIN chany_top_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.08 97.435 70.22 97.92 ;
    END
  END chany_top_in[3]
  PIN chany_top_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.18 97.435 63.32 97.92 ;
    END
  END chany_top_in[4]
  PIN chany_top_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.78 97.435 67.92 97.92 ;
    END
  END chany_top_in[5]
  PIN chany_top_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.14 97.435 52.28 97.92 ;
    END
  END chany_top_in[6]
  PIN chany_top_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.06 97.435 53.2 97.92 ;
    END
  END chany_top_in[7]
  PIN chany_top_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.7 97.435 45.84 97.92 ;
    END
  END chany_top_in[8]
  PIN chany_top_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.94 97.435 66.08 97.92 ;
    END
  END chany_top_in[9]
  PIN chany_top_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.1 97.435 64.24 97.92 ;
    END
  END chany_top_in[10]
  PIN chany_top_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.68 97.435 74.82 97.92 ;
    END
  END chany_top_in[11]
  PIN chany_top_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.26 97.435 62.4 97.92 ;
    END
  END chany_top_in[12]
  PIN chany_top_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.84 97.435 72.98 97.92 ;
    END
  END chany_top_in[13]
  PIN chany_top_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.98 97.435 54.12 97.92 ;
    END
  END chany_top_in[14]
  PIN chany_top_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.12 97.435 58.26 97.92 ;
    END
  END chany_top_in[15]
  PIN chany_top_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.46 97.435 48.6 97.92 ;
    END
  END chany_top_in[16]
  PIN chany_top_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.76 97.435 73.9 97.92 ;
    END
  END chany_top_in[17]
  PIN chany_top_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.78 97.435 44.92 97.92 ;
    END
  END chany_top_in[18]
  PIN chany_top_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.16 97.435 69.3 97.92 ;
    END
  END chany_top_in[19]
  PIN top_left_grid_pin_42_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.5 86.555 13.64 87.04 ;
    END
  END top_left_grid_pin_42_[0]
  PIN top_left_grid_pin_43_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.66 86.555 11.8 87.04 ;
    END
  END top_left_grid_pin_43_[0]
  PIN top_left_grid_pin_44_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.44 86.555 8.58 87.04 ;
    END
  END top_left_grid_pin_44_[0]
  PIN top_left_grid_pin_45_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.58 86.555 12.72 87.04 ;
    END
  END top_left_grid_pin_45_[0]
  PIN top_left_grid_pin_46_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.28 86.555 10.42 87.04 ;
    END
  END top_left_grid_pin_46_[0]
  PIN top_left_grid_pin_47_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.3 86.555 4.44 87.04 ;
    END
  END top_left_grid_pin_47_[0]
  PIN top_left_grid_pin_48_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.36 86.555 9.5 87.04 ;
    END
  END top_left_grid_pin_48_[0]
  PIN top_left_grid_pin_49_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.06 86.555 7.2 87.04 ;
    END
  END top_left_grid_pin_49_[0]
  PIN top_right_grid_pin_1_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.44 97.435 31.58 97.92 ;
    END
  END top_right_grid_pin_1_[0]
  PIN chanx_left_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 36.91 0.8 37.21 ;
    END
  END chanx_left_in[0]
  PIN chanx_left_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 21.27 0.8 21.57 ;
    END
  END chanx_left_in[1]
  PIN chanx_left_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 63.43 0.8 63.73 ;
    END
  END chanx_left_in[2]
  PIN chanx_left_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 47.11 0.8 47.41 ;
    END
  END chanx_left_in[3]
  PIN chanx_left_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 45.75 0.8 46.05 ;
    END
  END chanx_left_in[4]
  PIN chanx_left_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 49.83 0.8 50.13 ;
    END
  END chanx_left_in[5]
  PIN chanx_left_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 60.71 0.8 61.01 ;
    END
  END chanx_left_in[6]
  PIN chanx_left_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 55.95 0.8 56.25 ;
    END
  END chanx_left_in[7]
  PIN chanx_left_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 64.79 0.8 65.09 ;
    END
  END chanx_left_in[8]
  PIN chanx_left_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 51.19 0.8 51.49 ;
    END
  END chanx_left_in[9]
  PIN chanx_left_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 29.43 0.8 29.73 ;
    END
  END chanx_left_in[10]
  PIN chanx_left_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 15.83 0.8 16.13 ;
    END
  END chanx_left_in[11]
  PIN chanx_left_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 68.19 0.8 68.49 ;
    END
  END chanx_left_in[12]
  PIN chanx_left_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 48.47 0.8 48.77 ;
    END
  END chanx_left_in[13]
  PIN chanx_left_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 38.27 0.8 38.57 ;
    END
  END chanx_left_in[14]
  PIN chanx_left_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 57.31 0.8 57.61 ;
    END
  END chanx_left_in[15]
  PIN chanx_left_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 62.07 0.8 62.37 ;
    END
  END chanx_left_in[16]
  PIN chanx_left_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 73.63 0.8 73.93 ;
    END
  END chanx_left_in[17]
  PIN chanx_left_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 59.35 0.8 59.65 ;
    END
  END chanx_left_in[18]
  PIN chanx_left_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 78.39 0.8 78.69 ;
    END
  END chanx_left_in[19]
  PIN left_bottom_grid_pin_1_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 26.71 0.8 27.01 ;
    END
  END left_bottom_grid_pin_1_[0]
  PIN left_bottom_grid_pin_3_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 25.35 0.8 25.65 ;
    END
  END left_bottom_grid_pin_3_[0]
  PIN left_bottom_grid_pin_5_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 14.47 0.8 14.77 ;
    END
  END left_bottom_grid_pin_5_[0]
  PIN left_bottom_grid_pin_7_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 32.83 0.8 33.13 ;
    END
  END left_bottom_grid_pin_7_[0]
  PIN left_bottom_grid_pin_9_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 13.11 0.8 13.41 ;
    END
  END left_bottom_grid_pin_9_[0]
  PIN left_bottom_grid_pin_11_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 23.99 0.8 24.29 ;
    END
  END left_bottom_grid_pin_11_[0]
  PIN left_bottom_grid_pin_13_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 22.63 0.8 22.93 ;
    END
  END left_bottom_grid_pin_13_[0]
  PIN left_bottom_grid_pin_15_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 11.75 0.8 12.05 ;
    END
  END left_bottom_grid_pin_15_[0]
  PIN left_bottom_grid_pin_17_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 19.91 0.8 20.21 ;
    END
  END left_bottom_grid_pin_17_[0]
  PIN ccff_head[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.52 97.435 30.66 97.92 ;
    END
  END ccff_head[0]
  PIN chany_top_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.52 97.435 76.66 97.92 ;
    END
  END chany_top_out[0]
  PIN chany_top_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.86 97.435 44 97.92 ;
    END
  END chany_top_out[1]
  PIN chany_top_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.6 97.435 75.74 97.92 ;
    END
  END chany_top_out[2]
  PIN chany_top_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.44 97.435 77.58 97.92 ;
    END
  END chany_top_out[3]
  PIN chany_top_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.96 97.435 60.1 97.92 ;
    END
  END chany_top_out[4]
  PIN chany_top_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.62 97.435 46.76 97.92 ;
    END
  END chany_top_out[5]
  PIN chany_top_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.9 97.435 55.04 97.92 ;
    END
  END chany_top_out[6]
  PIN chany_top_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.36 97.435 78.5 97.92 ;
    END
  END chany_top_out[7]
  PIN chany_top_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.86 97.435 67 97.92 ;
    END
  END chany_top_out[8]
  PIN chany_top_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.82 97.435 55.96 97.92 ;
    END
  END chany_top_out[9]
  PIN chany_top_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.54 97.435 47.68 97.92 ;
    END
  END chany_top_out[10]
  PIN chany_top_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.34 97.435 61.48 97.92 ;
    END
  END chany_top_out[11]
  PIN chany_top_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.34 97.435 38.48 97.92 ;
    END
  END chany_top_out[12]
  PIN chany_top_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.28 97.435 79.42 97.92 ;
    END
  END chany_top_out[13]
  PIN chany_top_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.76 97.435 50.9 97.92 ;
    END
  END chany_top_out[14]
  PIN chany_top_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.84 97.435 49.98 97.92 ;
    END
  END chany_top_out[15]
  PIN chany_top_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.36 97.435 32.5 97.92 ;
    END
  END chany_top_out[16]
  PIN chany_top_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.92 97.435 72.06 97.92 ;
    END
  END chany_top_out[17]
  PIN chany_top_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.28 97.435 33.42 97.92 ;
    END
  END chany_top_out[18]
  PIN chany_top_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71 97.435 71.14 97.92 ;
    END
  END chany_top_out[19]
  PIN chanx_left_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 53.23 0.8 53.53 ;
    END
  END chanx_left_out[0]
  PIN chanx_left_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 74.99 0.8 75.29 ;
    END
  END chanx_left_out[1]
  PIN chanx_left_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 54.59 0.8 54.89 ;
    END
  END chanx_left_out[2]
  PIN chanx_left_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 44.39 0.8 44.69 ;
    END
  END chanx_left_out[3]
  PIN chanx_left_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 77.03 0.8 77.33 ;
    END
  END chanx_left_out[4]
  PIN chanx_left_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 31.47 0.8 31.77 ;
    END
  END chanx_left_out[5]
  PIN chanx_left_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 69.55 0.8 69.85 ;
    END
  END chanx_left_out[6]
  PIN chanx_left_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 18.55 0.8 18.85 ;
    END
  END chanx_left_out[7]
  PIN chanx_left_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 34.19 0.8 34.49 ;
    END
  END chanx_left_out[8]
  PIN chanx_left_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 66.83 0.8 67.13 ;
    END
  END chanx_left_out[9]
  PIN chanx_left_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 43.03 0.8 43.33 ;
    END
  END chanx_left_out[10]
  PIN chanx_left_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 39.63 0.8 39.93 ;
    END
  END chanx_left_out[11]
  PIN chanx_left_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 35.55 0.8 35.85 ;
    END
  END chanx_left_out[12]
  PIN chanx_left_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 72.27 0.8 72.57 ;
    END
  END chanx_left_out[13]
  PIN chanx_left_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 79.75 0.8 80.05 ;
    END
  END chanx_left_out[14]
  PIN chanx_left_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 83.15 0.8 83.45 ;
    END
  END chanx_left_out[15]
  PIN chanx_left_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 17.19 0.8 17.49 ;
    END
  END chanx_left_out[16]
  PIN chanx_left_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 28.07 0.8 28.37 ;
    END
  END chanx_left_out[17]
  PIN chanx_left_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 41.67 0.8 41.97 ;
    END
  END chanx_left_out[18]
  PIN chanx_left_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 70.91 0.8 71.21 ;
    END
  END chanx_left_out[19]
  PIN ccff_tail[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 81.11 0.8 81.41 ;
    END
  END ccff_tail[0]
  PIN prog_clk_0_N_in
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER met2 ;
        RECT 37.42 97.435 37.56 97.92 ;
    END
  END prog_clk_0_N_in
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0 11.32 3.2 14.52 ;
        RECT 88.8 11.32 92 14.52 ;
        RECT 0 52.12 3.2 55.32 ;
        RECT 88.8 52.12 92 55.32 ;
      LAYER met4 ;
        RECT 36.5 0 37.1 0.6 ;
        RECT 65.94 0 66.54 0.6 ;
        RECT 36.5 97.32 37.1 97.92 ;
        RECT 65.94 97.32 66.54 97.92 ;
      LAYER met1 ;
        RECT 0 2.48 0.48 2.96 ;
        RECT 91.52 2.48 92 2.96 ;
        RECT 0 7.92 0.48 8.4 ;
        RECT 91.52 7.92 92 8.4 ;
        RECT 0 13.36 0.48 13.84 ;
        RECT 91.52 13.36 92 13.84 ;
        RECT 0 18.8 0.48 19.28 ;
        RECT 91.52 18.8 92 19.28 ;
        RECT 0 24.24 0.48 24.72 ;
        RECT 91.52 24.24 92 24.72 ;
        RECT 0 29.68 0.48 30.16 ;
        RECT 91.52 29.68 92 30.16 ;
        RECT 0 35.12 0.48 35.6 ;
        RECT 91.52 35.12 92 35.6 ;
        RECT 0 40.56 0.48 41.04 ;
        RECT 91.52 40.56 92 41.04 ;
        RECT 0 46 0.48 46.48 ;
        RECT 91.52 46 92 46.48 ;
        RECT 0 51.44 0.48 51.92 ;
        RECT 91.52 51.44 92 51.92 ;
        RECT 0 56.88 0.48 57.36 ;
        RECT 91.52 56.88 92 57.36 ;
        RECT 0 62.32 0.48 62.8 ;
        RECT 91.52 62.32 92 62.8 ;
        RECT 0 67.76 0.48 68.24 ;
        RECT 91.52 67.76 92 68.24 ;
        RECT 0 73.2 0.48 73.68 ;
        RECT 91.52 73.2 92 73.68 ;
        RECT 0 78.64 0.48 79.12 ;
        RECT 91.52 78.64 92 79.12 ;
        RECT 0 84.08 0.48 84.56 ;
        RECT 91.52 84.08 92 84.56 ;
        RECT 25.76 89.52 26.24 90 ;
        RECT 91.52 89.52 92 90 ;
        RECT 25.76 94.96 26.24 95.44 ;
        RECT 91.52 94.96 92 95.44 ;
    END
  END VDD
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 10.74 0 11.34 0.6 ;
        RECT 51.22 0 51.82 0.6 ;
        RECT 80.66 0 81.26 0.6 ;
        RECT 10.74 86.44 11.34 87.04 ;
        RECT 51.22 97.32 51.82 97.92 ;
        RECT 80.66 97.32 81.26 97.92 ;
      LAYER met5 ;
        RECT 0 31.72 3.2 34.92 ;
        RECT 88.8 31.72 92 34.92 ;
        RECT 0 72.52 3.2 75.72 ;
        RECT 88.8 72.52 92 75.72 ;
      LAYER met1 ;
        RECT 0 0 45.4 0.24 ;
        RECT 46.6 0 92 0.24 ;
        RECT 0 5.2 0.48 5.68 ;
        RECT 91.52 5.2 92 5.68 ;
        RECT 0 10.64 0.48 11.12 ;
        RECT 91.52 10.64 92 11.12 ;
        RECT 0 16.08 0.48 16.56 ;
        RECT 91.52 16.08 92 16.56 ;
        RECT 0 21.52 0.48 22 ;
        RECT 91.52 21.52 92 22 ;
        RECT 0 26.96 0.48 27.44 ;
        RECT 91.52 26.96 92 27.44 ;
        RECT 0 32.4 0.48 32.88 ;
        RECT 91.52 32.4 92 32.88 ;
        RECT 0 37.84 0.48 38.32 ;
        RECT 91.52 37.84 92 38.32 ;
        RECT 0 43.28 0.48 43.76 ;
        RECT 91.52 43.28 92 43.76 ;
        RECT 0 48.72 0.48 49.2 ;
        RECT 91.52 48.72 92 49.2 ;
        RECT 0 54.16 0.48 54.64 ;
        RECT 91.52 54.16 92 54.64 ;
        RECT 0 59.6 0.48 60.08 ;
        RECT 91.52 59.6 92 60.08 ;
        RECT 0 65.04 0.48 65.52 ;
        RECT 91.52 65.04 92 65.52 ;
        RECT 0 70.48 0.48 70.96 ;
        RECT 91.52 70.48 92 70.96 ;
        RECT 0 75.92 0.48 76.4 ;
        RECT 91.52 75.92 92 76.4 ;
        RECT 0 81.36 0.48 81.84 ;
        RECT 91.52 81.36 92 81.84 ;
        RECT 0 86.8 45.4 87.28 ;
        RECT 91.52 86.8 92 87.28 ;
        RECT 25.76 92.24 26.24 92.72 ;
        RECT 91.52 92.24 92 92.72 ;
        RECT 25.76 97.68 45.4 97.92 ;
        RECT 46.6 97.68 92 97.92 ;
    END
  END VSS
  OBS
    LAYER met2 ;
      RECT 80.82 97.735 81.1 98.105 ;
      RECT 51.38 97.735 51.66 98.105 ;
      RECT 10.9 86.855 11.18 87.225 ;
      RECT 80.82 -0.185 81.1 0.185 ;
      RECT 51.38 -0.185 51.66 0.185 ;
      RECT 10.9 -0.185 11.18 0.185 ;
      POLYGON 91.72 97.64 91.72 0.28 0.28 0.28 0.28 86.76 4.02 86.76 4.02 86.275 4.72 86.275 4.72 86.76 6.78 86.76 6.78 86.275 7.48 86.275 7.48 86.76 8.16 86.76 8.16 86.275 8.86 86.275 8.86 86.76 9.08 86.76 9.08 86.275 9.78 86.275 9.78 86.76 10 86.76 10 86.275 10.7 86.275 10.7 86.76 11.38 86.76 11.38 86.275 12.08 86.275 12.08 86.76 12.3 86.76 12.3 86.275 13 86.275 13 86.76 13.22 86.76 13.22 86.275 13.92 86.275 13.92 86.76 26.04 86.76 26.04 97.64 30.24 97.64 30.24 97.155 30.94 97.155 30.94 97.64 31.16 97.64 31.16 97.155 31.86 97.155 31.86 97.64 32.08 97.64 32.08 97.155 32.78 97.155 32.78 97.64 33 97.64 33 97.155 33.7 97.155 33.7 97.64 37.14 97.64 37.14 97.155 37.84 97.155 37.84 97.64 38.06 97.64 38.06 97.155 38.76 97.155 38.76 97.64 43.58 97.64 43.58 97.155 44.28 97.155 44.28 97.64 44.5 97.64 44.5 97.155 45.2 97.155 45.2 97.64 45.42 97.64 45.42 97.155 46.12 97.155 46.12 97.64 46.34 97.64 46.34 97.155 47.04 97.155 47.04 97.64 47.26 97.64 47.26 97.155 47.96 97.155 47.96 97.64 48.18 97.64 48.18 97.155 48.88 97.155 48.88 97.64 49.56 97.64 49.56 97.155 50.26 97.155 50.26 97.64 50.48 97.64 50.48 97.155 51.18 97.155 51.18 97.64 51.86 97.64 51.86 97.155 52.56 97.155 52.56 97.64 52.78 97.64 52.78 97.155 53.48 97.155 53.48 97.64 53.7 97.64 53.7 97.155 54.4 97.155 54.4 97.64 54.62 97.64 54.62 97.155 55.32 97.155 55.32 97.64 55.54 97.64 55.54 97.155 56.24 97.155 56.24 97.64 56.46 97.64 56.46 97.155 57.16 97.155 57.16 97.64 57.84 97.64 57.84 97.155 58.54 97.155 58.54 97.64 58.76 97.64 58.76 97.155 59.46 97.155 59.46 97.64 59.68 97.64 59.68 97.155 60.38 97.155 60.38 97.64 61.06 97.64 61.06 97.155 61.76 97.155 61.76 97.64 61.98 97.64 61.98 97.155 62.68 97.155 62.68 97.64 62.9 97.64 62.9 97.155 63.6 97.155 63.6 97.64 63.82 97.64 63.82 97.155 64.52 97.155 64.52 97.64 64.74 97.64 64.74 97.155 65.44 97.155 65.44 97.64 65.66 97.64 65.66 97.155 66.36 97.155 66.36 97.64 66.58 97.64 66.58 97.155 67.28 97.155 67.28 97.64 67.5 97.64 67.5 97.155 68.2 97.155 68.2 97.64 68.88 97.64 68.88 97.155 69.58 97.155 69.58 97.64 69.8 97.64 69.8 97.155 70.5 97.155 70.5 97.64 70.72 97.64 70.72 97.155 71.42 97.155 71.42 97.64 71.64 97.64 71.64 97.155 72.34 97.155 72.34 97.64 72.56 97.64 72.56 97.155 73.26 97.155 73.26 97.64 73.48 97.64 73.48 97.155 74.18 97.155 74.18 97.64 74.4 97.64 74.4 97.155 75.1 97.155 75.1 97.64 75.32 97.64 75.32 97.155 76.02 97.155 76.02 97.64 76.24 97.64 76.24 97.155 76.94 97.155 76.94 97.64 77.16 97.64 77.16 97.155 77.86 97.155 77.86 97.64 78.08 97.64 78.08 97.155 78.78 97.155 78.78 97.64 79 97.64 79 97.155 79.7 97.155 79.7 97.64 ;
    LAYER met3 ;
      POLYGON 81.125 98.085 81.125 98.08 81.34 98.08 81.34 97.76 81.125 97.76 81.125 97.755 80.795 97.755 80.795 97.76 80.58 97.76 80.58 98.08 80.795 98.08 80.795 98.085 ;
      POLYGON 51.685 98.085 51.685 98.08 51.9 98.08 51.9 97.76 51.685 97.76 51.685 97.755 51.355 97.755 51.355 97.76 51.14 97.76 51.14 98.08 51.355 98.08 51.355 98.085 ;
      POLYGON 11.205 87.205 11.205 87.2 11.42 87.2 11.42 86.88 11.205 86.88 11.205 86.875 10.875 86.875 10.875 86.88 10.66 86.88 10.66 87.2 10.875 87.2 10.875 87.205 ;
      POLYGON 81.125 0.165 81.125 0.16 81.34 0.16 81.34 -0.16 81.125 -0.16 81.125 -0.165 80.795 -0.165 80.795 -0.16 80.58 -0.16 80.58 0.16 80.795 0.16 80.795 0.165 ;
      POLYGON 51.685 0.165 51.685 0.16 51.9 0.16 51.9 -0.16 51.685 -0.16 51.685 -0.165 51.355 -0.165 51.355 -0.16 51.14 -0.16 51.14 0.16 51.355 0.16 51.355 0.165 ;
      POLYGON 11.205 0.165 11.205 0.16 11.42 0.16 11.42 -0.16 11.205 -0.16 11.205 -0.165 10.875 -0.165 10.875 -0.16 10.66 -0.16 10.66 0.16 10.875 0.16 10.875 0.165 ;
      POLYGON 91.6 97.52 91.6 0.4 0.4 0.4 0.4 11.35 1.2 11.35 1.2 12.45 0.4 12.45 0.4 12.71 1.2 12.71 1.2 13.81 0.4 13.81 0.4 14.07 1.2 14.07 1.2 15.17 0.4 15.17 0.4 15.43 1.2 15.43 1.2 16.53 0.4 16.53 0.4 16.79 1.2 16.79 1.2 17.89 0.4 17.89 0.4 18.15 1.2 18.15 1.2 19.25 0.4 19.25 0.4 19.51 1.2 19.51 1.2 20.61 0.4 20.61 0.4 20.87 1.2 20.87 1.2 21.97 0.4 21.97 0.4 22.23 1.2 22.23 1.2 23.33 0.4 23.33 0.4 23.59 1.2 23.59 1.2 24.69 0.4 24.69 0.4 24.95 1.2 24.95 1.2 26.05 0.4 26.05 0.4 26.31 1.2 26.31 1.2 27.41 0.4 27.41 0.4 27.67 1.2 27.67 1.2 28.77 0.4 28.77 0.4 29.03 1.2 29.03 1.2 30.13 0.4 30.13 0.4 31.07 1.2 31.07 1.2 32.17 0.4 32.17 0.4 32.43 1.2 32.43 1.2 33.53 0.4 33.53 0.4 33.79 1.2 33.79 1.2 34.89 0.4 34.89 0.4 35.15 1.2 35.15 1.2 36.25 0.4 36.25 0.4 36.51 1.2 36.51 1.2 37.61 0.4 37.61 0.4 37.87 1.2 37.87 1.2 38.97 0.4 38.97 0.4 39.23 1.2 39.23 1.2 40.33 0.4 40.33 0.4 41.27 1.2 41.27 1.2 42.37 0.4 42.37 0.4 42.63 1.2 42.63 1.2 43.73 0.4 43.73 0.4 43.99 1.2 43.99 1.2 45.09 0.4 45.09 0.4 45.35 1.2 45.35 1.2 46.45 0.4 46.45 0.4 46.71 1.2 46.71 1.2 47.81 0.4 47.81 0.4 48.07 1.2 48.07 1.2 49.17 0.4 49.17 0.4 49.43 1.2 49.43 1.2 50.53 0.4 50.53 0.4 50.79 1.2 50.79 1.2 51.89 0.4 51.89 0.4 52.83 1.2 52.83 1.2 53.93 0.4 53.93 0.4 54.19 1.2 54.19 1.2 55.29 0.4 55.29 0.4 55.55 1.2 55.55 1.2 56.65 0.4 56.65 0.4 56.91 1.2 56.91 1.2 58.01 0.4 58.01 0.4 58.95 1.2 58.95 1.2 60.05 0.4 60.05 0.4 60.31 1.2 60.31 1.2 61.41 0.4 61.41 0.4 61.67 1.2 61.67 1.2 62.77 0.4 62.77 0.4 63.03 1.2 63.03 1.2 64.13 0.4 64.13 0.4 64.39 1.2 64.39 1.2 65.49 0.4 65.49 0.4 66.43 1.2 66.43 1.2 67.53 0.4 67.53 0.4 67.79 1.2 67.79 1.2 68.89 0.4 68.89 0.4 69.15 1.2 69.15 1.2 70.25 0.4 70.25 0.4 70.51 1.2 70.51 1.2 71.61 0.4 71.61 0.4 71.87 1.2 71.87 1.2 72.97 0.4 72.97 0.4 73.23 1.2 73.23 1.2 74.33 0.4 74.33 0.4 74.59 1.2 74.59 1.2 75.69 0.4 75.69 0.4 76.63 1.2 76.63 1.2 77.73 0.4 77.73 0.4 77.99 1.2 77.99 1.2 79.09 0.4 79.09 0.4 79.35 1.2 79.35 1.2 80.45 0.4 80.45 0.4 80.71 1.2 80.71 1.2 81.81 0.4 81.81 0.4 82.75 1.2 82.75 1.2 83.85 0.4 83.85 0.4 86.64 26.16 86.64 26.16 97.52 ;
    LAYER met1 ;
      RECT 45.68 97.68 46.32 98.16 ;
      RECT 41.01 87.42 41.33 87.68 ;
      POLYGON 32.59 86.66 32.59 86.4 32.27 86.4 32.27 86.46 32.115 86.46 32.115 86.415 31.825 86.415 31.825 86.645 32.115 86.645 32.115 86.6 32.27 86.6 32.27 86.66 ;
      POLYGON 43.155 86.645 43.155 86.6 43.54 86.6 43.54 86.12 43.4 86.12 43.4 86.46 43.155 86.46 43.155 86.415 42.865 86.415 42.865 86.645 ;
      RECT 45.68 -0.24 46.32 0.24 ;
      POLYGON 46.32 97.64 46.32 97.4 91.72 97.4 91.72 95.72 91.24 95.72 91.24 94.68 91.72 94.68 91.72 93 91.24 93 91.24 91.96 91.72 91.96 91.72 90.28 91.24 90.28 91.24 89.24 91.72 89.24 91.72 87.56 91.24 87.56 91.24 86.52 91.72 86.52 91.72 84.84 91.24 84.84 91.24 83.8 91.72 83.8 91.72 82.12 91.24 82.12 91.24 81.08 91.72 81.08 91.72 79.4 91.24 79.4 91.24 78.36 91.72 78.36 91.72 76.68 91.24 76.68 91.24 75.64 91.72 75.64 91.72 73.96 91.24 73.96 91.24 72.92 91.72 72.92 91.72 71.24 91.24 71.24 91.24 70.2 91.72 70.2 91.72 68.52 91.24 68.52 91.24 67.48 91.72 67.48 91.72 65.8 91.24 65.8 91.24 64.76 91.72 64.76 91.72 63.08 91.24 63.08 91.24 62.04 91.72 62.04 91.72 60.36 91.24 60.36 91.24 59.32 91.72 59.32 91.72 57.64 91.24 57.64 91.24 56.6 91.72 56.6 91.72 54.92 91.24 54.92 91.24 53.88 91.72 53.88 91.72 52.2 91.24 52.2 91.24 51.16 91.72 51.16 91.72 49.48 91.24 49.48 91.24 48.44 91.72 48.44 91.72 46.76 91.24 46.76 91.24 45.72 91.72 45.72 91.72 44.04 91.24 44.04 91.24 43 91.72 43 91.72 41.32 91.24 41.32 91.24 40.28 91.72 40.28 91.72 38.6 91.24 38.6 91.24 37.56 91.72 37.56 91.72 35.88 91.24 35.88 91.24 34.84 91.72 34.84 91.72 33.16 91.24 33.16 91.24 32.12 91.72 32.12 91.72 30.44 91.24 30.44 91.24 29.4 91.72 29.4 91.72 27.72 91.24 27.72 91.24 26.68 91.72 26.68 91.72 25 91.24 25 91.24 23.96 91.72 23.96 91.72 22.28 91.24 22.28 91.24 21.24 91.72 21.24 91.72 19.56 91.24 19.56 91.24 18.52 91.72 18.52 91.72 16.84 91.24 16.84 91.24 15.8 91.72 15.8 91.72 14.12 91.24 14.12 91.24 13.08 91.72 13.08 91.72 11.4 91.24 11.4 91.24 10.36 91.72 10.36 91.72 8.68 91.24 8.68 91.24 7.64 91.72 7.64 91.72 5.96 91.24 5.96 91.24 4.92 91.72 4.92 91.72 3.24 91.24 3.24 91.24 2.2 91.72 2.2 91.72 0.52 46.32 0.52 46.32 0.28 45.68 0.28 45.68 0.52 0.28 0.52 0.28 2.2 0.76 2.2 0.76 3.24 0.28 3.24 0.28 4.92 0.76 4.92 0.76 5.96 0.28 5.96 0.28 7.64 0.76 7.64 0.76 8.68 0.28 8.68 0.28 10.36 0.76 10.36 0.76 11.4 0.28 11.4 0.28 13.08 0.76 13.08 0.76 14.12 0.28 14.12 0.28 15.8 0.76 15.8 0.76 16.84 0.28 16.84 0.28 18.52 0.76 18.52 0.76 19.56 0.28 19.56 0.28 21.24 0.76 21.24 0.76 22.28 0.28 22.28 0.28 23.96 0.76 23.96 0.76 25 0.28 25 0.28 26.68 0.76 26.68 0.76 27.72 0.28 27.72 0.28 29.4 0.76 29.4 0.76 30.44 0.28 30.44 0.28 32.12 0.76 32.12 0.76 33.16 0.28 33.16 0.28 34.84 0.76 34.84 0.76 35.88 0.28 35.88 0.28 37.56 0.76 37.56 0.76 38.6 0.28 38.6 0.28 40.28 0.76 40.28 0.76 41.32 0.28 41.32 0.28 43 0.76 43 0.76 44.04 0.28 44.04 0.28 45.72 0.76 45.72 0.76 46.76 0.28 46.76 0.28 48.44 0.76 48.44 0.76 49.48 0.28 49.48 0.28 51.16 0.76 51.16 0.76 52.2 0.28 52.2 0.28 53.88 0.76 53.88 0.76 54.92 0.28 54.92 0.28 56.6 0.76 56.6 0.76 57.64 0.28 57.64 0.28 59.32 0.76 59.32 0.76 60.36 0.28 60.36 0.28 62.04 0.76 62.04 0.76 63.08 0.28 63.08 0.28 64.76 0.76 64.76 0.76 65.8 0.28 65.8 0.28 67.48 0.76 67.48 0.76 68.52 0.28 68.52 0.28 70.2 0.76 70.2 0.76 71.24 0.28 71.24 0.28 72.92 0.76 72.92 0.76 73.96 0.28 73.96 0.28 75.64 0.76 75.64 0.76 76.68 0.28 76.68 0.28 78.36 0.76 78.36 0.76 79.4 0.28 79.4 0.28 81.08 0.76 81.08 0.76 82.12 0.28 82.12 0.28 83.8 0.76 83.8 0.76 84.84 0.28 84.84 0.28 86.52 45.68 86.52 45.68 87.56 26.04 87.56 26.04 89.24 26.52 89.24 26.52 90.28 26.04 90.28 26.04 91.96 26.52 91.96 26.52 93 26.04 93 26.04 94.68 26.52 94.68 26.52 95.72 26.04 95.72 26.04 97.4 45.68 97.4 45.68 97.64 ;
    LAYER met4 ;
      POLYGON 91.6 97.52 91.6 0.4 81.66 0.4 81.66 1 80.26 1 80.26 0.4 66.94 0.4 66.94 1 65.54 1 65.54 0.4 52.22 0.4 52.22 1 50.82 1 50.82 0.4 37.5 0.4 37.5 1 36.1 1 36.1 0.4 11.74 0.4 11.74 1 10.34 1 10.34 0.4 0.4 0.4 0.4 86.64 10.34 86.64 10.34 86.04 11.74 86.04 11.74 86.64 26.16 86.64 26.16 97.52 36.1 97.52 36.1 96.92 37.5 96.92 37.5 97.52 50.82 97.52 50.82 96.92 52.22 96.92 52.22 97.52 65.54 97.52 65.54 96.92 66.94 96.92 66.94 97.52 80.26 97.52 80.26 96.92 81.66 96.92 81.66 97.52 ;
    LAYER met5 ;
      POLYGON 90.4 96.32 90.4 77.32 87.2 77.32 87.2 70.92 90.4 70.92 90.4 56.92 87.2 56.92 87.2 50.52 90.4 50.52 90.4 36.52 87.2 36.52 87.2 30.12 90.4 30.12 90.4 16.12 87.2 16.12 87.2 9.72 90.4 9.72 90.4 1.6 1.6 1.6 1.6 9.72 4.8 9.72 4.8 16.12 1.6 16.12 1.6 30.12 4.8 30.12 4.8 36.52 1.6 36.52 1.6 50.52 4.8 50.52 4.8 56.92 1.6 56.92 1.6 70.92 4.8 70.92 4.8 77.32 1.6 77.32 1.6 85.44 27.36 85.44 27.36 96.32 ;
    LAYER li1 ;
      RECT 25.76 97.835 92 98.005 ;
      RECT 88.32 95.115 92 95.285 ;
      RECT 25.76 95.115 29.44 95.285 ;
      RECT 91.54 92.395 92 92.565 ;
      RECT 25.76 92.395 27.6 92.565 ;
      RECT 91.08 89.675 92 89.845 ;
      RECT 25.76 89.675 27.6 89.845 ;
      RECT 88.32 86.955 92 87.125 ;
      RECT 0 86.955 27.6 87.125 ;
      RECT 88.32 84.235 92 84.405 ;
      RECT 0 84.235 3.68 84.405 ;
      RECT 91.08 81.515 92 81.685 ;
      RECT 0 81.515 3.68 81.685 ;
      RECT 91.08 78.795 92 78.965 ;
      RECT 0 78.795 3.68 78.965 ;
      RECT 88.32 76.075 92 76.245 ;
      RECT 0 76.075 3.68 76.245 ;
      RECT 88.32 73.355 92 73.525 ;
      RECT 0 73.355 3.68 73.525 ;
      RECT 90.16 70.635 92 70.805 ;
      RECT 0 70.635 3.68 70.805 ;
      RECT 90.16 67.915 92 68.085 ;
      RECT 0 67.915 1.84 68.085 ;
      RECT 91.08 65.195 92 65.365 ;
      RECT 0 65.195 1.84 65.365 ;
      RECT 91.54 62.475 92 62.645 ;
      RECT 0 62.475 1.84 62.645 ;
      RECT 91.08 59.755 92 59.925 ;
      RECT 0 59.755 3.68 59.925 ;
      RECT 91.08 57.035 92 57.205 ;
      RECT 0 57.035 3.68 57.205 ;
      RECT 88.32 54.315 92 54.485 ;
      RECT 0 54.315 3.68 54.485 ;
      RECT 88.32 51.595 92 51.765 ;
      RECT 0 51.595 3.68 51.765 ;
      RECT 91.08 48.875 92 49.045 ;
      RECT 0 48.875 3.68 49.045 ;
      RECT 91.08 46.155 92 46.325 ;
      RECT 0 46.155 1.84 46.325 ;
      RECT 91.54 43.435 92 43.605 ;
      RECT 0 43.435 3.68 43.605 ;
      RECT 91.08 40.715 92 40.885 ;
      RECT 0 40.715 3.68 40.885 ;
      RECT 91.08 37.995 92 38.165 ;
      RECT 0 37.995 3.68 38.165 ;
      RECT 90.16 35.275 92 35.445 ;
      RECT 0 35.275 3.68 35.445 ;
      RECT 90.16 32.555 92 32.725 ;
      RECT 0 32.555 3.68 32.725 ;
      RECT 91.54 29.835 92 30.005 ;
      RECT 0 29.835 3.68 30.005 ;
      RECT 91.08 27.115 92 27.285 ;
      RECT 0 27.115 1.84 27.285 ;
      RECT 91.08 24.395 92 24.565 ;
      RECT 0 24.395 3.68 24.565 ;
      RECT 91.08 21.675 92 21.845 ;
      RECT 0 21.675 3.68 21.845 ;
      RECT 91.08 18.955 92 19.125 ;
      RECT 0 18.955 3.68 19.125 ;
      RECT 91.54 16.235 92 16.405 ;
      RECT 0 16.235 3.68 16.405 ;
      RECT 91.54 13.515 92 13.685 ;
      RECT 0 13.515 3.68 13.685 ;
      RECT 88.32 10.795 92 10.965 ;
      RECT 0 10.795 3.68 10.965 ;
      RECT 88.32 8.075 92 8.245 ;
      RECT 0 8.075 3.68 8.245 ;
      RECT 88.32 5.355 92 5.525 ;
      RECT 0 5.355 3.68 5.525 ;
      RECT 88.32 2.635 92 2.805 ;
      RECT 0 2.635 3.68 2.805 ;
      RECT 0 -0.085 92 0.085 ;
      POLYGON 91.83 97.75 91.83 0.17 0.17 0.17 0.17 86.87 25.93 86.87 25.93 97.75 ;
    LAYER mcon ;
      RECT 41.085 87.465 41.255 87.635 ;
      RECT 42.925 86.445 43.095 86.615 ;
      RECT 31.885 86.445 32.055 86.615 ;
    LAYER via ;
      RECT 80.885 97.845 81.035 97.995 ;
      RECT 51.445 97.845 51.595 97.995 ;
      RECT 41.095 87.475 41.245 87.625 ;
      RECT 10.965 86.965 11.115 87.115 ;
      RECT 32.355 86.455 32.505 86.605 ;
      RECT 80.885 -0.075 81.035 0.075 ;
      RECT 51.445 -0.075 51.595 0.075 ;
      RECT 10.965 -0.075 11.115 0.075 ;
    LAYER via2 ;
      RECT 80.86 97.82 81.06 98.02 ;
      RECT 51.42 97.82 51.62 98.02 ;
      RECT 10.94 86.94 11.14 87.14 ;
      RECT 1.05 68.24 1.25 68.44 ;
      RECT 1.05 54.64 1.25 54.84 ;
      RECT 80.86 -0.1 81.06 0.1 ;
      RECT 51.42 -0.1 51.62 0.1 ;
      RECT 10.94 -0.1 11.14 0.1 ;
    LAYER via3 ;
      RECT 80.86 97.82 81.06 98.02 ;
      RECT 51.42 97.82 51.62 98.02 ;
      RECT 10.94 86.94 11.14 87.14 ;
      RECT 80.86 -0.1 81.06 0.1 ;
      RECT 51.42 -0.1 51.62 0.1 ;
      RECT 10.94 -0.1 11.14 0.1 ;
    LAYER OVERLAP ;
      POLYGON 0 0 0 87.04 25.76 87.04 25.76 97.92 92 97.92 92 0 ;
  END
END sb_2__0_

END LIBRARY
