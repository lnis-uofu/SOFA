VERSION 5.7 ;
BUSBITCHARS "[]" ;

UNITS
  DATABASE MICRONS 1000 ;
END UNITS

MANUFACTURINGGRID 0.005 ;

LAYER li1
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.46 ;
  WIDTH 0.17 ;
END li1

LAYER mcon
  TYPE CUT ;
END mcon

LAYER met1
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.34 ;
  WIDTH 0.14 ;
END met1

LAYER via
  TYPE CUT ;
END via

LAYER met2
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.46 ;
  WIDTH 0.14 ;
END met2

LAYER via2
  TYPE CUT ;
END via2

LAYER met3
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.68 ;
  WIDTH 0.3 ;
END met3

LAYER via3
  TYPE CUT ;
END via3

LAYER met4
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.92 ;
  WIDTH 0.3 ;
END met4

LAYER via4
  TYPE CUT ;
END via4

LAYER met5
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 3.4 ;
  WIDTH 1.6 ;
END met5

LAYER nwell
  TYPE MASTERSLICE ;
END nwell

LAYER pwell
  TYPE MASTERSLICE ;
END pwell

LAYER OVERLAP
  TYPE OVERLAP ;
END OVERLAP

VIA L1M1_PR
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.145 -0.115 0.145 0.115 ;
END L1M1_PR

VIA L1M1_PR_R
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.115 -0.145 0.115 0.145 ;
END L1M1_PR_R

VIA L1M1_PR_M
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.115 -0.145 0.115 0.145 ;
END L1M1_PR_M

VIA L1M1_PR_MR
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.145 -0.115 0.145 0.115 ;
END L1M1_PR_MR

VIA L1M1_PR_C
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.145 -0.145 0.145 0.145 ;
END L1M1_PR_C

VIA M1M2_PR
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR

VIA M1M2_PR_Enc
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_Enc

VIA M1M2_PR_R
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_R

VIA M1M2_PR_R_Enc
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR_R_Enc

VIA M1M2_PR_M
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_M

VIA M1M2_PR_M_Enc
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR_M_Enc

VIA M1M2_PR_MR
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR_MR

VIA M1M2_PR_MR_Enc
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_MR_Enc

VIA M1M2_PR_C
  LAYER met1 ;
    RECT -0.16 -0.16 0.16 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.16 0.16 0.16 ;
END M1M2_PR_C

VIA M2M3_PR
  LAYER met2 ;
    RECT -0.14 -0.185 0.14 0.185 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR

VIA M2M3_PR_R
  LAYER met2 ;
    RECT -0.185 -0.14 0.185 0.14 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_R

VIA M2M3_PR_M
  LAYER met2 ;
    RECT -0.14 -0.185 0.14 0.185 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_M

VIA M2M3_PR_MR
  LAYER met2 ;
    RECT -0.185 -0.14 0.185 0.14 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_MR

VIA M2M3_PR_C
  LAYER met2 ;
    RECT -0.185 -0.185 0.185 0.185 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_C

VIA M3M4_PR
  LAYER met3 ;
    RECT -0.19 -0.16 0.19 0.16 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR

VIA M3M4_PR_R
  LAYER met3 ;
    RECT -0.16 -0.19 0.16 0.19 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_R

VIA M3M4_PR_M
  LAYER met3 ;
    RECT -0.19 -0.16 0.19 0.16 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_M

VIA M3M4_PR_MR
  LAYER met3 ;
    RECT -0.16 -0.19 0.16 0.19 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_MR

VIA M3M4_PR_C
  LAYER met3 ;
    RECT -0.19 -0.19 0.19 0.19 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_C

VIA M4M5_PR
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR

VIA M4M5_PR_R
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_R

VIA M4M5_PR_M
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_M

VIA M4M5_PR_MR
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_MR

VIA M4M5_PR_C
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_C

SITE unit
  CLASS CORE ;
  SYMMETRY Y ;
  SIZE 0.46 BY 2.72 ;
END unit

SITE unithddbl
  CLASS CORE ;
  SIZE 0.46 BY 5.44 ;
END unithddbl

MACRO sb_2__0_
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  SIZE 95.68 BY 97.92 ;
  SYMMETRY X Y ;
  PIN prog_clk[0]
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER met3 ;
        RECT 0 13.45 1.38 13.75 ;
    END
  END prog_clk[0]
  PIN chany_top_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.11 96.56 61.25 97.92 ;
    END
  END chany_top_in[0]
  PIN chany_top_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 63.33 96.56 63.63 97.92 ;
    END
  END chany_top_in[1]
  PIN chany_top_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 61.49 96.56 61.79 97.92 ;
    END
  END chany_top_in[2]
  PIN chany_top_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.91 96.56 52.05 97.92 ;
    END
  END chany_top_in[3]
  PIN chany_top_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.43 96.56 57.57 97.92 ;
    END
  END chany_top_in[4]
  PIN chany_top_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.03 96.56 62.17 97.92 ;
    END
  END chany_top_in[5]
  PIN chany_top_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.01 96.56 68.15 97.92 ;
    END
  END chany_top_in[6]
  PIN chany_top_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.15 96.56 49.29 97.92 ;
    END
  END chany_top_in[7]
  PIN chany_top_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.17 96.56 66.31 97.92 ;
    END
  END chany_top_in[8]
  PIN chany_top_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 45.85 96.56 46.15 97.92 ;
    END
  END chany_top_in[9]
  PIN chany_top_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 44.01 96.56 44.31 97.92 ;
    END
  END chany_top_in[10]
  PIN chany_top_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.13 96.56 78.27 97.92 ;
    END
  END chany_top_in[11]
  PIN chany_top_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.35 96.56 58.49 97.92 ;
    END
  END chany_top_in[12]
  PIN chany_top_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.27 96.56 59.41 97.92 ;
    END
  END chany_top_in[13]
  PIN chany_top_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.77 96.56 70.91 97.92 ;
    END
  END chany_top_in[14]
  PIN chany_top_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.33 96.56 64.47 97.92 ;
    END
  END chany_top_in[15]
  PIN chany_top_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.89 96.56 81.03 97.92 ;
    END
  END chany_top_in[16]
  PIN chany_top_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.97 96.56 80.11 97.92 ;
    END
  END chany_top_in[17]
  PIN chany_top_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.19 96.56 60.33 97.92 ;
    END
  END chany_top_in[18]
  PIN chany_top_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.05 96.56 79.19 97.92 ;
    END
  END chany_top_in[19]
  PIN top_left_grid_pin_42_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.87 85.68 18.01 87.04 ;
    END
  END top_left_grid_pin_42_[0]
  PIN top_left_grid_pin_43_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.81 85.68 12.95 87.04 ;
    END
  END top_left_grid_pin_43_[0]
  PIN top_left_grid_pin_44_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.21 85.68 8.35 87.04 ;
    END
  END top_left_grid_pin_44_[0]
  PIN top_left_grid_pin_45_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.89 85.68 12.03 87.04 ;
    END
  END top_left_grid_pin_45_[0]
  PIN top_left_grid_pin_46_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.37 85.68 6.51 87.04 ;
    END
  END top_left_grid_pin_46_[0]
  PIN top_left_grid_pin_47_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.97 85.68 11.11 87.04 ;
    END
  END top_left_grid_pin_47_[0]
  PIN top_left_grid_pin_48_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.29 85.68 7.43 87.04 ;
    END
  END top_left_grid_pin_48_[0]
  PIN top_left_grid_pin_49_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.45 85.68 5.59 87.04 ;
    END
  END top_left_grid_pin_49_[0]
  PIN top_right_grid_pin_1_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.55 96.56 44.69 97.92 ;
    END
  END top_right_grid_pin_1_[0]
  PIN chanx_left_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 76.69 1.38 76.99 ;
    END
  END chanx_left_in[0]
  PIN chanx_left_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 63.77 1.38 64.07 ;
    END
  END chanx_left_in[1]
  PIN chanx_left_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 58.33 1.38 58.63 ;
    END
  END chanx_left_in[2]
  PIN chanx_left_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 73.97 1.38 74.27 ;
    END
  END chanx_left_in[3]
  PIN chanx_left_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 23.65 1.38 23.95 ;
    END
  END chanx_left_in[4]
  PIN chanx_left_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 36.57 1.38 36.87 ;
    END
  END chanx_left_in[5]
  PIN chanx_left_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 55.61 1.38 55.91 ;
    END
  END chanx_left_in[6]
  PIN chanx_left_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 29.77 1.38 30.07 ;
    END
  END chanx_left_in[7]
  PIN chanx_left_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 26.37 1.38 26.67 ;
    END
  END chanx_left_in[8]
  PIN chanx_left_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 10.05 1.38 10.35 ;
    END
  END chanx_left_in[9]
  PIN chanx_left_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 50.17 1.38 50.47 ;
    END
  END chanx_left_in[10]
  PIN chanx_left_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 33.85 1.38 34.15 ;
    END
  END chanx_left_in[11]
  PIN chanx_left_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 62.41 1.38 62.71 ;
    END
  END chanx_left_in[12]
  PIN chanx_left_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 72.61 1.38 72.91 ;
    END
  END chanx_left_in[13]
  PIN chanx_left_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 18.89 1.38 19.19 ;
    END
  END chanx_left_in[14]
  PIN chanx_left_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 39.29 1.38 39.59 ;
    END
  END chanx_left_in[15]
  PIN chanx_left_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 43.37 1.38 43.67 ;
    END
  END chanx_left_in[16]
  PIN chanx_left_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 32.49 1.38 32.79 ;
    END
  END chanx_left_in[17]
  PIN chanx_left_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 31.13 1.38 31.43 ;
    END
  END chanx_left_in[18]
  PIN chanx_left_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 17.53 1.38 17.83 ;
    END
  END chanx_left_in[19]
  PIN left_bottom_grid_pin_1_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 54.25 1.38 54.55 ;
    END
  END left_bottom_grid_pin_1_[0]
  PIN left_bottom_grid_pin_3_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 51.53 1.38 51.83 ;
    END
  END left_bottom_grid_pin_3_[0]
  PIN left_bottom_grid_pin_5_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 40.65 1.38 40.95 ;
    END
  END left_bottom_grid_pin_5_[0]
  PIN left_bottom_grid_pin_7_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 67.85 1.38 68.15 ;
    END
  END left_bottom_grid_pin_7_[0]
  PIN left_bottom_grid_pin_9_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 42.01 1.38 42.31 ;
    END
  END left_bottom_grid_pin_9_[0]
  PIN left_bottom_grid_pin_11_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 48.13 1.38 48.43 ;
    END
  END left_bottom_grid_pin_11_[0]
  PIN ccff_head[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.35 96.56 35.49 97.92 ;
    END
  END ccff_head[0]
  PIN chany_top_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.29 96.56 53.43 97.92 ;
    END
  END chany_top_out[0]
  PIN chany_top_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.99 96.56 51.13 97.92 ;
    END
  END chany_top_out[1]
  PIN chany_top_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.13 96.56 55.27 97.92 ;
    END
  END chany_top_out[2]
  PIN chany_top_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.03 96.56 39.17 97.92 ;
    END
  END chany_top_out[3]
  PIN chany_top_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.79 96.56 41.93 97.92 ;
    END
  END chany_top_out[4]
  PIN chany_top_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.95 96.56 40.09 97.92 ;
    END
  END chany_top_out[5]
  PIN chany_top_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.21 96.56 77.35 97.92 ;
    END
  END chany_top_out[6]
  PIN chany_top_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.11 96.56 38.25 97.92 ;
    END
  END chany_top_out[7]
  PIN chany_top_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.25 96.56 65.39 97.92 ;
    END
  END chany_top_out[8]
  PIN chany_top_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.41 96.56 63.55 97.92 ;
    END
  END chany_top_out[9]
  PIN chany_top_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.23 96.56 48.37 97.92 ;
    END
  END chany_top_out[10]
  PIN chany_top_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.19 96.56 37.33 97.92 ;
    END
  END chany_top_out[11]
  PIN chany_top_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.07 96.56 50.21 97.92 ;
    END
  END chany_top_out[12]
  PIN chany_top_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.31 96.56 47.45 97.92 ;
    END
  END chany_top_out[13]
  PIN chany_top_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.09 96.56 67.23 97.92 ;
    END
  END chany_top_out[14]
  PIN chany_top_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.71 96.56 42.85 97.92 ;
    END
  END chany_top_out[15]
  PIN chany_top_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.63 96.56 43.77 97.92 ;
    END
  END chany_top_out[16]
  PIN chany_top_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.87 96.56 41.01 97.92 ;
    END
  END chany_top_out[17]
  PIN chany_top_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.39 96.56 46.53 97.92 ;
    END
  END chany_top_out[18]
  PIN chany_top_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.47 96.56 45.61 97.92 ;
    END
  END chany_top_out[19]
  PIN chanx_left_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 44.73 1.38 45.03 ;
    END
  END chanx_left_out[0]
  PIN chanx_left_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 56.97 1.38 57.27 ;
    END
  END chanx_left_out[1]
  PIN chanx_left_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 59.69 1.38 59.99 ;
    END
  END chanx_left_out[2]
  PIN chanx_left_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 75.33 1.38 75.63 ;
    END
  END chanx_left_out[3]
  PIN chanx_left_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 20.25 1.38 20.55 ;
    END
  END chanx_left_out[4]
  PIN chanx_left_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 61.05 1.38 61.35 ;
    END
  END chanx_left_out[5]
  PIN chanx_left_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 78.73 1.38 79.03 ;
    END
  END chanx_left_out[6]
  PIN chanx_left_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 8.69 1.38 8.99 ;
    END
  END chanx_left_out[7]
  PIN chanx_left_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 35.21 1.38 35.51 ;
    END
  END chanx_left_out[8]
  PIN chanx_left_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 52.89 1.38 53.19 ;
    END
  END chanx_left_out[9]
  PIN chanx_left_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 46.09 1.38 46.39 ;
    END
  END chanx_left_out[10]
  PIN chanx_left_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 82.81 1.38 83.11 ;
    END
  END chanx_left_out[11]
  PIN chanx_left_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 65.13 1.38 65.43 ;
    END
  END chanx_left_out[12]
  PIN chanx_left_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 16.17 1.38 16.47 ;
    END
  END chanx_left_out[13]
  PIN chanx_left_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 28.41 1.38 28.71 ;
    END
  END chanx_left_out[14]
  PIN chanx_left_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 37.93 1.38 38.23 ;
    END
  END chanx_left_out[15]
  PIN chanx_left_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 25.01 1.38 25.31 ;
    END
  END chanx_left_out[16]
  PIN chanx_left_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 69.21 1.38 69.51 ;
    END
  END chanx_left_out[17]
  PIN chanx_left_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 66.49 1.38 66.79 ;
    END
  END chanx_left_out[18]
  PIN chanx_left_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 71.25 1.38 71.55 ;
    END
  END chanx_left_out[19]
  PIN ccff_tail[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 11.41 1.38 11.71 ;
    END
  END ccff_tail[0]
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 0.48 2.96 ;
        RECT 95.2 2.48 95.68 2.96 ;
        RECT 0 7.92 0.48 8.4 ;
        RECT 95.2 7.92 95.68 8.4 ;
        RECT 0 13.36 0.48 13.84 ;
        RECT 95.2 13.36 95.68 13.84 ;
        RECT 0 18.8 0.48 19.28 ;
        RECT 95.2 18.8 95.68 19.28 ;
        RECT 0 24.24 0.48 24.72 ;
        RECT 95.2 24.24 95.68 24.72 ;
        RECT 0 29.68 0.48 30.16 ;
        RECT 95.2 29.68 95.68 30.16 ;
        RECT 0 35.12 0.48 35.6 ;
        RECT 95.2 35.12 95.68 35.6 ;
        RECT 0 40.56 0.48 41.04 ;
        RECT 95.2 40.56 95.68 41.04 ;
        RECT 0 46 0.48 46.48 ;
        RECT 95.2 46 95.68 46.48 ;
        RECT 0 51.44 0.48 51.92 ;
        RECT 95.2 51.44 95.68 51.92 ;
        RECT 0 56.88 0.48 57.36 ;
        RECT 95.2 56.88 95.68 57.36 ;
        RECT 0 62.32 0.48 62.8 ;
        RECT 95.2 62.32 95.68 62.8 ;
        RECT 0 67.76 0.48 68.24 ;
        RECT 95.2 67.76 95.68 68.24 ;
        RECT 0 73.2 0.48 73.68 ;
        RECT 95.2 73.2 95.68 73.68 ;
        RECT 0 78.64 0.48 79.12 ;
        RECT 95.2 78.64 95.68 79.12 ;
        RECT 0 84.08 0.48 84.56 ;
        RECT 95.2 84.08 95.68 84.56 ;
        RECT 27.6 89.52 28.08 90 ;
        RECT 95.2 89.52 95.68 90 ;
        RECT 27.6 94.96 28.08 95.44 ;
        RECT 95.2 94.96 95.68 95.44 ;
      LAYER met4 ;
        RECT 39.26 0 39.86 0.6 ;
        RECT 68.7 0 69.3 0.6 ;
        RECT 39.26 97.32 39.86 97.92 ;
        RECT 68.7 97.32 69.3 97.92 ;
      LAYER met5 ;
        RECT 0 11.32 3.2 14.52 ;
        RECT 92.48 11.32 95.68 14.52 ;
        RECT 0 52.12 3.2 55.32 ;
        RECT 92.48 52.12 95.68 55.32 ;
    END
  END VDD
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 0 95.68 0.24 ;
        RECT 0 5.2 0.48 5.68 ;
        RECT 95.2 5.2 95.68 5.68 ;
        RECT 0 10.64 0.48 11.12 ;
        RECT 95.2 10.64 95.68 11.12 ;
        RECT 0 16.08 0.48 16.56 ;
        RECT 95.2 16.08 95.68 16.56 ;
        RECT 0 21.52 0.48 22 ;
        RECT 95.2 21.52 95.68 22 ;
        RECT 0 26.96 0.48 27.44 ;
        RECT 95.2 26.96 95.68 27.44 ;
        RECT 0 32.4 0.48 32.88 ;
        RECT 95.2 32.4 95.68 32.88 ;
        RECT 0 37.84 0.48 38.32 ;
        RECT 95.2 37.84 95.68 38.32 ;
        RECT 0 43.28 0.48 43.76 ;
        RECT 95.2 43.28 95.68 43.76 ;
        RECT 0 48.72 0.48 49.2 ;
        RECT 95.2 48.72 95.68 49.2 ;
        RECT 0 54.16 0.48 54.64 ;
        RECT 95.2 54.16 95.68 54.64 ;
        RECT 0 59.6 0.48 60.08 ;
        RECT 95.2 59.6 95.68 60.08 ;
        RECT 0 65.04 0.48 65.52 ;
        RECT 95.2 65.04 95.68 65.52 ;
        RECT 0 70.48 0.48 70.96 ;
        RECT 95.2 70.48 95.68 70.96 ;
        RECT 0 75.92 0.48 76.4 ;
        RECT 95.2 75.92 95.68 76.4 ;
        RECT 0 81.36 0.48 81.84 ;
        RECT 95.2 81.36 95.68 81.84 ;
        RECT 0 86.8 95.68 87.28 ;
        RECT 27.6 92.24 28.08 92.72 ;
        RECT 95.2 92.24 95.68 92.72 ;
        RECT 27.6 97.68 95.68 97.92 ;
      LAYER met4 ;
        RECT 9.82 0 10.42 0.6 ;
        RECT 53.98 0 54.58 0.6 ;
        RECT 83.42 0 84.02 0.6 ;
        RECT 9.82 86.44 10.42 87.04 ;
        RECT 53.98 97.32 54.58 97.92 ;
        RECT 83.42 97.32 84.02 97.92 ;
      LAYER met5 ;
        RECT 0 31.72 3.2 34.92 ;
        RECT 92.48 31.72 95.68 34.92 ;
        RECT 0 72.52 3.2 75.72 ;
        RECT 92.48 72.52 95.68 75.72 ;
    END
  END VSS
  OBS
    LAYER li1 ;
      RECT 27.6 97.835 95.68 98.005 ;
      RECT 92 95.115 95.68 95.285 ;
      RECT 27.6 95.115 31.28 95.285 ;
      RECT 92 92.395 95.68 92.565 ;
      RECT 27.6 92.395 31.28 92.565 ;
      RECT 95.22 89.675 95.68 89.845 ;
      RECT 27.6 89.675 31.28 89.845 ;
      RECT 95.22 86.955 95.68 87.125 ;
      RECT 0 86.955 29.44 87.125 ;
      RECT 95.22 84.235 95.68 84.405 ;
      RECT 0 84.235 3.68 84.405 ;
      RECT 94.76 81.515 95.68 81.685 ;
      RECT 0 81.515 1.84 81.685 ;
      RECT 94.76 78.795 95.68 78.965 ;
      RECT 0 78.795 1.84 78.965 ;
      RECT 94.76 76.075 95.68 76.245 ;
      RECT 0 76.075 1.84 76.245 ;
      RECT 94.76 73.355 95.68 73.525 ;
      RECT 0 73.355 1.84 73.525 ;
      RECT 95.22 70.635 95.68 70.805 ;
      RECT 0 70.635 1.84 70.805 ;
      RECT 94.76 67.915 95.68 68.085 ;
      RECT 0 67.915 1.84 68.085 ;
      RECT 94.76 65.195 95.68 65.365 ;
      RECT 0 65.195 1.84 65.365 ;
      RECT 95.22 62.475 95.68 62.645 ;
      RECT 0 62.475 1.84 62.645 ;
      RECT 92 59.755 95.68 59.925 ;
      RECT 0 59.755 1.84 59.925 ;
      RECT 92 57.035 95.68 57.205 ;
      RECT 0 57.035 1.84 57.205 ;
      RECT 93.84 54.315 95.68 54.485 ;
      RECT 0 54.315 3.68 54.485 ;
      RECT 95.22 51.595 95.68 51.765 ;
      RECT 0 51.595 3.68 51.765 ;
      RECT 95.22 48.875 95.68 49.045 ;
      RECT 0 48.875 1.84 49.045 ;
      RECT 92 46.155 95.68 46.325 ;
      RECT 0 46.155 1.84 46.325 ;
      RECT 92 43.435 95.68 43.605 ;
      RECT 0 43.435 1.84 43.605 ;
      RECT 93.84 40.715 95.68 40.885 ;
      RECT 0 40.715 1.84 40.885 ;
      RECT 93.84 37.995 95.68 38.165 ;
      RECT 0 37.995 1.84 38.165 ;
      RECT 95.22 35.275 95.68 35.445 ;
      RECT 0 35.275 1.84 35.445 ;
      RECT 95.22 32.555 95.68 32.725 ;
      RECT 0 32.555 1.84 32.725 ;
      RECT 95.22 29.835 95.68 30.005 ;
      RECT 0 29.835 1.84 30.005 ;
      RECT 95.22 27.115 95.68 27.285 ;
      RECT 0 27.115 1.84 27.285 ;
      RECT 95.22 24.395 95.68 24.565 ;
      RECT 0 24.395 1.84 24.565 ;
      RECT 95.22 21.675 95.68 21.845 ;
      RECT 0 21.675 1.84 21.845 ;
      RECT 95.22 18.955 95.68 19.125 ;
      RECT 0 18.955 1.84 19.125 ;
      RECT 95.22 16.235 95.68 16.405 ;
      RECT 0 16.235 1.84 16.405 ;
      RECT 95.22 13.515 95.68 13.685 ;
      RECT 0 13.515 1.84 13.685 ;
      RECT 95.22 10.795 95.68 10.965 ;
      RECT 0 10.795 1.84 10.965 ;
      RECT 95.22 8.075 95.68 8.245 ;
      RECT 0 8.075 3.68 8.245 ;
      RECT 95.22 5.355 95.68 5.525 ;
      RECT 0 5.355 3.68 5.525 ;
      RECT 95.22 2.635 95.68 2.805 ;
      RECT 0 2.635 3.68 2.805 ;
      RECT 0 -0.085 95.68 0.085 ;
    LAYER met3 ;
      POLYGON 83.885 98.085 83.885 98.08 84.1 98.08 84.1 97.76 83.885 97.76 83.885 97.755 83.555 97.755 83.555 97.76 83.34 97.76 83.34 98.08 83.555 98.08 83.555 98.085 ;
      POLYGON 54.445 98.085 54.445 98.08 54.66 98.08 54.66 97.76 54.445 97.76 54.445 97.755 54.115 97.755 54.115 97.76 53.9 97.76 53.9 98.08 54.115 98.08 54.115 98.085 ;
      POLYGON 10.285 87.205 10.285 87.2 10.5 87.2 10.5 86.88 10.285 86.88 10.285 86.875 9.955 86.875 9.955 86.88 9.74 86.88 9.74 87.2 9.955 87.2 9.955 87.205 ;
      POLYGON 11.65 66.11 11.65 65.81 1.99 65.81 1.99 65.13 1.78 65.13 1.78 65.83 1.69 65.83 1.69 66.11 ;
      POLYGON 7.51 59.31 7.51 59.01 1.78 59.01 1.78 59.03 1.23 59.03 1.23 59.31 ;
      POLYGON 1.99 45.03 1.99 44.35 6.59 44.35 6.59 44.05 1.69 44.05 1.69 44.33 1.78 44.33 1.78 45.03 ;
      POLYGON 1.99 39.59 1.99 38.91 21.77 38.91 21.77 38.61 1.69 38.61 1.69 38.89 1.78 38.89 1.78 39.59 ;
      POLYGON 2.005 28.045 2.005 28.03 15.79 28.03 15.79 27.73 2.005 27.73 2.005 27.715 1.675 27.715 1.675 28.045 ;
      POLYGON 6.59 25.99 6.59 25.69 1.99 25.69 1.99 25.01 1.78 25.01 1.78 25.71 1.69 25.71 1.69 25.99 ;
      POLYGON 83.885 0.165 83.885 0.16 84.1 0.16 84.1 -0.16 83.885 -0.16 83.885 -0.165 83.555 -0.165 83.555 -0.16 83.34 -0.16 83.34 0.16 83.555 0.16 83.555 0.165 ;
      POLYGON 54.445 0.165 54.445 0.16 54.66 0.16 54.66 -0.16 54.445 -0.16 54.445 -0.165 54.115 -0.165 54.115 -0.16 53.9 -0.16 53.9 0.16 54.115 0.16 54.115 0.165 ;
      POLYGON 10.285 0.165 10.285 0.16 10.5 0.16 10.5 -0.16 10.285 -0.16 10.285 -0.165 9.955 -0.165 9.955 -0.16 9.74 -0.16 9.74 0.16 9.955 0.16 9.955 0.165 ;
      POLYGON 95.28 97.52 95.28 0.4 0.4 0.4 0.4 8.29 1.78 8.29 1.78 9.39 0.4 9.39 0.4 9.65 1.78 9.65 1.78 10.75 0.4 10.75 0.4 11.01 1.78 11.01 1.78 12.11 0.4 12.11 0.4 13.05 1.78 13.05 1.78 14.15 0.4 14.15 0.4 15.77 1.78 15.77 1.78 16.87 0.4 16.87 0.4 17.13 1.78 17.13 1.78 18.23 0.4 18.23 0.4 18.49 1.78 18.49 1.78 19.59 0.4 19.59 0.4 19.85 1.78 19.85 1.78 20.95 0.4 20.95 0.4 23.25 1.78 23.25 1.78 24.35 0.4 24.35 0.4 24.61 1.78 24.61 1.78 25.71 0.4 25.71 0.4 25.97 1.78 25.97 1.78 27.07 0.4 27.07 0.4 28.01 1.78 28.01 1.78 29.11 0.4 29.11 0.4 29.37 1.78 29.37 1.78 30.47 0.4 30.47 0.4 30.73 1.78 30.73 1.78 31.83 0.4 31.83 0.4 32.09 1.78 32.09 1.78 33.19 0.4 33.19 0.4 33.45 1.78 33.45 1.78 34.55 0.4 34.55 0.4 34.81 1.78 34.81 1.78 35.91 0.4 35.91 0.4 36.17 1.78 36.17 1.78 37.27 0.4 37.27 0.4 37.53 1.78 37.53 1.78 38.63 0.4 38.63 0.4 38.89 1.78 38.89 1.78 39.99 0.4 39.99 0.4 40.25 1.78 40.25 1.78 41.35 0.4 41.35 0.4 41.61 1.78 41.61 1.78 42.71 0.4 42.71 0.4 42.97 1.78 42.97 1.78 44.07 0.4 44.07 0.4 44.33 1.78 44.33 1.78 45.43 0.4 45.43 0.4 45.69 1.78 45.69 1.78 46.79 0.4 46.79 0.4 47.73 1.78 47.73 1.78 48.83 0.4 48.83 0.4 49.77 1.78 49.77 1.78 50.87 0.4 50.87 0.4 51.13 1.78 51.13 1.78 52.23 0.4 52.23 0.4 52.49 1.78 52.49 1.78 53.59 0.4 53.59 0.4 53.85 1.78 53.85 1.78 54.95 0.4 54.95 0.4 55.21 1.78 55.21 1.78 56.31 0.4 56.31 0.4 56.57 1.78 56.57 1.78 57.67 0.4 57.67 0.4 57.93 1.78 57.93 1.78 59.03 0.4 59.03 0.4 59.29 1.78 59.29 1.78 60.39 0.4 60.39 0.4 60.65 1.78 60.65 1.78 61.75 0.4 61.75 0.4 62.01 1.78 62.01 1.78 63.11 0.4 63.11 0.4 63.37 1.78 63.37 1.78 64.47 0.4 64.47 0.4 64.73 1.78 64.73 1.78 65.83 0.4 65.83 0.4 66.09 1.78 66.09 1.78 67.19 0.4 67.19 0.4 67.45 1.78 67.45 1.78 68.55 0.4 68.55 0.4 68.81 1.78 68.81 1.78 69.91 0.4 69.91 0.4 70.85 1.78 70.85 1.78 71.95 0.4 71.95 0.4 72.21 1.78 72.21 1.78 73.31 0.4 73.31 0.4 73.57 1.78 73.57 1.78 74.67 0.4 74.67 0.4 74.93 1.78 74.93 1.78 76.03 0.4 76.03 0.4 76.29 1.78 76.29 1.78 77.39 0.4 77.39 0.4 78.33 1.78 78.33 1.78 79.43 0.4 79.43 0.4 82.41 1.78 82.41 1.78 83.51 0.4 83.51 0.4 86.64 28 86.64 28 97.52 ;
    LAYER met2 ;
      RECT 83.58 97.735 83.86 98.105 ;
      RECT 54.14 97.735 54.42 98.105 ;
      RECT 68.41 96.06 68.67 96.38 ;
      RECT 49.55 96.06 49.81 96.38 ;
      RECT 9.98 86.855 10.26 87.225 ;
      RECT 83.58 -0.185 83.86 0.185 ;
      RECT 54.14 -0.185 54.42 0.185 ;
      RECT 9.98 -0.185 10.26 0.185 ;
      POLYGON 95.4 97.64 95.4 0.28 0.28 0.28 0.28 86.76 5.17 86.76 5.17 85.4 5.87 85.4 5.87 86.76 6.09 86.76 6.09 85.4 6.79 85.4 6.79 86.76 7.01 86.76 7.01 85.4 7.71 85.4 7.71 86.76 7.93 86.76 7.93 85.4 8.63 85.4 8.63 86.76 10.69 86.76 10.69 85.4 11.39 85.4 11.39 86.76 11.61 86.76 11.61 85.4 12.31 85.4 12.31 86.76 12.53 86.76 12.53 85.4 13.23 85.4 13.23 86.76 17.59 86.76 17.59 85.4 18.29 85.4 18.29 86.76 27.88 86.76 27.88 97.64 35.07 97.64 35.07 96.28 35.77 96.28 35.77 97.64 36.91 97.64 36.91 96.28 37.61 96.28 37.61 97.64 37.83 97.64 37.83 96.28 38.53 96.28 38.53 97.64 38.75 97.64 38.75 96.28 39.45 96.28 39.45 97.64 39.67 97.64 39.67 96.28 40.37 96.28 40.37 97.64 40.59 97.64 40.59 96.28 41.29 96.28 41.29 97.64 41.51 97.64 41.51 96.28 42.21 96.28 42.21 97.64 42.43 97.64 42.43 96.28 43.13 96.28 43.13 97.64 43.35 97.64 43.35 96.28 44.05 96.28 44.05 97.64 44.27 97.64 44.27 96.28 44.97 96.28 44.97 97.64 45.19 97.64 45.19 96.28 45.89 96.28 45.89 97.64 46.11 97.64 46.11 96.28 46.81 96.28 46.81 97.64 47.03 97.64 47.03 96.28 47.73 96.28 47.73 97.64 47.95 97.64 47.95 96.28 48.65 96.28 48.65 97.64 48.87 97.64 48.87 96.28 49.57 96.28 49.57 97.64 49.79 97.64 49.79 96.28 50.49 96.28 50.49 97.64 50.71 97.64 50.71 96.28 51.41 96.28 51.41 97.64 51.63 97.64 51.63 96.28 52.33 96.28 52.33 97.64 53.01 97.64 53.01 96.28 53.71 96.28 53.71 97.64 54.85 97.64 54.85 96.28 55.55 96.28 55.55 97.64 57.15 97.64 57.15 96.28 57.85 96.28 57.85 97.64 58.07 97.64 58.07 96.28 58.77 96.28 58.77 97.64 58.99 97.64 58.99 96.28 59.69 96.28 59.69 97.64 59.91 97.64 59.91 96.28 60.61 96.28 60.61 97.64 60.83 97.64 60.83 96.28 61.53 96.28 61.53 97.64 61.75 97.64 61.75 96.28 62.45 96.28 62.45 97.64 63.13 97.64 63.13 96.28 63.83 96.28 63.83 97.64 64.05 97.64 64.05 96.28 64.75 96.28 64.75 97.64 64.97 97.64 64.97 96.28 65.67 96.28 65.67 97.64 65.89 97.64 65.89 96.28 66.59 96.28 66.59 97.64 66.81 97.64 66.81 96.28 67.51 96.28 67.51 97.64 67.73 97.64 67.73 96.28 68.43 96.28 68.43 97.64 70.49 97.64 70.49 96.28 71.19 96.28 71.19 97.64 76.93 97.64 76.93 96.28 77.63 96.28 77.63 97.64 77.85 97.64 77.85 96.28 78.55 96.28 78.55 97.64 78.77 97.64 78.77 96.28 79.47 96.28 79.47 97.64 79.69 97.64 79.69 96.28 80.39 96.28 80.39 97.64 80.61 97.64 80.61 96.28 81.31 96.28 81.31 97.64 ;
    LAYER met4 ;
      POLYGON 95.28 97.52 95.28 0.4 84.42 0.4 84.42 1 83.02 1 83.02 0.4 69.7 0.4 69.7 1 68.3 1 68.3 0.4 54.98 0.4 54.98 1 53.58 1 53.58 0.4 40.26 0.4 40.26 1 38.86 1 38.86 0.4 10.82 0.4 10.82 1 9.42 1 9.42 0.4 0.4 0.4 0.4 86.64 9.42 86.64 9.42 86.04 10.82 86.04 10.82 86.64 28 86.64 28 97.52 38.86 97.52 38.86 96.92 40.26 96.92 40.26 97.52 43.61 97.52 43.61 96.16 44.71 96.16 44.71 97.52 45.45 97.52 45.45 96.16 46.55 96.16 46.55 97.52 53.58 97.52 53.58 96.92 54.98 96.92 54.98 97.52 61.09 97.52 61.09 96.16 62.19 96.16 62.19 97.52 62.93 97.52 62.93 96.16 64.03 96.16 64.03 97.52 68.3 97.52 68.3 96.92 69.7 96.92 69.7 97.52 83.02 97.52 83.02 96.92 84.42 96.92 84.42 97.52 ;
    LAYER met5 ;
      POLYGON 94.08 96.32 94.08 77.32 90.88 77.32 90.88 70.92 94.08 70.92 94.08 56.92 90.88 56.92 90.88 50.52 94.08 50.52 94.08 36.52 90.88 36.52 90.88 30.12 94.08 30.12 94.08 16.12 90.88 16.12 90.88 9.72 94.08 9.72 94.08 1.6 1.6 1.6 1.6 9.72 4.8 9.72 4.8 16.12 1.6 16.12 1.6 30.12 4.8 30.12 4.8 36.52 1.6 36.52 1.6 50.52 4.8 50.52 4.8 56.92 1.6 56.92 1.6 70.92 4.8 70.92 4.8 77.32 1.6 77.32 1.6 85.44 29.2 85.44 29.2 96.32 ;
    LAYER met1 ;
      POLYGON 95.4 97.4 95.4 95.72 94.92 95.72 94.92 94.68 95.4 94.68 95.4 93 94.92 93 94.92 91.96 95.4 91.96 95.4 90.28 94.92 90.28 94.92 89.24 95.4 89.24 95.4 87.56 27.88 87.56 27.88 89.24 28.36 89.24 28.36 90.28 27.88 90.28 27.88 91.96 28.36 91.96 28.36 93 27.88 93 27.88 94.68 28.36 94.68 28.36 95.72 27.88 95.72 27.88 97.4 ;
      POLYGON 95.4 86.52 95.4 84.84 94.92 84.84 94.92 83.8 95.4 83.8 95.4 82.12 94.92 82.12 94.92 81.08 95.4 81.08 95.4 79.4 94.92 79.4 94.92 78.36 95.4 78.36 95.4 76.68 94.92 76.68 94.92 75.64 95.4 75.64 95.4 73.96 94.92 73.96 94.92 72.92 95.4 72.92 95.4 71.24 94.92 71.24 94.92 70.2 95.4 70.2 95.4 68.52 94.92 68.52 94.92 67.48 95.4 67.48 95.4 65.8 94.92 65.8 94.92 64.76 95.4 64.76 95.4 63.08 94.92 63.08 94.92 62.04 95.4 62.04 95.4 60.36 94.92 60.36 94.92 59.32 95.4 59.32 95.4 57.64 94.92 57.64 94.92 56.6 95.4 56.6 95.4 54.92 94.92 54.92 94.92 53.88 95.4 53.88 95.4 52.2 94.92 52.2 94.92 51.16 95.4 51.16 95.4 49.48 94.92 49.48 94.92 48.44 95.4 48.44 95.4 46.76 94.92 46.76 94.92 45.72 95.4 45.72 95.4 44.04 94.92 44.04 94.92 43 95.4 43 95.4 41.32 94.92 41.32 94.92 40.28 95.4 40.28 95.4 38.6 94.92 38.6 94.92 37.56 95.4 37.56 95.4 35.88 94.92 35.88 94.92 34.84 95.4 34.84 95.4 33.16 94.92 33.16 94.92 32.12 95.4 32.12 95.4 30.44 94.92 30.44 94.92 29.4 95.4 29.4 95.4 27.72 94.92 27.72 94.92 26.68 95.4 26.68 95.4 25 94.92 25 94.92 23.96 95.4 23.96 95.4 22.28 94.92 22.28 94.92 21.24 95.4 21.24 95.4 19.56 94.92 19.56 94.92 18.52 95.4 18.52 95.4 16.84 94.92 16.84 94.92 15.8 95.4 15.8 95.4 14.12 94.92 14.12 94.92 13.08 95.4 13.08 95.4 11.4 94.92 11.4 94.92 10.36 95.4 10.36 95.4 8.68 94.92 8.68 94.92 7.64 95.4 7.64 95.4 5.96 94.92 5.96 94.92 4.92 95.4 4.92 95.4 3.24 94.92 3.24 94.92 2.2 95.4 2.2 95.4 0.52 0.28 0.52 0.28 2.2 0.76 2.2 0.76 3.24 0.28 3.24 0.28 4.92 0.76 4.92 0.76 5.96 0.28 5.96 0.28 7.64 0.76 7.64 0.76 8.68 0.28 8.68 0.28 10.36 0.76 10.36 0.76 11.4 0.28 11.4 0.28 13.08 0.76 13.08 0.76 14.12 0.28 14.12 0.28 15.8 0.76 15.8 0.76 16.84 0.28 16.84 0.28 18.52 0.76 18.52 0.76 19.56 0.28 19.56 0.28 21.24 0.76 21.24 0.76 22.28 0.28 22.28 0.28 23.96 0.76 23.96 0.76 25 0.28 25 0.28 26.68 0.76 26.68 0.76 27.72 0.28 27.72 0.28 29.4 0.76 29.4 0.76 30.44 0.28 30.44 0.28 32.12 0.76 32.12 0.76 33.16 0.28 33.16 0.28 34.84 0.76 34.84 0.76 35.88 0.28 35.88 0.28 37.56 0.76 37.56 0.76 38.6 0.28 38.6 0.28 40.28 0.76 40.28 0.76 41.32 0.28 41.32 0.28 43 0.76 43 0.76 44.04 0.28 44.04 0.28 45.72 0.76 45.72 0.76 46.76 0.28 46.76 0.28 48.44 0.76 48.44 0.76 49.48 0.28 49.48 0.28 51.16 0.76 51.16 0.76 52.2 0.28 52.2 0.28 53.88 0.76 53.88 0.76 54.92 0.28 54.92 0.28 56.6 0.76 56.6 0.76 57.64 0.28 57.64 0.28 59.32 0.76 59.32 0.76 60.36 0.28 60.36 0.28 62.04 0.76 62.04 0.76 63.08 0.28 63.08 0.28 64.76 0.76 64.76 0.76 65.8 0.28 65.8 0.28 67.48 0.76 67.48 0.76 68.52 0.28 68.52 0.28 70.2 0.76 70.2 0.76 71.24 0.28 71.24 0.28 72.92 0.76 72.92 0.76 73.96 0.28 73.96 0.28 75.64 0.76 75.64 0.76 76.68 0.28 76.68 0.28 78.36 0.76 78.36 0.76 79.4 0.28 79.4 0.28 81.08 0.76 81.08 0.76 82.12 0.28 82.12 0.28 83.8 0.76 83.8 0.76 84.84 0.28 84.84 0.28 86.52 ;
    LAYER li1 ;
      POLYGON 95.51 97.75 95.51 0.17 0.17 0.17 0.17 86.87 27.77 86.87 27.77 97.75 ;
    LAYER mcon ;
      RECT 95.365 97.835 95.535 98.005 ;
      RECT 94.905 97.835 95.075 98.005 ;
      RECT 94.445 97.835 94.615 98.005 ;
      RECT 93.985 97.835 94.155 98.005 ;
      RECT 93.525 97.835 93.695 98.005 ;
      RECT 93.065 97.835 93.235 98.005 ;
      RECT 92.605 97.835 92.775 98.005 ;
      RECT 92.145 97.835 92.315 98.005 ;
      RECT 91.685 97.835 91.855 98.005 ;
      RECT 91.225 97.835 91.395 98.005 ;
      RECT 90.765 97.835 90.935 98.005 ;
      RECT 90.305 97.835 90.475 98.005 ;
      RECT 89.845 97.835 90.015 98.005 ;
      RECT 89.385 97.835 89.555 98.005 ;
      RECT 88.925 97.835 89.095 98.005 ;
      RECT 88.465 97.835 88.635 98.005 ;
      RECT 88.005 97.835 88.175 98.005 ;
      RECT 87.545 97.835 87.715 98.005 ;
      RECT 87.085 97.835 87.255 98.005 ;
      RECT 86.625 97.835 86.795 98.005 ;
      RECT 86.165 97.835 86.335 98.005 ;
      RECT 85.705 97.835 85.875 98.005 ;
      RECT 85.245 97.835 85.415 98.005 ;
      RECT 84.785 97.835 84.955 98.005 ;
      RECT 84.325 97.835 84.495 98.005 ;
      RECT 83.865 97.835 84.035 98.005 ;
      RECT 83.405 97.835 83.575 98.005 ;
      RECT 82.945 97.835 83.115 98.005 ;
      RECT 82.485 97.835 82.655 98.005 ;
      RECT 82.025 97.835 82.195 98.005 ;
      RECT 81.565 97.835 81.735 98.005 ;
      RECT 81.105 97.835 81.275 98.005 ;
      RECT 80.645 97.835 80.815 98.005 ;
      RECT 80.185 97.835 80.355 98.005 ;
      RECT 79.725 97.835 79.895 98.005 ;
      RECT 79.265 97.835 79.435 98.005 ;
      RECT 78.805 97.835 78.975 98.005 ;
      RECT 78.345 97.835 78.515 98.005 ;
      RECT 77.885 97.835 78.055 98.005 ;
      RECT 77.425 97.835 77.595 98.005 ;
      RECT 76.965 97.835 77.135 98.005 ;
      RECT 76.505 97.835 76.675 98.005 ;
      RECT 76.045 97.835 76.215 98.005 ;
      RECT 75.585 97.835 75.755 98.005 ;
      RECT 75.125 97.835 75.295 98.005 ;
      RECT 74.665 97.835 74.835 98.005 ;
      RECT 74.205 97.835 74.375 98.005 ;
      RECT 73.745 97.835 73.915 98.005 ;
      RECT 73.285 97.835 73.455 98.005 ;
      RECT 72.825 97.835 72.995 98.005 ;
      RECT 72.365 97.835 72.535 98.005 ;
      RECT 71.905 97.835 72.075 98.005 ;
      RECT 71.445 97.835 71.615 98.005 ;
      RECT 70.985 97.835 71.155 98.005 ;
      RECT 70.525 97.835 70.695 98.005 ;
      RECT 70.065 97.835 70.235 98.005 ;
      RECT 69.605 97.835 69.775 98.005 ;
      RECT 69.145 97.835 69.315 98.005 ;
      RECT 68.685 97.835 68.855 98.005 ;
      RECT 68.225 97.835 68.395 98.005 ;
      RECT 67.765 97.835 67.935 98.005 ;
      RECT 67.305 97.835 67.475 98.005 ;
      RECT 66.845 97.835 67.015 98.005 ;
      RECT 66.385 97.835 66.555 98.005 ;
      RECT 65.925 97.835 66.095 98.005 ;
      RECT 65.465 97.835 65.635 98.005 ;
      RECT 65.005 97.835 65.175 98.005 ;
      RECT 64.545 97.835 64.715 98.005 ;
      RECT 64.085 97.835 64.255 98.005 ;
      RECT 63.625 97.835 63.795 98.005 ;
      RECT 63.165 97.835 63.335 98.005 ;
      RECT 62.705 97.835 62.875 98.005 ;
      RECT 62.245 97.835 62.415 98.005 ;
      RECT 61.785 97.835 61.955 98.005 ;
      RECT 61.325 97.835 61.495 98.005 ;
      RECT 60.865 97.835 61.035 98.005 ;
      RECT 60.405 97.835 60.575 98.005 ;
      RECT 59.945 97.835 60.115 98.005 ;
      RECT 59.485 97.835 59.655 98.005 ;
      RECT 59.025 97.835 59.195 98.005 ;
      RECT 58.565 97.835 58.735 98.005 ;
      RECT 58.105 97.835 58.275 98.005 ;
      RECT 57.645 97.835 57.815 98.005 ;
      RECT 57.185 97.835 57.355 98.005 ;
      RECT 56.725 97.835 56.895 98.005 ;
      RECT 56.265 97.835 56.435 98.005 ;
      RECT 55.805 97.835 55.975 98.005 ;
      RECT 55.345 97.835 55.515 98.005 ;
      RECT 54.885 97.835 55.055 98.005 ;
      RECT 54.425 97.835 54.595 98.005 ;
      RECT 53.965 97.835 54.135 98.005 ;
      RECT 53.505 97.835 53.675 98.005 ;
      RECT 53.045 97.835 53.215 98.005 ;
      RECT 52.585 97.835 52.755 98.005 ;
      RECT 52.125 97.835 52.295 98.005 ;
      RECT 51.665 97.835 51.835 98.005 ;
      RECT 51.205 97.835 51.375 98.005 ;
      RECT 50.745 97.835 50.915 98.005 ;
      RECT 50.285 97.835 50.455 98.005 ;
      RECT 49.825 97.835 49.995 98.005 ;
      RECT 49.365 97.835 49.535 98.005 ;
      RECT 48.905 97.835 49.075 98.005 ;
      RECT 48.445 97.835 48.615 98.005 ;
      RECT 47.985 97.835 48.155 98.005 ;
      RECT 47.525 97.835 47.695 98.005 ;
      RECT 47.065 97.835 47.235 98.005 ;
      RECT 46.605 97.835 46.775 98.005 ;
      RECT 46.145 97.835 46.315 98.005 ;
      RECT 45.685 97.835 45.855 98.005 ;
      RECT 45.225 97.835 45.395 98.005 ;
      RECT 44.765 97.835 44.935 98.005 ;
      RECT 44.305 97.835 44.475 98.005 ;
      RECT 43.845 97.835 44.015 98.005 ;
      RECT 43.385 97.835 43.555 98.005 ;
      RECT 42.925 97.835 43.095 98.005 ;
      RECT 42.465 97.835 42.635 98.005 ;
      RECT 42.005 97.835 42.175 98.005 ;
      RECT 41.545 97.835 41.715 98.005 ;
      RECT 41.085 97.835 41.255 98.005 ;
      RECT 40.625 97.835 40.795 98.005 ;
      RECT 40.165 97.835 40.335 98.005 ;
      RECT 39.705 97.835 39.875 98.005 ;
      RECT 39.245 97.835 39.415 98.005 ;
      RECT 38.785 97.835 38.955 98.005 ;
      RECT 38.325 97.835 38.495 98.005 ;
      RECT 37.865 97.835 38.035 98.005 ;
      RECT 37.405 97.835 37.575 98.005 ;
      RECT 36.945 97.835 37.115 98.005 ;
      RECT 36.485 97.835 36.655 98.005 ;
      RECT 36.025 97.835 36.195 98.005 ;
      RECT 35.565 97.835 35.735 98.005 ;
      RECT 35.105 97.835 35.275 98.005 ;
      RECT 34.645 97.835 34.815 98.005 ;
      RECT 34.185 97.835 34.355 98.005 ;
      RECT 33.725 97.835 33.895 98.005 ;
      RECT 33.265 97.835 33.435 98.005 ;
      RECT 32.805 97.835 32.975 98.005 ;
      RECT 32.345 97.835 32.515 98.005 ;
      RECT 31.885 97.835 32.055 98.005 ;
      RECT 31.425 97.835 31.595 98.005 ;
      RECT 30.965 97.835 31.135 98.005 ;
      RECT 30.505 97.835 30.675 98.005 ;
      RECT 30.045 97.835 30.215 98.005 ;
      RECT 29.585 97.835 29.755 98.005 ;
      RECT 29.125 97.835 29.295 98.005 ;
      RECT 28.665 97.835 28.835 98.005 ;
      RECT 28.205 97.835 28.375 98.005 ;
      RECT 27.745 97.835 27.915 98.005 ;
      RECT 95.365 95.115 95.535 95.285 ;
      RECT 94.905 95.115 95.075 95.285 ;
      RECT 28.205 95.115 28.375 95.285 ;
      RECT 27.745 95.115 27.915 95.285 ;
      RECT 95.365 92.395 95.535 92.565 ;
      RECT 94.905 92.395 95.075 92.565 ;
      RECT 28.205 92.395 28.375 92.565 ;
      RECT 27.745 92.395 27.915 92.565 ;
      RECT 95.365 89.675 95.535 89.845 ;
      RECT 94.905 89.675 95.075 89.845 ;
      RECT 28.205 89.675 28.375 89.845 ;
      RECT 27.745 89.675 27.915 89.845 ;
      RECT 95.365 86.955 95.535 87.125 ;
      RECT 94.905 86.955 95.075 87.125 ;
      RECT 94.445 86.955 94.615 87.125 ;
      RECT 93.985 86.955 94.155 87.125 ;
      RECT 93.525 86.955 93.695 87.125 ;
      RECT 93.065 86.955 93.235 87.125 ;
      RECT 92.605 86.955 92.775 87.125 ;
      RECT 92.145 86.955 92.315 87.125 ;
      RECT 91.685 86.955 91.855 87.125 ;
      RECT 91.225 86.955 91.395 87.125 ;
      RECT 90.765 86.955 90.935 87.125 ;
      RECT 90.305 86.955 90.475 87.125 ;
      RECT 89.845 86.955 90.015 87.125 ;
      RECT 89.385 86.955 89.555 87.125 ;
      RECT 88.925 86.955 89.095 87.125 ;
      RECT 88.465 86.955 88.635 87.125 ;
      RECT 88.005 86.955 88.175 87.125 ;
      RECT 87.545 86.955 87.715 87.125 ;
      RECT 87.085 86.955 87.255 87.125 ;
      RECT 86.625 86.955 86.795 87.125 ;
      RECT 86.165 86.955 86.335 87.125 ;
      RECT 85.705 86.955 85.875 87.125 ;
      RECT 85.245 86.955 85.415 87.125 ;
      RECT 84.785 86.955 84.955 87.125 ;
      RECT 84.325 86.955 84.495 87.125 ;
      RECT 83.865 86.955 84.035 87.125 ;
      RECT 83.405 86.955 83.575 87.125 ;
      RECT 82.945 86.955 83.115 87.125 ;
      RECT 82.485 86.955 82.655 87.125 ;
      RECT 82.025 86.955 82.195 87.125 ;
      RECT 81.565 86.955 81.735 87.125 ;
      RECT 81.105 86.955 81.275 87.125 ;
      RECT 80.645 86.955 80.815 87.125 ;
      RECT 80.185 86.955 80.355 87.125 ;
      RECT 79.725 86.955 79.895 87.125 ;
      RECT 79.265 86.955 79.435 87.125 ;
      RECT 78.805 86.955 78.975 87.125 ;
      RECT 78.345 86.955 78.515 87.125 ;
      RECT 77.885 86.955 78.055 87.125 ;
      RECT 77.425 86.955 77.595 87.125 ;
      RECT 76.965 86.955 77.135 87.125 ;
      RECT 76.505 86.955 76.675 87.125 ;
      RECT 76.045 86.955 76.215 87.125 ;
      RECT 75.585 86.955 75.755 87.125 ;
      RECT 75.125 86.955 75.295 87.125 ;
      RECT 74.665 86.955 74.835 87.125 ;
      RECT 74.205 86.955 74.375 87.125 ;
      RECT 73.745 86.955 73.915 87.125 ;
      RECT 73.285 86.955 73.455 87.125 ;
      RECT 72.825 86.955 72.995 87.125 ;
      RECT 72.365 86.955 72.535 87.125 ;
      RECT 71.905 86.955 72.075 87.125 ;
      RECT 71.445 86.955 71.615 87.125 ;
      RECT 70.985 86.955 71.155 87.125 ;
      RECT 70.525 86.955 70.695 87.125 ;
      RECT 70.065 86.955 70.235 87.125 ;
      RECT 69.605 86.955 69.775 87.125 ;
      RECT 69.145 86.955 69.315 87.125 ;
      RECT 68.685 86.955 68.855 87.125 ;
      RECT 68.225 86.955 68.395 87.125 ;
      RECT 67.765 86.955 67.935 87.125 ;
      RECT 67.305 86.955 67.475 87.125 ;
      RECT 66.845 86.955 67.015 87.125 ;
      RECT 66.385 86.955 66.555 87.125 ;
      RECT 65.925 86.955 66.095 87.125 ;
      RECT 65.465 86.955 65.635 87.125 ;
      RECT 65.005 86.955 65.175 87.125 ;
      RECT 64.545 86.955 64.715 87.125 ;
      RECT 64.085 86.955 64.255 87.125 ;
      RECT 63.625 86.955 63.795 87.125 ;
      RECT 63.165 86.955 63.335 87.125 ;
      RECT 62.705 86.955 62.875 87.125 ;
      RECT 62.245 86.955 62.415 87.125 ;
      RECT 61.785 86.955 61.955 87.125 ;
      RECT 61.325 86.955 61.495 87.125 ;
      RECT 60.865 86.955 61.035 87.125 ;
      RECT 60.405 86.955 60.575 87.125 ;
      RECT 59.945 86.955 60.115 87.125 ;
      RECT 59.485 86.955 59.655 87.125 ;
      RECT 59.025 86.955 59.195 87.125 ;
      RECT 58.565 86.955 58.735 87.125 ;
      RECT 58.105 86.955 58.275 87.125 ;
      RECT 57.645 86.955 57.815 87.125 ;
      RECT 57.185 86.955 57.355 87.125 ;
      RECT 56.725 86.955 56.895 87.125 ;
      RECT 56.265 86.955 56.435 87.125 ;
      RECT 55.805 86.955 55.975 87.125 ;
      RECT 55.345 86.955 55.515 87.125 ;
      RECT 54.885 86.955 55.055 87.125 ;
      RECT 54.425 86.955 54.595 87.125 ;
      RECT 53.965 86.955 54.135 87.125 ;
      RECT 53.505 86.955 53.675 87.125 ;
      RECT 53.045 86.955 53.215 87.125 ;
      RECT 52.585 86.955 52.755 87.125 ;
      RECT 52.125 86.955 52.295 87.125 ;
      RECT 51.665 86.955 51.835 87.125 ;
      RECT 51.205 86.955 51.375 87.125 ;
      RECT 50.745 86.955 50.915 87.125 ;
      RECT 50.285 86.955 50.455 87.125 ;
      RECT 49.825 86.955 49.995 87.125 ;
      RECT 49.365 86.955 49.535 87.125 ;
      RECT 48.905 86.955 49.075 87.125 ;
      RECT 48.445 86.955 48.615 87.125 ;
      RECT 47.985 86.955 48.155 87.125 ;
      RECT 47.525 86.955 47.695 87.125 ;
      RECT 47.065 86.955 47.235 87.125 ;
      RECT 46.605 86.955 46.775 87.125 ;
      RECT 46.145 86.955 46.315 87.125 ;
      RECT 45.685 86.955 45.855 87.125 ;
      RECT 45.225 86.955 45.395 87.125 ;
      RECT 44.765 86.955 44.935 87.125 ;
      RECT 44.305 86.955 44.475 87.125 ;
      RECT 43.845 86.955 44.015 87.125 ;
      RECT 43.385 86.955 43.555 87.125 ;
      RECT 42.925 86.955 43.095 87.125 ;
      RECT 42.465 86.955 42.635 87.125 ;
      RECT 42.005 86.955 42.175 87.125 ;
      RECT 41.545 86.955 41.715 87.125 ;
      RECT 41.085 86.955 41.255 87.125 ;
      RECT 40.625 86.955 40.795 87.125 ;
      RECT 40.165 86.955 40.335 87.125 ;
      RECT 39.705 86.955 39.875 87.125 ;
      RECT 39.245 86.955 39.415 87.125 ;
      RECT 38.785 86.955 38.955 87.125 ;
      RECT 38.325 86.955 38.495 87.125 ;
      RECT 37.865 86.955 38.035 87.125 ;
      RECT 37.405 86.955 37.575 87.125 ;
      RECT 36.945 86.955 37.115 87.125 ;
      RECT 36.485 86.955 36.655 87.125 ;
      RECT 36.025 86.955 36.195 87.125 ;
      RECT 35.565 86.955 35.735 87.125 ;
      RECT 35.105 86.955 35.275 87.125 ;
      RECT 34.645 86.955 34.815 87.125 ;
      RECT 34.185 86.955 34.355 87.125 ;
      RECT 33.725 86.955 33.895 87.125 ;
      RECT 33.265 86.955 33.435 87.125 ;
      RECT 32.805 86.955 32.975 87.125 ;
      RECT 32.345 86.955 32.515 87.125 ;
      RECT 31.885 86.955 32.055 87.125 ;
      RECT 31.425 86.955 31.595 87.125 ;
      RECT 30.965 86.955 31.135 87.125 ;
      RECT 30.505 86.955 30.675 87.125 ;
      RECT 30.045 86.955 30.215 87.125 ;
      RECT 29.585 86.955 29.755 87.125 ;
      RECT 29.125 86.955 29.295 87.125 ;
      RECT 28.665 86.955 28.835 87.125 ;
      RECT 28.205 86.955 28.375 87.125 ;
      RECT 27.745 86.955 27.915 87.125 ;
      RECT 27.285 86.955 27.455 87.125 ;
      RECT 26.825 86.955 26.995 87.125 ;
      RECT 26.365 86.955 26.535 87.125 ;
      RECT 25.905 86.955 26.075 87.125 ;
      RECT 25.445 86.955 25.615 87.125 ;
      RECT 24.985 86.955 25.155 87.125 ;
      RECT 24.525 86.955 24.695 87.125 ;
      RECT 24.065 86.955 24.235 87.125 ;
      RECT 23.605 86.955 23.775 87.125 ;
      RECT 23.145 86.955 23.315 87.125 ;
      RECT 22.685 86.955 22.855 87.125 ;
      RECT 22.225 86.955 22.395 87.125 ;
      RECT 21.765 86.955 21.935 87.125 ;
      RECT 21.305 86.955 21.475 87.125 ;
      RECT 20.845 86.955 21.015 87.125 ;
      RECT 20.385 86.955 20.555 87.125 ;
      RECT 19.925 86.955 20.095 87.125 ;
      RECT 19.465 86.955 19.635 87.125 ;
      RECT 19.005 86.955 19.175 87.125 ;
      RECT 18.545 86.955 18.715 87.125 ;
      RECT 18.085 86.955 18.255 87.125 ;
      RECT 17.625 86.955 17.795 87.125 ;
      RECT 17.165 86.955 17.335 87.125 ;
      RECT 16.705 86.955 16.875 87.125 ;
      RECT 16.245 86.955 16.415 87.125 ;
      RECT 15.785 86.955 15.955 87.125 ;
      RECT 15.325 86.955 15.495 87.125 ;
      RECT 14.865 86.955 15.035 87.125 ;
      RECT 14.405 86.955 14.575 87.125 ;
      RECT 13.945 86.955 14.115 87.125 ;
      RECT 13.485 86.955 13.655 87.125 ;
      RECT 13.025 86.955 13.195 87.125 ;
      RECT 12.565 86.955 12.735 87.125 ;
      RECT 12.105 86.955 12.275 87.125 ;
      RECT 11.645 86.955 11.815 87.125 ;
      RECT 11.185 86.955 11.355 87.125 ;
      RECT 10.725 86.955 10.895 87.125 ;
      RECT 10.265 86.955 10.435 87.125 ;
      RECT 9.805 86.955 9.975 87.125 ;
      RECT 9.345 86.955 9.515 87.125 ;
      RECT 8.885 86.955 9.055 87.125 ;
      RECT 8.425 86.955 8.595 87.125 ;
      RECT 7.965 86.955 8.135 87.125 ;
      RECT 7.505 86.955 7.675 87.125 ;
      RECT 7.045 86.955 7.215 87.125 ;
      RECT 6.585 86.955 6.755 87.125 ;
      RECT 6.125 86.955 6.295 87.125 ;
      RECT 5.665 86.955 5.835 87.125 ;
      RECT 5.205 86.955 5.375 87.125 ;
      RECT 4.745 86.955 4.915 87.125 ;
      RECT 4.285 86.955 4.455 87.125 ;
      RECT 3.825 86.955 3.995 87.125 ;
      RECT 3.365 86.955 3.535 87.125 ;
      RECT 2.905 86.955 3.075 87.125 ;
      RECT 2.445 86.955 2.615 87.125 ;
      RECT 1.985 86.955 2.155 87.125 ;
      RECT 1.525 86.955 1.695 87.125 ;
      RECT 1.065 86.955 1.235 87.125 ;
      RECT 0.605 86.955 0.775 87.125 ;
      RECT 0.145 86.955 0.315 87.125 ;
      RECT 95.365 84.235 95.535 84.405 ;
      RECT 94.905 84.235 95.075 84.405 ;
      RECT 0.605 84.235 0.775 84.405 ;
      RECT 0.145 84.235 0.315 84.405 ;
      RECT 95.365 81.515 95.535 81.685 ;
      RECT 94.905 81.515 95.075 81.685 ;
      RECT 0.605 81.515 0.775 81.685 ;
      RECT 0.145 81.515 0.315 81.685 ;
      RECT 95.365 78.795 95.535 78.965 ;
      RECT 94.905 78.795 95.075 78.965 ;
      RECT 0.605 78.795 0.775 78.965 ;
      RECT 0.145 78.795 0.315 78.965 ;
      RECT 95.365 76.075 95.535 76.245 ;
      RECT 94.905 76.075 95.075 76.245 ;
      RECT 0.605 76.075 0.775 76.245 ;
      RECT 0.145 76.075 0.315 76.245 ;
      RECT 95.365 73.355 95.535 73.525 ;
      RECT 94.905 73.355 95.075 73.525 ;
      RECT 0.605 73.355 0.775 73.525 ;
      RECT 0.145 73.355 0.315 73.525 ;
      RECT 95.365 70.635 95.535 70.805 ;
      RECT 94.905 70.635 95.075 70.805 ;
      RECT 0.605 70.635 0.775 70.805 ;
      RECT 0.145 70.635 0.315 70.805 ;
      RECT 95.365 67.915 95.535 68.085 ;
      RECT 94.905 67.915 95.075 68.085 ;
      RECT 0.605 67.915 0.775 68.085 ;
      RECT 0.145 67.915 0.315 68.085 ;
      RECT 95.365 65.195 95.535 65.365 ;
      RECT 94.905 65.195 95.075 65.365 ;
      RECT 0.605 65.195 0.775 65.365 ;
      RECT 0.145 65.195 0.315 65.365 ;
      RECT 95.365 62.475 95.535 62.645 ;
      RECT 94.905 62.475 95.075 62.645 ;
      RECT 0.605 62.475 0.775 62.645 ;
      RECT 0.145 62.475 0.315 62.645 ;
      RECT 95.365 59.755 95.535 59.925 ;
      RECT 94.905 59.755 95.075 59.925 ;
      RECT 0.605 59.755 0.775 59.925 ;
      RECT 0.145 59.755 0.315 59.925 ;
      RECT 95.365 57.035 95.535 57.205 ;
      RECT 94.905 57.035 95.075 57.205 ;
      RECT 0.605 57.035 0.775 57.205 ;
      RECT 0.145 57.035 0.315 57.205 ;
      RECT 95.365 54.315 95.535 54.485 ;
      RECT 94.905 54.315 95.075 54.485 ;
      RECT 0.605 54.315 0.775 54.485 ;
      RECT 0.145 54.315 0.315 54.485 ;
      RECT 95.365 51.595 95.535 51.765 ;
      RECT 94.905 51.595 95.075 51.765 ;
      RECT 0.605 51.595 0.775 51.765 ;
      RECT 0.145 51.595 0.315 51.765 ;
      RECT 95.365 48.875 95.535 49.045 ;
      RECT 94.905 48.875 95.075 49.045 ;
      RECT 0.605 48.875 0.775 49.045 ;
      RECT 0.145 48.875 0.315 49.045 ;
      RECT 95.365 46.155 95.535 46.325 ;
      RECT 94.905 46.155 95.075 46.325 ;
      RECT 0.605 46.155 0.775 46.325 ;
      RECT 0.145 46.155 0.315 46.325 ;
      RECT 95.365 43.435 95.535 43.605 ;
      RECT 94.905 43.435 95.075 43.605 ;
      RECT 0.605 43.435 0.775 43.605 ;
      RECT 0.145 43.435 0.315 43.605 ;
      RECT 95.365 40.715 95.535 40.885 ;
      RECT 94.905 40.715 95.075 40.885 ;
      RECT 0.605 40.715 0.775 40.885 ;
      RECT 0.145 40.715 0.315 40.885 ;
      RECT 95.365 37.995 95.535 38.165 ;
      RECT 94.905 37.995 95.075 38.165 ;
      RECT 0.605 37.995 0.775 38.165 ;
      RECT 0.145 37.995 0.315 38.165 ;
      RECT 95.365 35.275 95.535 35.445 ;
      RECT 94.905 35.275 95.075 35.445 ;
      RECT 0.605 35.275 0.775 35.445 ;
      RECT 0.145 35.275 0.315 35.445 ;
      RECT 95.365 32.555 95.535 32.725 ;
      RECT 94.905 32.555 95.075 32.725 ;
      RECT 0.605 32.555 0.775 32.725 ;
      RECT 0.145 32.555 0.315 32.725 ;
      RECT 95.365 29.835 95.535 30.005 ;
      RECT 94.905 29.835 95.075 30.005 ;
      RECT 0.605 29.835 0.775 30.005 ;
      RECT 0.145 29.835 0.315 30.005 ;
      RECT 95.365 27.115 95.535 27.285 ;
      RECT 94.905 27.115 95.075 27.285 ;
      RECT 0.605 27.115 0.775 27.285 ;
      RECT 0.145 27.115 0.315 27.285 ;
      RECT 95.365 24.395 95.535 24.565 ;
      RECT 94.905 24.395 95.075 24.565 ;
      RECT 0.605 24.395 0.775 24.565 ;
      RECT 0.145 24.395 0.315 24.565 ;
      RECT 95.365 21.675 95.535 21.845 ;
      RECT 94.905 21.675 95.075 21.845 ;
      RECT 0.605 21.675 0.775 21.845 ;
      RECT 0.145 21.675 0.315 21.845 ;
      RECT 95.365 18.955 95.535 19.125 ;
      RECT 94.905 18.955 95.075 19.125 ;
      RECT 0.605 18.955 0.775 19.125 ;
      RECT 0.145 18.955 0.315 19.125 ;
      RECT 95.365 16.235 95.535 16.405 ;
      RECT 94.905 16.235 95.075 16.405 ;
      RECT 0.605 16.235 0.775 16.405 ;
      RECT 0.145 16.235 0.315 16.405 ;
      RECT 95.365 13.515 95.535 13.685 ;
      RECT 94.905 13.515 95.075 13.685 ;
      RECT 0.605 13.515 0.775 13.685 ;
      RECT 0.145 13.515 0.315 13.685 ;
      RECT 95.365 10.795 95.535 10.965 ;
      RECT 94.905 10.795 95.075 10.965 ;
      RECT 0.605 10.795 0.775 10.965 ;
      RECT 0.145 10.795 0.315 10.965 ;
      RECT 95.365 8.075 95.535 8.245 ;
      RECT 94.905 8.075 95.075 8.245 ;
      RECT 0.605 8.075 0.775 8.245 ;
      RECT 0.145 8.075 0.315 8.245 ;
      RECT 95.365 5.355 95.535 5.525 ;
      RECT 94.905 5.355 95.075 5.525 ;
      RECT 0.605 5.355 0.775 5.525 ;
      RECT 0.145 5.355 0.315 5.525 ;
      RECT 95.365 2.635 95.535 2.805 ;
      RECT 94.905 2.635 95.075 2.805 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 95.365 -0.085 95.535 0.085 ;
      RECT 94.905 -0.085 95.075 0.085 ;
      RECT 94.445 -0.085 94.615 0.085 ;
      RECT 93.985 -0.085 94.155 0.085 ;
      RECT 93.525 -0.085 93.695 0.085 ;
      RECT 93.065 -0.085 93.235 0.085 ;
      RECT 92.605 -0.085 92.775 0.085 ;
      RECT 92.145 -0.085 92.315 0.085 ;
      RECT 91.685 -0.085 91.855 0.085 ;
      RECT 91.225 -0.085 91.395 0.085 ;
      RECT 90.765 -0.085 90.935 0.085 ;
      RECT 90.305 -0.085 90.475 0.085 ;
      RECT 89.845 -0.085 90.015 0.085 ;
      RECT 89.385 -0.085 89.555 0.085 ;
      RECT 88.925 -0.085 89.095 0.085 ;
      RECT 88.465 -0.085 88.635 0.085 ;
      RECT 88.005 -0.085 88.175 0.085 ;
      RECT 87.545 -0.085 87.715 0.085 ;
      RECT 87.085 -0.085 87.255 0.085 ;
      RECT 86.625 -0.085 86.795 0.085 ;
      RECT 86.165 -0.085 86.335 0.085 ;
      RECT 85.705 -0.085 85.875 0.085 ;
      RECT 85.245 -0.085 85.415 0.085 ;
      RECT 84.785 -0.085 84.955 0.085 ;
      RECT 84.325 -0.085 84.495 0.085 ;
      RECT 83.865 -0.085 84.035 0.085 ;
      RECT 83.405 -0.085 83.575 0.085 ;
      RECT 82.945 -0.085 83.115 0.085 ;
      RECT 82.485 -0.085 82.655 0.085 ;
      RECT 82.025 -0.085 82.195 0.085 ;
      RECT 81.565 -0.085 81.735 0.085 ;
      RECT 81.105 -0.085 81.275 0.085 ;
      RECT 80.645 -0.085 80.815 0.085 ;
      RECT 80.185 -0.085 80.355 0.085 ;
      RECT 79.725 -0.085 79.895 0.085 ;
      RECT 79.265 -0.085 79.435 0.085 ;
      RECT 78.805 -0.085 78.975 0.085 ;
      RECT 78.345 -0.085 78.515 0.085 ;
      RECT 77.885 -0.085 78.055 0.085 ;
      RECT 77.425 -0.085 77.595 0.085 ;
      RECT 76.965 -0.085 77.135 0.085 ;
      RECT 76.505 -0.085 76.675 0.085 ;
      RECT 76.045 -0.085 76.215 0.085 ;
      RECT 75.585 -0.085 75.755 0.085 ;
      RECT 75.125 -0.085 75.295 0.085 ;
      RECT 74.665 -0.085 74.835 0.085 ;
      RECT 74.205 -0.085 74.375 0.085 ;
      RECT 73.745 -0.085 73.915 0.085 ;
      RECT 73.285 -0.085 73.455 0.085 ;
      RECT 72.825 -0.085 72.995 0.085 ;
      RECT 72.365 -0.085 72.535 0.085 ;
      RECT 71.905 -0.085 72.075 0.085 ;
      RECT 71.445 -0.085 71.615 0.085 ;
      RECT 70.985 -0.085 71.155 0.085 ;
      RECT 70.525 -0.085 70.695 0.085 ;
      RECT 70.065 -0.085 70.235 0.085 ;
      RECT 69.605 -0.085 69.775 0.085 ;
      RECT 69.145 -0.085 69.315 0.085 ;
      RECT 68.685 -0.085 68.855 0.085 ;
      RECT 68.225 -0.085 68.395 0.085 ;
      RECT 67.765 -0.085 67.935 0.085 ;
      RECT 67.305 -0.085 67.475 0.085 ;
      RECT 66.845 -0.085 67.015 0.085 ;
      RECT 66.385 -0.085 66.555 0.085 ;
      RECT 65.925 -0.085 66.095 0.085 ;
      RECT 65.465 -0.085 65.635 0.085 ;
      RECT 65.005 -0.085 65.175 0.085 ;
      RECT 64.545 -0.085 64.715 0.085 ;
      RECT 64.085 -0.085 64.255 0.085 ;
      RECT 63.625 -0.085 63.795 0.085 ;
      RECT 63.165 -0.085 63.335 0.085 ;
      RECT 62.705 -0.085 62.875 0.085 ;
      RECT 62.245 -0.085 62.415 0.085 ;
      RECT 61.785 -0.085 61.955 0.085 ;
      RECT 61.325 -0.085 61.495 0.085 ;
      RECT 60.865 -0.085 61.035 0.085 ;
      RECT 60.405 -0.085 60.575 0.085 ;
      RECT 59.945 -0.085 60.115 0.085 ;
      RECT 59.485 -0.085 59.655 0.085 ;
      RECT 59.025 -0.085 59.195 0.085 ;
      RECT 58.565 -0.085 58.735 0.085 ;
      RECT 58.105 -0.085 58.275 0.085 ;
      RECT 57.645 -0.085 57.815 0.085 ;
      RECT 57.185 -0.085 57.355 0.085 ;
      RECT 56.725 -0.085 56.895 0.085 ;
      RECT 56.265 -0.085 56.435 0.085 ;
      RECT 55.805 -0.085 55.975 0.085 ;
      RECT 55.345 -0.085 55.515 0.085 ;
      RECT 54.885 -0.085 55.055 0.085 ;
      RECT 54.425 -0.085 54.595 0.085 ;
      RECT 53.965 -0.085 54.135 0.085 ;
      RECT 53.505 -0.085 53.675 0.085 ;
      RECT 53.045 -0.085 53.215 0.085 ;
      RECT 52.585 -0.085 52.755 0.085 ;
      RECT 52.125 -0.085 52.295 0.085 ;
      RECT 51.665 -0.085 51.835 0.085 ;
      RECT 51.205 -0.085 51.375 0.085 ;
      RECT 50.745 -0.085 50.915 0.085 ;
      RECT 50.285 -0.085 50.455 0.085 ;
      RECT 49.825 -0.085 49.995 0.085 ;
      RECT 49.365 -0.085 49.535 0.085 ;
      RECT 48.905 -0.085 49.075 0.085 ;
      RECT 48.445 -0.085 48.615 0.085 ;
      RECT 47.985 -0.085 48.155 0.085 ;
      RECT 47.525 -0.085 47.695 0.085 ;
      RECT 47.065 -0.085 47.235 0.085 ;
      RECT 46.605 -0.085 46.775 0.085 ;
      RECT 46.145 -0.085 46.315 0.085 ;
      RECT 45.685 -0.085 45.855 0.085 ;
      RECT 45.225 -0.085 45.395 0.085 ;
      RECT 44.765 -0.085 44.935 0.085 ;
      RECT 44.305 -0.085 44.475 0.085 ;
      RECT 43.845 -0.085 44.015 0.085 ;
      RECT 43.385 -0.085 43.555 0.085 ;
      RECT 42.925 -0.085 43.095 0.085 ;
      RECT 42.465 -0.085 42.635 0.085 ;
      RECT 42.005 -0.085 42.175 0.085 ;
      RECT 41.545 -0.085 41.715 0.085 ;
      RECT 41.085 -0.085 41.255 0.085 ;
      RECT 40.625 -0.085 40.795 0.085 ;
      RECT 40.165 -0.085 40.335 0.085 ;
      RECT 39.705 -0.085 39.875 0.085 ;
      RECT 39.245 -0.085 39.415 0.085 ;
      RECT 38.785 -0.085 38.955 0.085 ;
      RECT 38.325 -0.085 38.495 0.085 ;
      RECT 37.865 -0.085 38.035 0.085 ;
      RECT 37.405 -0.085 37.575 0.085 ;
      RECT 36.945 -0.085 37.115 0.085 ;
      RECT 36.485 -0.085 36.655 0.085 ;
      RECT 36.025 -0.085 36.195 0.085 ;
      RECT 35.565 -0.085 35.735 0.085 ;
      RECT 35.105 -0.085 35.275 0.085 ;
      RECT 34.645 -0.085 34.815 0.085 ;
      RECT 34.185 -0.085 34.355 0.085 ;
      RECT 33.725 -0.085 33.895 0.085 ;
      RECT 33.265 -0.085 33.435 0.085 ;
      RECT 32.805 -0.085 32.975 0.085 ;
      RECT 32.345 -0.085 32.515 0.085 ;
      RECT 31.885 -0.085 32.055 0.085 ;
      RECT 31.425 -0.085 31.595 0.085 ;
      RECT 30.965 -0.085 31.135 0.085 ;
      RECT 30.505 -0.085 30.675 0.085 ;
      RECT 30.045 -0.085 30.215 0.085 ;
      RECT 29.585 -0.085 29.755 0.085 ;
      RECT 29.125 -0.085 29.295 0.085 ;
      RECT 28.665 -0.085 28.835 0.085 ;
      RECT 28.205 -0.085 28.375 0.085 ;
      RECT 27.745 -0.085 27.915 0.085 ;
      RECT 27.285 -0.085 27.455 0.085 ;
      RECT 26.825 -0.085 26.995 0.085 ;
      RECT 26.365 -0.085 26.535 0.085 ;
      RECT 25.905 -0.085 26.075 0.085 ;
      RECT 25.445 -0.085 25.615 0.085 ;
      RECT 24.985 -0.085 25.155 0.085 ;
      RECT 24.525 -0.085 24.695 0.085 ;
      RECT 24.065 -0.085 24.235 0.085 ;
      RECT 23.605 -0.085 23.775 0.085 ;
      RECT 23.145 -0.085 23.315 0.085 ;
      RECT 22.685 -0.085 22.855 0.085 ;
      RECT 22.225 -0.085 22.395 0.085 ;
      RECT 21.765 -0.085 21.935 0.085 ;
      RECT 21.305 -0.085 21.475 0.085 ;
      RECT 20.845 -0.085 21.015 0.085 ;
      RECT 20.385 -0.085 20.555 0.085 ;
      RECT 19.925 -0.085 20.095 0.085 ;
      RECT 19.465 -0.085 19.635 0.085 ;
      RECT 19.005 -0.085 19.175 0.085 ;
      RECT 18.545 -0.085 18.715 0.085 ;
      RECT 18.085 -0.085 18.255 0.085 ;
      RECT 17.625 -0.085 17.795 0.085 ;
      RECT 17.165 -0.085 17.335 0.085 ;
      RECT 16.705 -0.085 16.875 0.085 ;
      RECT 16.245 -0.085 16.415 0.085 ;
      RECT 15.785 -0.085 15.955 0.085 ;
      RECT 15.325 -0.085 15.495 0.085 ;
      RECT 14.865 -0.085 15.035 0.085 ;
      RECT 14.405 -0.085 14.575 0.085 ;
      RECT 13.945 -0.085 14.115 0.085 ;
      RECT 13.485 -0.085 13.655 0.085 ;
      RECT 13.025 -0.085 13.195 0.085 ;
      RECT 12.565 -0.085 12.735 0.085 ;
      RECT 12.105 -0.085 12.275 0.085 ;
      RECT 11.645 -0.085 11.815 0.085 ;
      RECT 11.185 -0.085 11.355 0.085 ;
      RECT 10.725 -0.085 10.895 0.085 ;
      RECT 10.265 -0.085 10.435 0.085 ;
      RECT 9.805 -0.085 9.975 0.085 ;
      RECT 9.345 -0.085 9.515 0.085 ;
      RECT 8.885 -0.085 9.055 0.085 ;
      RECT 8.425 -0.085 8.595 0.085 ;
      RECT 7.965 -0.085 8.135 0.085 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.145 -0.085 0.315 0.085 ;
    LAYER via ;
      RECT 83.645 97.845 83.795 97.995 ;
      RECT 54.205 97.845 54.355 97.995 ;
      RECT 67.085 96.145 67.235 96.295 ;
      RECT 46.385 96.145 46.535 96.295 ;
      RECT 38.105 96.145 38.255 96.295 ;
      RECT 83.645 86.965 83.795 87.115 ;
      RECT 54.205 86.965 54.355 87.115 ;
      RECT 10.045 86.965 10.195 87.115 ;
      RECT 8.205 85.265 8.355 85.415 ;
      RECT 83.645 -0.075 83.795 0.075 ;
      RECT 54.205 -0.075 54.355 0.075 ;
      RECT 10.045 -0.075 10.195 0.075 ;
    LAYER via2 ;
      RECT 83.62 97.82 83.82 98.02 ;
      RECT 54.18 97.82 54.38 98.02 ;
      RECT 10.02 86.94 10.22 87.14 ;
      RECT 1.28 76.74 1.48 76.94 ;
      RECT 1.74 74.02 1.94 74.22 ;
      RECT 1.74 61.1 1.94 61.3 ;
      RECT 1.28 57.02 1.48 57.22 ;
      RECT 1.28 52.94 1.48 53.14 ;
      RECT 1.28 33.9 1.48 34.1 ;
      RECT 1.28 26.42 1.48 26.62 ;
      RECT 1.74 20.3 1.94 20.5 ;
      RECT 1.28 13.5 1.48 13.7 ;
      RECT 83.62 -0.1 83.82 0.1 ;
      RECT 54.18 -0.1 54.38 0.1 ;
      RECT 10.02 -0.1 10.22 0.1 ;
    LAYER via3 ;
      RECT 83.62 97.82 83.82 98.02 ;
      RECT 54.18 97.82 54.38 98.02 ;
      RECT 10.02 86.94 10.22 87.14 ;
      RECT 83.62 -0.1 83.82 0.1 ;
      RECT 54.18 -0.1 54.38 0.1 ;
      RECT 10.02 -0.1 10.22 0.1 ;
    LAYER OVERLAP ;
      POLYGON 0 0 0 87.04 27.6 87.04 27.6 97.92 95.68 97.92 95.68 0 ;
  END
END sb_2__0_

END LIBRARY
