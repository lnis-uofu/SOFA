VERSION 5.7 ;
BUSBITCHARS "[]" ;

UNITS
  DATABASE MICRONS 1000 ;
END UNITS

MANUFACTURINGGRID 0.005 ;

LAYER li1
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.46 ;
  WIDTH 0.17 ;
END li1

LAYER mcon
  TYPE CUT ;
END mcon

LAYER met1
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.34 ;
  WIDTH 0.14 ;
END met1

LAYER via
  TYPE CUT ;
END via

LAYER met2
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.46 ;
  WIDTH 0.14 ;
END met2

LAYER via2
  TYPE CUT ;
END via2

LAYER met3
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.68 ;
  WIDTH 0.3 ;
END met3

LAYER via3
  TYPE CUT ;
END via3

LAYER met4
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.92 ;
  WIDTH 0.3 ;
END met4

LAYER via4
  TYPE CUT ;
END via4

LAYER met5
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 3.4 ;
  WIDTH 1.6 ;
END met5

LAYER nwell
  TYPE MASTERSLICE ;
END nwell

LAYER pwell
  TYPE MASTERSLICE ;
END pwell

LAYER OVERLAP
  TYPE OVERLAP ;
END OVERLAP

VIA L1M1_PR
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.145 -0.115 0.145 0.115 ;
END L1M1_PR

VIA L1M1_PR_R
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.115 -0.145 0.115 0.145 ;
END L1M1_PR_R

VIA L1M1_PR_M
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.115 -0.145 0.115 0.145 ;
END L1M1_PR_M

VIA L1M1_PR_MR
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.145 -0.115 0.145 0.115 ;
END L1M1_PR_MR

VIA L1M1_PR_C
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.145 -0.145 0.145 0.145 ;
END L1M1_PR_C

VIA M1M2_PR
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR

VIA M1M2_PR_Enc
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_Enc

VIA M1M2_PR_R
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_R

VIA M1M2_PR_R_Enc
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR_R_Enc

VIA M1M2_PR_M
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_M

VIA M1M2_PR_M_Enc
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR_M_Enc

VIA M1M2_PR_MR
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR_MR

VIA M1M2_PR_MR_Enc
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_MR_Enc

VIA M1M2_PR_C
  LAYER met1 ;
    RECT -0.16 -0.16 0.16 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.16 0.16 0.16 ;
END M1M2_PR_C

VIA M2M3_PR
  LAYER met2 ;
    RECT -0.14 -0.185 0.14 0.185 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR

VIA M2M3_PR_R
  LAYER met2 ;
    RECT -0.185 -0.14 0.185 0.14 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_R

VIA M2M3_PR_M
  LAYER met2 ;
    RECT -0.14 -0.185 0.14 0.185 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_M

VIA M2M3_PR_MR
  LAYER met2 ;
    RECT -0.185 -0.14 0.185 0.14 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_MR

VIA M2M3_PR_C
  LAYER met2 ;
    RECT -0.185 -0.185 0.185 0.185 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_C

VIA M3M4_PR
  LAYER met3 ;
    RECT -0.19 -0.16 0.19 0.16 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR

VIA M3M4_PR_R
  LAYER met3 ;
    RECT -0.16 -0.19 0.16 0.19 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_R

VIA M3M4_PR_M
  LAYER met3 ;
    RECT -0.19 -0.16 0.19 0.16 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_M

VIA M3M4_PR_MR
  LAYER met3 ;
    RECT -0.16 -0.19 0.16 0.19 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_MR

VIA M3M4_PR_C
  LAYER met3 ;
    RECT -0.19 -0.19 0.19 0.19 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_C

VIA M4M5_PR
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR

VIA M4M5_PR_R
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_R

VIA M4M5_PR_M
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_M

VIA M4M5_PR_MR
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_MR

VIA M4M5_PR_C
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_C

SITE unit
  CLASS CORE ;
  SYMMETRY Y ;
  SIZE 0.46 BY 2.72 ;
END unit

SITE unithddbl
  CLASS CORE ;
  SIZE 0.46 BY 5.44 ;
END unithddbl

MACRO cby_2__1_
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  SIZE 73.6 BY 119.68 ;
  SYMMETRY X Y ;
  PIN pReset[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 64.02 0.595 64.16 ;
    END
  END pReset[0]
  PIN chany_bottom_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.6 0 52.74 0.485 ;
    END
  END chany_bottom_in[0]
  PIN chany_bottom_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.52 0 53.66 0.485 ;
    END
  END chany_bottom_in[1]
  PIN chany_bottom_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.36 0 55.5 0.485 ;
    END
  END chany_bottom_in[2]
  PIN chany_bottom_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.44 0 54.58 0.485 ;
    END
  END chany_bottom_in[3]
  PIN chany_bottom_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.26 0 16.4 0.485 ;
    END
  END chany_bottom_in[4]
  PIN chany_bottom_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 6.75 0 7.05 0.8 ;
    END
  END chany_bottom_in[5]
  PIN chany_bottom_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.66 0 34.8 0.485 ;
    END
  END chany_bottom_in[6]
  PIN chany_bottom_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.42 0 14.56 0.485 ;
    END
  END chany_bottom_in[7]
  PIN chany_bottom_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.68 0 28.82 0.485 ;
    END
  END chany_bottom_in[8]
  PIN chany_bottom_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.26 0 62.4 0.485 ;
    END
  END chany_bottom_in[9]
  PIN chany_bottom_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.28 0 10.42 0.485 ;
    END
  END chany_bottom_in[10]
  PIN chany_bottom_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.58 0 35.72 0.485 ;
    END
  END chany_bottom_in[11]
  PIN chany_bottom_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.02 0 65.16 0.485 ;
    END
  END chany_bottom_in[12]
  PIN chany_bottom_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.34 0 15.48 0.485 ;
    END
  END chany_bottom_in[13]
  PIN chany_bottom_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.74 0 33.88 0.485 ;
    END
  END chany_bottom_in[14]
  PIN chany_bottom_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.08 0 24.22 0.485 ;
    END
  END chany_bottom_in[15]
  PIN chany_bottom_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.6 0 6.74 0.485 ;
    END
  END chany_bottom_in[16]
  PIN chany_bottom_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.86 0 44 0.485 ;
    END
  END chany_bottom_in[17]
  PIN chany_bottom_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.68 0 51.82 0.485 ;
    END
  END chany_bottom_in[18]
  PIN chany_bottom_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.94 0 20.08 0.485 ;
    END
  END chany_bottom_in[19]
  PIN chany_bottom_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.7 0 22.84 0.485 ;
    END
  END chany_bottom_in[20]
  PIN chany_bottom_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.56 0 18.7 0.485 ;
    END
  END chany_bottom_in[21]
  PIN chany_bottom_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.9 0 32.04 0.485 ;
    END
  END chany_bottom_in[22]
  PIN chany_bottom_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.5 0 36.64 0.485 ;
    END
  END chany_bottom_in[23]
  PIN chany_bottom_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.28 0 56.42 0.485 ;
    END
  END chany_bottom_in[24]
  PIN chany_bottom_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.64 0 17.78 0.485 ;
    END
  END chany_bottom_in[25]
  PIN chany_bottom_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.76 0 27.9 0.485 ;
    END
  END chany_bottom_in[26]
  PIN chany_bottom_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.78 0 21.92 0.485 ;
    END
  END chany_bottom_in[27]
  PIN chany_bottom_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.44 0 8.58 0.485 ;
    END
  END chany_bottom_in[28]
  PIN chany_bottom_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.08 0 47.22 0.485 ;
    END
  END chany_bottom_in[29]
  PIN chany_top_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.52 119.195 53.66 119.68 ;
    END
  END chany_top_in[0]
  PIN chany_top_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.94 119.195 43.08 119.68 ;
    END
  END chany_top_in[1]
  PIN chany_top_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.84 119.195 3.98 119.68 ;
    END
  END chany_top_in[2]
  PIN chany_top_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.6 119.195 52.74 119.68 ;
    END
  END chany_top_in[3]
  PIN chany_top_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.98 119.195 31.12 119.68 ;
    END
  END chany_top_in[4]
  PIN chany_top_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.94 119.195 66.08 119.68 ;
    END
  END chany_top_in[5]
  PIN chany_top_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.36 119.195 9.5 119.68 ;
    END
  END chany_top_in[6]
  PIN chany_top_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.26 119.195 16.4 119.68 ;
    END
  END chany_top_in[7]
  PIN chany_top_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.18 119.195 40.32 119.68 ;
    END
  END chany_top_in[8]
  PIN chany_top_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.3 119.195 27.44 119.68 ;
    END
  END chany_top_in[9]
  PIN chany_top_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.52 119.195 7.66 119.68 ;
    END
  END chany_top_in[10]
  PIN chany_top_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.5 119.195 36.64 119.68 ;
    END
  END chany_top_in[11]
  PIN chany_top_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.18 119.195 17.32 119.68 ;
    END
  END chany_top_in[12]
  PIN chany_top_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.1 119.195 18.24 119.68 ;
    END
  END chany_top_in[13]
  PIN chany_top_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.76 119.195 50.9 119.68 ;
    END
  END chany_top_in[14]
  PIN chany_top_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.62 119.195 23.76 119.68 ;
    END
  END chany_top_in[15]
  PIN chany_top_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.7 119.195 22.84 119.68 ;
    END
  END chany_top_in[16]
  PIN chany_top_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.16 119.195 46.3 119.68 ;
    END
  END chany_top_in[17]
  PIN chany_top_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.22 119.195 28.36 119.68 ;
    END
  END chany_top_in[18]
  PIN chany_top_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.94 119.195 20.08 119.68 ;
    END
  END chany_top_in[19]
  PIN chany_top_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.02 119.195 19.16 119.68 ;
    END
  END chany_top_in[20]
  PIN chany_top_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.78 119.195 21.92 119.68 ;
    END
  END chany_top_in[21]
  PIN chany_top_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.44 119.195 8.58 119.68 ;
    END
  END chany_top_in[22]
  PIN chany_top_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.34 119.195 38.48 119.68 ;
    END
  END chany_top_in[23]
  PIN chany_top_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.42 119.195 60.56 119.68 ;
    END
  END chany_top_in[24]
  PIN chany_top_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.36 119.195 55.5 119.68 ;
    END
  END chany_top_in[25]
  PIN chany_top_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.74 119.195 33.88 119.68 ;
    END
  END chany_top_in[26]
  PIN chany_top_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.38 119.195 26.52 119.68 ;
    END
  END chany_top_in[27]
  PIN chany_top_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.54 119.195 24.68 119.68 ;
    END
  END chany_top_in[28]
  PIN chany_top_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48 119.195 48.14 119.68 ;
    END
  END chany_top_in[29]
  PIN ccff_head[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 17.44 0.595 17.58 ;
    END
  END ccff_head[0]
  PIN chany_bottom_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.02 0 42.16 0.485 ;
    END
  END chany_bottom_out[0]
  PIN chany_bottom_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 30.67 0 30.97 0.8 ;
    END
  END chany_bottom_out[1]
  PIN chany_bottom_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.92 0 3.06 0.485 ;
    END
  END chany_bottom_out[2]
  PIN chany_bottom_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.84 0 26.98 0.485 ;
    END
  END chany_bottom_out[3]
  PIN chany_bottom_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.86 0 21 0.485 ;
    END
  END chany_bottom_out[4]
  PIN chany_bottom_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.98 0 31.12 0.485 ;
    END
  END chany_bottom_out[5]
  PIN chany_bottom_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25 0 25.14 0.485 ;
    END
  END chany_bottom_out[6]
  PIN chany_bottom_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.26 0 39.4 0.485 ;
    END
  END chany_bottom_out[7]
  PIN chany_bottom_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.94 0 43.08 0.485 ;
    END
  END chany_bottom_out[8]
  PIN chany_bottom_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.34 0 38.48 0.485 ;
    END
  END chany_bottom_out[9]
  PIN chany_bottom_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.42 0 60.56 0.485 ;
    END
  END chany_bottom_out[10]
  PIN chany_bottom_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48 0 48.14 0.485 ;
    END
  END chany_bottom_out[11]
  PIN chany_bottom_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.1 0 41.24 0.485 ;
    END
  END chany_bottom_out[12]
  PIN chany_bottom_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.42 0 37.56 0.485 ;
    END
  END chany_bottom_out[13]
  PIN chany_bottom_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.16 0 46.3 0.485 ;
    END
  END chany_bottom_out[14]
  PIN chany_bottom_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.1 0 64.24 0.485 ;
    END
  END chany_bottom_out[15]
  PIN chany_bottom_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.18 0 40.32 0.485 ;
    END
  END chany_bottom_out[16]
  PIN chany_bottom_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.5 0 59.64 0.485 ;
    END
  END chany_bottom_out[17]
  PIN chany_bottom_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.66 0 57.8 0.485 ;
    END
  END chany_bottom_out[18]
  PIN chany_bottom_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.18 0 63.32 0.485 ;
    END
  END chany_bottom_out[19]
  PIN chany_bottom_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.78 0 44.92 0.485 ;
    END
  END chany_bottom_out[20]
  PIN chany_bottom_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.92 0 26.06 0.485 ;
    END
  END chany_bottom_out[21]
  PIN chany_bottom_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.52 0 7.66 0.485 ;
    END
  END chany_bottom_out[22]
  PIN chany_bottom_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.5 0 13.64 0.485 ;
    END
  END chany_bottom_out[23]
  PIN chany_bottom_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.84 0 3.98 0.485 ;
    END
  END chany_bottom_out[24]
  PIN chany_bottom_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.58 0 12.72 0.485 ;
    END
  END chany_bottom_out[25]
  PIN chany_bottom_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.34 0 61.48 0.485 ;
    END
  END chany_bottom_out[26]
  PIN chany_bottom_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.76 0 50.9 0.485 ;
    END
  END chany_bottom_out[27]
  PIN chany_bottom_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.84 0 49.98 0.485 ;
    END
  END chany_bottom_out[28]
  PIN chany_bottom_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.92 0 49.06 0.485 ;
    END
  END chany_bottom_out[29]
  PIN chany_top_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.68 119.195 51.82 119.68 ;
    END
  END chany_top_out[0]
  PIN chany_top_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.68 119.195 5.82 119.68 ;
    END
  END chany_top_out[1]
  PIN chany_top_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.84 119.195 49.98 119.68 ;
    END
  END chany_top_out[2]
  PIN chany_top_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 24.23 118.88 24.53 119.68 ;
    END
  END chany_top_out[3]
  PIN chany_top_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.02 119.195 65.16 119.68 ;
    END
  END chany_top_out[4]
  PIN chany_top_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.32 119.195 44.46 119.68 ;
    END
  END chany_top_out[5]
  PIN chany_top_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.9 119.195 32.04 119.68 ;
    END
  END chany_top_out[6]
  PIN chany_top_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.1 119.195 41.24 119.68 ;
    END
  END chany_top_out[7]
  PIN chany_top_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.34 119.195 61.48 119.68 ;
    END
  END chany_top_out[8]
  PIN chany_top_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.66 119.195 34.8 119.68 ;
    END
  END chany_top_out[9]
  PIN chany_top_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.58 119.195 35.72 119.68 ;
    END
  END chany_top_out[10]
  PIN chany_top_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.08 119.195 47.22 119.68 ;
    END
  END chany_top_out[11]
  PIN chany_top_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.06 119.195 30.2 119.68 ;
    END
  END chany_top_out[12]
  PIN chany_top_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.1 119.195 64.24 119.68 ;
    END
  END chany_top_out[13]
  PIN chany_top_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.18 119.195 63.32 119.68 ;
    END
  END chany_top_out[14]
  PIN chany_top_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.28 119.195 56.42 119.68 ;
    END
  END chany_top_out[15]
  PIN chany_top_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.42 119.195 37.56 119.68 ;
    END
  END chany_top_out[16]
  PIN chany_top_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.24 119.195 45.38 119.68 ;
    END
  END chany_top_out[17]
  PIN chany_top_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.5 119.195 59.64 119.68 ;
    END
  END chany_top_out[18]
  PIN chany_top_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.26 119.195 39.4 119.68 ;
    END
  END chany_top_out[19]
  PIN chany_top_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.26 119.195 62.4 119.68 ;
    END
  END chany_top_out[20]
  PIN chany_top_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.92 119.195 49.06 119.68 ;
    END
  END chany_top_out[21]
  PIN chany_top_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.82 119.195 32.96 119.68 ;
    END
  END chany_top_out[22]
  PIN chany_top_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 30.67 118.88 30.97 119.68 ;
    END
  END chany_top_out[23]
  PIN chany_top_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.76 119.195 4.9 119.68 ;
    END
  END chany_top_out[24]
  PIN chany_top_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.66 119.195 57.8 119.68 ;
    END
  END chany_top_out[25]
  PIN chany_top_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.46 119.195 25.6 119.68 ;
    END
  END chany_top_out[26]
  PIN chany_top_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.86 119.195 21 119.68 ;
    END
  END chany_top_out[27]
  PIN chany_top_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.02 119.195 42.16 119.68 ;
    END
  END chany_top_out[28]
  PIN chany_top_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.44 119.195 54.58 119.68 ;
    END
  END chany_top_out[29]
  PIN right_grid_pin_0_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 39.87 0 40.17 0.8 ;
    END
  END right_grid_pin_0_[0]
  PIN left_grid_pin_16_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 63.34 0.595 63.48 ;
    END
  END left_grid_pin_16_[0]
  PIN left_grid_pin_17_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 105.16 0.595 105.3 ;
    END
  END left_grid_pin_17_[0]
  PIN left_grid_pin_18_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 83.4 0.595 83.54 ;
    END
  END left_grid_pin_18_[0]
  PIN left_grid_pin_19_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 85.1 0.595 85.24 ;
    END
  END left_grid_pin_19_[0]
  PIN left_grid_pin_20_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 41.58 0.595 41.72 ;
    END
  END left_grid_pin_20_[0]
  PIN left_grid_pin_21_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 39.88 0.595 40.02 ;
    END
  END left_grid_pin_21_[0]
  PIN left_grid_pin_22_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 42.26 0.595 42.4 ;
    END
  END left_grid_pin_22_[0]
  PIN left_grid_pin_23_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 61.64 0.595 61.78 ;
    END
  END left_grid_pin_23_[0]
  PIN left_grid_pin_24_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 37.16 0.595 37.3 ;
    END
  END left_grid_pin_24_[0]
  PIN left_grid_pin_25_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 60.96 0.595 61.1 ;
    END
  END left_grid_pin_25_[0]
  PIN left_grid_pin_26_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 19.82 0.595 19.96 ;
    END
  END left_grid_pin_26_[0]
  PIN left_grid_pin_27_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 39.2 0.595 39.34 ;
    END
  END left_grid_pin_27_[0]
  PIN left_grid_pin_28_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 4.52 0.595 4.66 ;
    END
  END left_grid_pin_28_[0]
  PIN left_grid_pin_29_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 3.84 0.595 3.98 ;
    END
  END left_grid_pin_29_[0]
  PIN left_grid_pin_30_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 18.12 0.595 18.26 ;
    END
  END left_grid_pin_30_[0]
  PIN left_grid_pin_31_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 20.5 0.595 20.64 ;
    END
  END left_grid_pin_31_[0]
  PIN ccff_tail[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.36 0 9.5 0.485 ;
    END
  END ccff_tail[0]
  PIN IO_ISOL_N[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 6.22 0.595 6.36 ;
    END
  END IO_ISOL_N[0]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 73.005 1.8 73.6 1.94 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[0]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 73.005 4.52 73.6 4.66 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[0]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 73.005 3.5 73.6 3.64 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[0]
  PIN left_width_0_height_0__pin_0_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 38.03 0 38.33 0.8 ;
    END
  END left_width_0_height_0__pin_0_[0]
  PIN left_width_0_height_0__pin_1_upper[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.46 119.195 2.6 119.68 ;
    END
  END left_width_0_height_0__pin_1_upper[0]
  PIN left_width_0_height_0__pin_1_lower[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.82 0 32.96 0.485 ;
    END
  END left_width_0_height_0__pin_1_lower[0]
  PIN pReset_S_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.22 0 5.36 0.485 ;
    END
  END pReset_S_in
  PIN prog_clk_0_W_in
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER met1 ;
        RECT 0 1.8 0.595 1.94 ;
    END
  END prog_clk_0_W_in
  PIN prog_clk_0_S_out
    DIRECTION OUTPUT ;
    USE CLOCK ;
    PORT
      LAYER met2 ;
        RECT 11.66 0 11.8 0.485 ;
    END
  END prog_clk_0_S_out
  PIN prog_clk_0_N_out
    DIRECTION OUTPUT ;
    USE CLOCK ;
    PORT
      LAYER met2 ;
        RECT 6.6 119.195 6.74 119.68 ;
    END
  END prog_clk_0_N_out
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0 7.24 3.2 10.44 ;
        RECT 70.4 7.24 73.6 10.44 ;
        RECT 0 48.04 3.2 51.24 ;
        RECT 70.4 48.04 73.6 51.24 ;
        RECT 0 88.84 3.2 92.04 ;
        RECT 70.4 88.84 73.6 92.04 ;
      LAYER met4 ;
        RECT 14.42 0 15.02 0.6 ;
        RECT 43.86 0 44.46 0.6 ;
        RECT 14.42 119.08 15.02 119.68 ;
        RECT 43.86 119.08 44.46 119.68 ;
      LAYER met1 ;
        RECT 0 2.48 0.48 2.96 ;
        RECT 73.12 2.48 73.6 2.96 ;
        RECT 0 7.92 0.48 8.4 ;
        RECT 73.12 7.92 73.6 8.4 ;
        RECT 0 13.36 0.48 13.84 ;
        RECT 73.12 13.36 73.6 13.84 ;
        RECT 0 18.8 0.48 19.28 ;
        RECT 73.12 18.8 73.6 19.28 ;
        RECT 0 24.24 0.48 24.72 ;
        RECT 73.12 24.24 73.6 24.72 ;
        RECT 0 29.68 0.48 30.16 ;
        RECT 73.12 29.68 73.6 30.16 ;
        RECT 0 35.12 0.48 35.6 ;
        RECT 73.12 35.12 73.6 35.6 ;
        RECT 0 40.56 0.48 41.04 ;
        RECT 73.12 40.56 73.6 41.04 ;
        RECT 0 46 0.48 46.48 ;
        RECT 73.12 46 73.6 46.48 ;
        RECT 0 51.44 0.48 51.92 ;
        RECT 73.12 51.44 73.6 51.92 ;
        RECT 0 56.88 0.48 57.36 ;
        RECT 73.12 56.88 73.6 57.36 ;
        RECT 0 62.32 0.48 62.8 ;
        RECT 73.12 62.32 73.6 62.8 ;
        RECT 0 67.76 0.48 68.24 ;
        RECT 73.12 67.76 73.6 68.24 ;
        RECT 0 73.2 0.48 73.68 ;
        RECT 73.12 73.2 73.6 73.68 ;
        RECT 0 78.64 0.48 79.12 ;
        RECT 73.12 78.64 73.6 79.12 ;
        RECT 0 84.08 0.48 84.56 ;
        RECT 73.12 84.08 73.6 84.56 ;
        RECT 0 89.52 0.48 90 ;
        RECT 73.12 89.52 73.6 90 ;
        RECT 0 94.96 0.48 95.44 ;
        RECT 73.12 94.96 73.6 95.44 ;
        RECT 0 100.4 0.48 100.88 ;
        RECT 73.12 100.4 73.6 100.88 ;
        RECT 0 105.84 0.48 106.32 ;
        RECT 73.12 105.84 73.6 106.32 ;
        RECT 0 111.28 0.48 111.76 ;
        RECT 73.12 111.28 73.6 111.76 ;
        RECT 0 116.72 0.48 117.2 ;
        RECT 73.12 116.72 73.6 117.2 ;
    END
  END VDD
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0 27.64 3.2 30.84 ;
        RECT 70.4 27.64 73.6 30.84 ;
        RECT 0 68.44 3.2 71.64 ;
        RECT 70.4 68.44 73.6 71.64 ;
        RECT 0 109.24 3.2 112.44 ;
        RECT 70.4 109.24 73.6 112.44 ;
      LAYER met4 ;
        RECT 29.14 0 29.74 0.6 ;
        RECT 58.58 0 59.18 0.6 ;
        RECT 29.14 119.08 29.74 119.68 ;
        RECT 58.58 119.08 59.18 119.68 ;
      LAYER met1 ;
        RECT 0 -0.24 0.48 0.24 ;
        RECT 73.12 -0.24 73.6 0.24 ;
        RECT 0 5.2 0.48 5.68 ;
        RECT 73.12 5.2 73.6 5.68 ;
        RECT 0 10.64 0.48 11.12 ;
        RECT 73.12 10.64 73.6 11.12 ;
        RECT 0 16.08 0.48 16.56 ;
        RECT 73.12 16.08 73.6 16.56 ;
        RECT 0 21.52 0.48 22 ;
        RECT 73.12 21.52 73.6 22 ;
        RECT 0 26.96 0.48 27.44 ;
        RECT 73.12 26.96 73.6 27.44 ;
        RECT 0 32.4 0.48 32.88 ;
        RECT 73.12 32.4 73.6 32.88 ;
        RECT 0 37.84 0.48 38.32 ;
        RECT 73.12 37.84 73.6 38.32 ;
        RECT 0 43.28 0.48 43.76 ;
        RECT 73.12 43.28 73.6 43.76 ;
        RECT 0 48.72 0.48 49.2 ;
        RECT 73.12 48.72 73.6 49.2 ;
        RECT 0 54.16 0.48 54.64 ;
        RECT 73.12 54.16 73.6 54.64 ;
        RECT 0 59.6 0.48 60.08 ;
        RECT 73.12 59.6 73.6 60.08 ;
        RECT 0 65.04 0.48 65.52 ;
        RECT 73.12 65.04 73.6 65.52 ;
        RECT 0 70.48 0.48 70.96 ;
        RECT 73.12 70.48 73.6 70.96 ;
        RECT 0 75.92 0.48 76.4 ;
        RECT 73.12 75.92 73.6 76.4 ;
        RECT 0 81.36 0.48 81.84 ;
        RECT 73.12 81.36 73.6 81.84 ;
        RECT 0 86.8 0.48 87.28 ;
        RECT 73.12 86.8 73.6 87.28 ;
        RECT 0 92.24 0.48 92.72 ;
        RECT 73.12 92.24 73.6 92.72 ;
        RECT 0 97.68 0.48 98.16 ;
        RECT 73.12 97.68 73.6 98.16 ;
        RECT 0 103.12 0.48 103.6 ;
        RECT 73.12 103.12 73.6 103.6 ;
        RECT 0 108.56 0.48 109.04 ;
        RECT 73.12 108.56 73.6 109.04 ;
        RECT 0 114 0.48 114.48 ;
        RECT 73.12 114 73.6 114.48 ;
        RECT 0 119.44 0.48 119.92 ;
        RECT 73.12 119.44 73.6 119.92 ;
    END
  END VSS
  OBS
    LAYER met1 ;
      POLYGON 72.84 119.92 72.84 119.44 59.04 119.44 59.04 119.43 58.72 119.43 58.72 119.44 29.6 119.44 29.6 119.43 29.28 119.43 29.28 119.44 0.76 119.44 0.76 119.92 ;
      POLYGON 59.04 0.25 59.04 0.24 72.84 0.24 72.84 -0.24 0.76 -0.24 0.76 0.24 29.28 0.24 29.28 0.25 29.6 0.25 29.6 0.24 58.72 0.24 58.72 0.25 ;
      POLYGON 72.84 119.4 72.84 119.16 73.32 119.16 73.32 117.48 72.84 117.48 72.84 116.44 73.32 116.44 73.32 114.76 72.84 114.76 72.84 113.72 73.32 113.72 73.32 112.04 72.84 112.04 72.84 111 73.32 111 73.32 109.32 72.84 109.32 72.84 108.28 73.32 108.28 73.32 106.6 72.84 106.6 72.84 105.56 73.32 105.56 73.32 103.88 72.84 103.88 72.84 102.84 73.32 102.84 73.32 101.16 72.84 101.16 72.84 100.12 73.32 100.12 73.32 98.44 72.84 98.44 72.84 97.4 73.32 97.4 73.32 95.72 72.84 95.72 72.84 94.68 73.32 94.68 73.32 93 72.84 93 72.84 91.96 73.32 91.96 73.32 90.28 72.84 90.28 72.84 89.24 73.32 89.24 73.32 87.56 72.84 87.56 72.84 86.52 73.32 86.52 73.32 84.84 72.84 84.84 72.84 83.8 73.32 83.8 73.32 82.12 72.84 82.12 72.84 81.08 73.32 81.08 73.32 79.4 72.84 79.4 72.84 78.36 73.32 78.36 73.32 76.68 72.84 76.68 72.84 75.64 73.32 75.64 73.32 73.96 72.84 73.96 72.84 72.92 73.32 72.92 73.32 71.24 72.84 71.24 72.84 70.2 73.32 70.2 73.32 68.52 72.84 68.52 72.84 67.48 73.32 67.48 73.32 65.8 72.84 65.8 72.84 64.76 73.32 64.76 73.32 63.08 72.84 63.08 72.84 62.04 73.32 62.04 73.32 60.36 72.84 60.36 72.84 59.32 73.32 59.32 73.32 57.64 72.84 57.64 72.84 56.6 73.32 56.6 73.32 54.92 72.84 54.92 72.84 53.88 73.32 53.88 73.32 52.2 72.84 52.2 72.84 51.16 73.32 51.16 73.32 49.48 72.84 49.48 72.84 48.44 73.32 48.44 73.32 46.76 72.84 46.76 72.84 45.72 73.32 45.72 73.32 44.04 72.84 44.04 72.84 43 73.32 43 73.32 41.32 72.84 41.32 72.84 40.28 73.32 40.28 73.32 38.6 72.84 38.6 72.84 37.56 73.32 37.56 73.32 35.88 72.84 35.88 72.84 34.84 73.32 34.84 73.32 33.16 72.84 33.16 72.84 32.12 73.32 32.12 73.32 30.44 72.84 30.44 72.84 29.4 73.32 29.4 73.32 27.72 72.84 27.72 72.84 26.68 73.32 26.68 73.32 25 72.84 25 72.84 23.96 73.32 23.96 73.32 22.28 72.84 22.28 72.84 21.24 73.32 21.24 73.32 19.56 72.84 19.56 72.84 18.52 73.32 18.52 73.32 16.84 72.84 16.84 72.84 15.8 73.32 15.8 73.32 14.12 72.84 14.12 72.84 13.08 73.32 13.08 73.32 11.4 72.84 11.4 72.84 10.36 73.32 10.36 73.32 8.68 72.84 8.68 72.84 7.64 73.32 7.64 73.32 5.96 72.84 5.96 72.84 4.94 72.725 4.94 72.725 4.24 73.32 4.24 73.32 3.92 72.725 3.92 72.725 3.22 72.84 3.22 72.84 2.22 72.725 2.22 72.725 1.52 73.32 1.52 73.32 0.52 72.84 0.52 72.84 0.28 0.76 0.28 0.76 0.52 0.28 0.52 0.28 1.52 0.875 1.52 0.875 2.22 0.76 2.22 0.76 3.24 0.28 3.24 0.28 3.56 0.875 3.56 0.875 4.94 0.76 4.94 0.76 5.94 0.875 5.94 0.875 6.64 0.28 6.64 0.28 7.64 0.76 7.64 0.76 8.68 0.28 8.68 0.28 10.36 0.76 10.36 0.76 11.4 0.28 11.4 0.28 13.08 0.76 13.08 0.76 14.12 0.28 14.12 0.28 15.8 0.76 15.8 0.76 16.84 0.28 16.84 0.28 17.16 0.875 17.16 0.875 18.54 0.76 18.54 0.76 19.54 0.875 19.54 0.875 20.92 0.28 20.92 0.28 21.24 0.76 21.24 0.76 22.28 0.28 22.28 0.28 23.96 0.76 23.96 0.76 25 0.28 25 0.28 26.68 0.76 26.68 0.76 27.72 0.28 27.72 0.28 29.4 0.76 29.4 0.76 30.44 0.28 30.44 0.28 32.12 0.76 32.12 0.76 33.16 0.28 33.16 0.28 34.84 0.76 34.84 0.76 35.88 0.28 35.88 0.28 36.88 0.875 36.88 0.875 37.58 0.76 37.58 0.76 38.6 0.28 38.6 0.28 38.92 0.875 38.92 0.875 40.3 0.76 40.3 0.76 41.3 0.875 41.3 0.875 42.68 0.28 42.68 0.28 43 0.76 43 0.76 44.04 0.28 44.04 0.28 45.72 0.76 45.72 0.76 46.76 0.28 46.76 0.28 48.44 0.76 48.44 0.76 49.48 0.28 49.48 0.28 51.16 0.76 51.16 0.76 52.2 0.28 52.2 0.28 53.88 0.76 53.88 0.76 54.92 0.28 54.92 0.28 56.6 0.76 56.6 0.76 57.64 0.28 57.64 0.28 59.32 0.76 59.32 0.76 60.36 0.28 60.36 0.28 60.68 0.875 60.68 0.875 62.06 0.76 62.06 0.76 63.06 0.875 63.06 0.875 64.44 0.28 64.44 0.28 64.76 0.76 64.76 0.76 65.8 0.28 65.8 0.28 67.48 0.76 67.48 0.76 68.52 0.28 68.52 0.28 70.2 0.76 70.2 0.76 71.24 0.28 71.24 0.28 72.92 0.76 72.92 0.76 73.96 0.28 73.96 0.28 75.64 0.76 75.64 0.76 76.68 0.28 76.68 0.28 78.36 0.76 78.36 0.76 79.4 0.28 79.4 0.28 81.08 0.76 81.08 0.76 82.12 0.28 82.12 0.28 83.12 0.875 83.12 0.875 83.82 0.76 83.82 0.76 84.82 0.875 84.82 0.875 85.52 0.28 85.52 0.28 86.52 0.76 86.52 0.76 87.56 0.28 87.56 0.28 89.24 0.76 89.24 0.76 90.28 0.28 90.28 0.28 91.96 0.76 91.96 0.76 93 0.28 93 0.28 94.68 0.76 94.68 0.76 95.72 0.28 95.72 0.28 97.4 0.76 97.4 0.76 98.44 0.28 98.44 0.28 100.12 0.76 100.12 0.76 101.16 0.28 101.16 0.28 102.84 0.76 102.84 0.76 103.88 0.28 103.88 0.28 104.88 0.875 104.88 0.875 105.58 0.76 105.58 0.76 106.6 0.28 106.6 0.28 108.28 0.76 108.28 0.76 109.32 0.28 109.32 0.28 111 0.76 111 0.76 112.04 0.28 112.04 0.28 113.72 0.76 113.72 0.76 114.76 0.28 114.76 0.28 116.44 0.76 116.44 0.76 117.48 0.28 117.48 0.28 119.16 0.76 119.16 0.76 119.4 ;
    LAYER met2 ;
      RECT 58.74 119.375 59.02 119.745 ;
      RECT 29.3 119.375 29.58 119.745 ;
      POLYGON 44.92 119.58 44.92 112.47 44.78 112.47 44.78 119.44 44.74 119.44 44.74 119.58 ;
      POLYGON 10.42 119.58 10.42 115.36 10.28 115.36 10.28 119.44 9.78 119.44 9.78 119.58 ;
      RECT 24.02 119.01 24.28 119.33 ;
      POLYGON 4.9 9.25 4.9 0.1 4.26 0.1 4.26 0.24 4.76 0.24 4.76 9.25 ;
      RECT 38.74 0.69 39 1.01 ;
      RECT 51.16 0.35 51.42 0.67 ;
      RECT 41.5 0.35 41.76 0.67 ;
      RECT 58.74 -0.065 59.02 0.305 ;
      RECT 29.3 -0.065 29.58 0.305 ;
      POLYGON 73.32 119.4 73.32 0.28 65.44 0.28 65.44 0.765 64.74 0.765 64.74 0.28 64.52 0.28 64.52 0.765 63.82 0.765 63.82 0.28 63.6 0.28 63.6 0.765 62.9 0.765 62.9 0.28 62.68 0.28 62.68 0.765 61.98 0.765 61.98 0.28 61.76 0.28 61.76 0.765 61.06 0.765 61.06 0.28 60.84 0.28 60.84 0.765 60.14 0.765 60.14 0.28 59.92 0.28 59.92 0.765 59.22 0.765 59.22 0.28 58.08 0.28 58.08 0.765 57.38 0.765 57.38 0.28 56.7 0.28 56.7 0.765 56 0.765 56 0.28 55.78 0.28 55.78 0.765 55.08 0.765 55.08 0.28 54.86 0.28 54.86 0.765 54.16 0.765 54.16 0.28 53.94 0.28 53.94 0.765 53.24 0.765 53.24 0.28 53.02 0.28 53.02 0.765 52.32 0.765 52.32 0.28 52.1 0.28 52.1 0.765 51.4 0.765 51.4 0.28 51.18 0.28 51.18 0.765 50.48 0.765 50.48 0.28 50.26 0.28 50.26 0.765 49.56 0.765 49.56 0.28 49.34 0.28 49.34 0.765 48.64 0.765 48.64 0.28 48.42 0.28 48.42 0.765 47.72 0.765 47.72 0.28 47.5 0.28 47.5 0.765 46.8 0.765 46.8 0.28 46.58 0.28 46.58 0.765 45.88 0.765 45.88 0.28 45.2 0.28 45.2 0.765 44.5 0.765 44.5 0.28 44.28 0.28 44.28 0.765 43.58 0.765 43.58 0.28 43.36 0.28 43.36 0.765 42.66 0.765 42.66 0.28 42.44 0.28 42.44 0.765 41.74 0.765 41.74 0.28 41.52 0.28 41.52 0.765 40.82 0.765 40.82 0.28 40.6 0.28 40.6 0.765 39.9 0.765 39.9 0.28 39.68 0.28 39.68 0.765 38.98 0.765 38.98 0.28 38.76 0.28 38.76 0.765 38.06 0.765 38.06 0.28 37.84 0.28 37.84 0.765 37.14 0.765 37.14 0.28 36.92 0.28 36.92 0.765 36.22 0.765 36.22 0.28 36 0.28 36 0.765 35.3 0.765 35.3 0.28 35.08 0.28 35.08 0.765 34.38 0.765 34.38 0.28 34.16 0.28 34.16 0.765 33.46 0.765 33.46 0.28 33.24 0.28 33.24 0.765 32.54 0.765 32.54 0.28 32.32 0.28 32.32 0.765 31.62 0.765 31.62 0.28 31.4 0.28 31.4 0.765 30.7 0.765 30.7 0.28 29.1 0.28 29.1 0.765 28.4 0.765 28.4 0.28 28.18 0.28 28.18 0.765 27.48 0.765 27.48 0.28 27.26 0.28 27.26 0.765 26.56 0.765 26.56 0.28 26.34 0.28 26.34 0.765 25.64 0.765 25.64 0.28 25.42 0.28 25.42 0.765 24.72 0.765 24.72 0.28 24.5 0.28 24.5 0.765 23.8 0.765 23.8 0.28 23.12 0.28 23.12 0.765 22.42 0.765 22.42 0.28 22.2 0.28 22.2 0.765 21.5 0.765 21.5 0.28 21.28 0.28 21.28 0.765 20.58 0.765 20.58 0.28 20.36 0.28 20.36 0.765 19.66 0.765 19.66 0.28 18.98 0.28 18.98 0.765 18.28 0.765 18.28 0.28 18.06 0.28 18.06 0.765 17.36 0.765 17.36 0.28 16.68 0.28 16.68 0.765 15.98 0.765 15.98 0.28 15.76 0.28 15.76 0.765 15.06 0.765 15.06 0.28 14.84 0.28 14.84 0.765 14.14 0.765 14.14 0.28 13.92 0.28 13.92 0.765 13.22 0.765 13.22 0.28 13 0.28 13 0.765 12.3 0.765 12.3 0.28 12.08 0.28 12.08 0.765 11.38 0.765 11.38 0.28 10.7 0.28 10.7 0.765 10 0.765 10 0.28 9.78 0.28 9.78 0.765 9.08 0.765 9.08 0.28 8.86 0.28 8.86 0.765 8.16 0.765 8.16 0.28 7.94 0.28 7.94 0.765 7.24 0.765 7.24 0.28 7.02 0.28 7.02 0.765 6.32 0.765 6.32 0.28 5.64 0.28 5.64 0.765 4.94 0.765 4.94 0.28 4.26 0.28 4.26 0.765 3.56 0.765 3.56 0.28 3.34 0.28 3.34 0.765 2.64 0.765 2.64 0.28 0.28 0.28 0.28 119.4 2.18 119.4 2.18 118.915 2.88 118.915 2.88 119.4 3.56 119.4 3.56 118.915 4.26 118.915 4.26 119.4 4.48 119.4 4.48 118.915 5.18 118.915 5.18 119.4 5.4 119.4 5.4 118.915 6.1 118.915 6.1 119.4 6.32 119.4 6.32 118.915 7.02 118.915 7.02 119.4 7.24 119.4 7.24 118.915 7.94 118.915 7.94 119.4 8.16 119.4 8.16 118.915 8.86 118.915 8.86 119.4 9.08 119.4 9.08 118.915 9.78 118.915 9.78 119.4 15.98 119.4 15.98 118.915 16.68 118.915 16.68 119.4 16.9 119.4 16.9 118.915 17.6 118.915 17.6 119.4 17.82 119.4 17.82 118.915 18.52 118.915 18.52 119.4 18.74 119.4 18.74 118.915 19.44 118.915 19.44 119.4 19.66 119.4 19.66 118.915 20.36 118.915 20.36 119.4 20.58 119.4 20.58 118.915 21.28 118.915 21.28 119.4 21.5 119.4 21.5 118.915 22.2 118.915 22.2 119.4 22.42 119.4 22.42 118.915 23.12 118.915 23.12 119.4 23.34 119.4 23.34 118.915 24.04 118.915 24.04 119.4 24.26 119.4 24.26 118.915 24.96 118.915 24.96 119.4 25.18 119.4 25.18 118.915 25.88 118.915 25.88 119.4 26.1 119.4 26.1 118.915 26.8 118.915 26.8 119.4 27.02 119.4 27.02 118.915 27.72 118.915 27.72 119.4 27.94 119.4 27.94 118.915 28.64 118.915 28.64 119.4 29.78 119.4 29.78 118.915 30.48 118.915 30.48 119.4 30.7 119.4 30.7 118.915 31.4 118.915 31.4 119.4 31.62 119.4 31.62 118.915 32.32 118.915 32.32 119.4 32.54 119.4 32.54 118.915 33.24 118.915 33.24 119.4 33.46 119.4 33.46 118.915 34.16 118.915 34.16 119.4 34.38 119.4 34.38 118.915 35.08 118.915 35.08 119.4 35.3 119.4 35.3 118.915 36 118.915 36 119.4 36.22 119.4 36.22 118.915 36.92 118.915 36.92 119.4 37.14 119.4 37.14 118.915 37.84 118.915 37.84 119.4 38.06 119.4 38.06 118.915 38.76 118.915 38.76 119.4 38.98 119.4 38.98 118.915 39.68 118.915 39.68 119.4 39.9 119.4 39.9 118.915 40.6 118.915 40.6 119.4 40.82 119.4 40.82 118.915 41.52 118.915 41.52 119.4 41.74 119.4 41.74 118.915 42.44 118.915 42.44 119.4 42.66 119.4 42.66 118.915 43.36 118.915 43.36 119.4 44.04 119.4 44.04 118.915 44.74 118.915 44.74 119.4 44.96 119.4 44.96 118.915 45.66 118.915 45.66 119.4 45.88 119.4 45.88 118.915 46.58 118.915 46.58 119.4 46.8 119.4 46.8 118.915 47.5 118.915 47.5 119.4 47.72 119.4 47.72 118.915 48.42 118.915 48.42 119.4 48.64 119.4 48.64 118.915 49.34 118.915 49.34 119.4 49.56 119.4 49.56 118.915 50.26 118.915 50.26 119.4 50.48 119.4 50.48 118.915 51.18 118.915 51.18 119.4 51.4 119.4 51.4 118.915 52.1 118.915 52.1 119.4 52.32 119.4 52.32 118.915 53.02 118.915 53.02 119.4 53.24 119.4 53.24 118.915 53.94 118.915 53.94 119.4 54.16 119.4 54.16 118.915 54.86 118.915 54.86 119.4 55.08 119.4 55.08 118.915 55.78 118.915 55.78 119.4 56 119.4 56 118.915 56.7 118.915 56.7 119.4 57.38 119.4 57.38 118.915 58.08 118.915 58.08 119.4 59.22 119.4 59.22 118.915 59.92 118.915 59.92 119.4 60.14 119.4 60.14 118.915 60.84 118.915 60.84 119.4 61.06 119.4 61.06 118.915 61.76 118.915 61.76 119.4 61.98 119.4 61.98 118.915 62.68 118.915 62.68 119.4 62.9 119.4 62.9 118.915 63.6 118.915 63.6 119.4 63.82 119.4 63.82 118.915 64.52 118.915 64.52 119.4 64.74 119.4 64.74 118.915 65.44 118.915 65.44 119.4 65.66 119.4 65.66 118.915 66.36 118.915 66.36 119.4 ;
    LAYER met4 ;
      POLYGON 36.505 119.505 36.505 119.175 36.49 119.175 36.49 87.91 36.19 87.91 36.19 119.175 36.175 119.175 36.175 119.505 ;
      POLYGON 26.385 119.505 26.385 119.175 26.37 119.175 26.37 83.83 26.07 83.83 26.07 119.175 26.055 119.175 26.055 119.505 ;
      POLYGON 73.2 119.28 73.2 0.4 59.58 0.4 59.58 1 58.18 1 58.18 0.4 44.86 0.4 44.86 1 43.46 1 43.46 0.4 40.57 0.4 40.57 1.2 39.47 1.2 39.47 0.4 38.73 0.4 38.73 1.2 37.63 1.2 37.63 0.4 31.37 0.4 31.37 1.2 30.27 1.2 30.27 0.4 30.14 0.4 30.14 1 28.74 1 28.74 0.4 15.42 0.4 15.42 1 14.02 1 14.02 0.4 7.45 0.4 7.45 1.2 6.35 1.2 6.35 0.4 0.4 0.4 0.4 119.28 14.02 119.28 14.02 118.68 15.42 118.68 15.42 119.28 23.83 119.28 23.83 118.48 24.93 118.48 24.93 119.28 28.74 119.28 28.74 118.68 30.14 118.68 30.14 119.28 30.27 119.28 30.27 118.48 31.37 118.48 31.37 119.28 43.46 119.28 43.46 118.68 44.86 118.68 44.86 119.28 58.18 119.28 58.18 118.68 59.58 118.68 59.58 119.28 ;
    LAYER met5 ;
      POLYGON 72 118.08 72 114.04 68.8 114.04 68.8 107.64 72 107.64 72 93.64 68.8 93.64 68.8 87.24 72 87.24 72 73.24 68.8 73.24 68.8 66.84 72 66.84 72 52.84 68.8 52.84 68.8 46.44 72 46.44 72 32.44 68.8 32.44 68.8 26.04 72 26.04 72 12.04 68.8 12.04 68.8 5.64 72 5.64 72 1.6 1.6 1.6 1.6 5.64 4.8 5.64 4.8 12.04 1.6 12.04 1.6 26.04 4.8 26.04 4.8 32.44 1.6 32.44 1.6 46.44 4.8 46.44 4.8 52.84 1.6 52.84 1.6 66.84 4.8 66.84 4.8 73.24 1.6 73.24 1.6 87.24 4.8 87.24 4.8 93.64 1.6 93.64 1.6 107.64 4.8 107.64 4.8 114.04 1.6 114.04 1.6 118.08 ;
    LAYER li1 ;
      POLYGON 73.6 119.765 73.6 119.595 69.905 119.595 69.905 118.795 69.575 118.795 69.575 119.595 69.065 119.595 69.065 119.115 68.735 119.115 68.735 119.595 68.225 119.595 68.225 119.115 67.895 119.115 67.895 119.595 67.385 119.595 67.385 119.115 67.055 119.115 67.055 119.595 66.545 119.595 66.545 119.115 66.215 119.115 66.215 119.595 65.705 119.595 65.705 119.115 65.375 119.115 65.375 119.595 63.925 119.595 63.925 118.795 63.595 118.795 63.595 119.595 63.085 119.595 63.085 119.115 62.755 119.115 62.755 119.595 62.245 119.595 62.245 119.115 61.915 119.115 61.915 119.595 61.405 119.595 61.405 119.115 61.075 119.115 61.075 119.595 60.565 119.595 60.565 119.115 60.235 119.115 60.235 119.595 59.725 119.595 59.725 119.115 59.395 119.115 59.395 119.595 57.485 119.595 57.485 118.795 57.155 118.795 57.155 119.595 56.645 119.595 56.645 119.115 56.315 119.115 56.315 119.595 55.805 119.595 55.805 119.115 55.475 119.115 55.475 119.595 54.965 119.595 54.965 119.115 54.635 119.115 54.635 119.595 54.125 119.595 54.125 119.115 53.795 119.115 53.795 119.595 53.285 119.595 53.285 119.115 52.955 119.115 52.955 119.595 51.465 119.595 51.465 119.115 51.135 119.115 51.135 119.595 50.625 119.595 50.625 119.115 50.295 119.115 50.295 119.595 49.785 119.595 49.785 119.115 49.455 119.115 49.455 119.595 48.945 119.595 48.945 119.115 48.615 119.115 48.615 119.595 48.105 119.595 48.105 119.115 47.775 119.115 47.775 119.595 47.265 119.595 47.265 118.795 46.935 118.795 46.935 119.595 45.065 119.595 45.065 118.795 44.735 118.795 44.735 119.595 44.225 119.595 44.225 119.115 43.895 119.115 43.895 119.595 43.385 119.595 43.385 119.115 43.055 119.115 43.055 119.595 42.545 119.595 42.545 119.115 42.215 119.115 42.215 119.595 41.705 119.595 41.705 119.115 41.375 119.115 41.375 119.595 40.865 119.595 40.865 119.115 40.535 119.115 40.535 119.595 39.085 119.595 39.085 118.795 38.755 118.795 38.755 119.595 38.245 119.595 38.245 119.115 37.915 119.115 37.915 119.595 37.405 119.595 37.405 119.115 37.075 119.115 37.075 119.595 36.565 119.595 36.565 119.115 36.235 119.115 36.235 119.595 35.725 119.595 35.725 119.115 35.395 119.115 35.395 119.595 34.885 119.595 34.885 119.115 34.555 119.115 34.555 119.595 32.645 119.595 32.645 118.795 32.315 118.795 32.315 119.595 31.805 119.595 31.805 119.115 31.475 119.115 31.475 119.595 30.965 119.595 30.965 119.115 30.635 119.115 30.635 119.595 30.125 119.595 30.125 119.115 29.795 119.115 29.795 119.595 29.285 119.595 29.285 119.115 28.955 119.115 28.955 119.595 28.445 119.595 28.445 119.115 28.115 119.115 28.115 119.595 26.665 119.595 26.665 118.795 26.335 118.795 26.335 119.595 25.825 119.595 25.825 119.115 25.495 119.115 25.495 119.595 24.985 119.595 24.985 119.115 24.655 119.115 24.655 119.595 24.145 119.595 24.145 119.115 23.815 119.115 23.815 119.595 23.305 119.595 23.305 119.115 22.975 119.115 22.975 119.595 22.465 119.595 22.465 119.115 22.135 119.115 22.135 119.595 20.225 119.595 20.225 118.795 19.895 118.795 19.895 119.595 19.385 119.595 19.385 119.115 19.055 119.115 19.055 119.595 18.545 119.595 18.545 119.115 18.215 119.115 18.215 119.595 17.705 119.595 17.705 119.115 17.375 119.115 17.375 119.595 16.865 119.595 16.865 119.115 16.535 119.115 16.535 119.595 16.025 119.595 16.025 119.115 15.695 119.115 15.695 119.595 14.245 119.595 14.245 118.795 13.915 118.795 13.915 119.595 13.405 119.595 13.405 119.115 13.075 119.115 13.075 119.595 12.565 119.595 12.565 119.115 12.235 119.115 12.235 119.595 11.725 119.595 11.725 119.115 11.395 119.115 11.395 119.595 10.885 119.595 10.885 119.115 10.555 119.115 10.555 119.595 10.045 119.595 10.045 119.115 9.715 119.115 9.715 119.595 8.265 119.595 8.265 118.795 7.935 118.795 7.935 119.595 7.425 119.595 7.425 119.115 7.095 119.115 7.095 119.595 6.585 119.595 6.585 119.115 6.255 119.115 6.255 119.595 5.745 119.595 5.745 119.115 5.415 119.115 5.415 119.595 4.905 119.595 4.905 119.115 4.575 119.115 4.575 119.595 4.065 119.595 4.065 119.115 3.735 119.115 3.735 119.595 0 119.595 0 119.765 ;
      RECT 72.68 116.875 73.6 117.045 ;
      RECT 0 116.875 3.68 117.045 ;
      RECT 72.68 114.155 73.6 114.325 ;
      RECT 0 114.155 3.68 114.325 ;
      RECT 73.14 111.435 73.6 111.605 ;
      RECT 0 111.435 3.68 111.605 ;
      RECT 73.14 108.715 73.6 108.885 ;
      RECT 0 108.715 3.68 108.885 ;
      RECT 72.68 105.995 73.6 106.165 ;
      RECT 0 105.995 1.84 106.165 ;
      RECT 72.68 103.275 73.6 103.445 ;
      RECT 0 103.275 1.84 103.445 ;
      RECT 72.68 100.555 73.6 100.725 ;
      RECT 0 100.555 1.84 100.725 ;
      RECT 72.68 97.835 73.6 98.005 ;
      RECT 0 97.835 1.84 98.005 ;
      RECT 72.68 95.115 73.6 95.285 ;
      RECT 0 95.115 3.68 95.285 ;
      RECT 72.68 92.395 73.6 92.565 ;
      RECT 0 92.395 3.68 92.565 ;
      RECT 72.68 89.675 73.6 89.845 ;
      RECT 0 89.675 3.68 89.845 ;
      RECT 72.68 86.955 73.6 87.125 ;
      RECT 0 86.955 3.68 87.125 ;
      RECT 72.68 84.235 73.6 84.405 ;
      RECT 0 84.235 1.84 84.405 ;
      RECT 72.68 81.515 73.6 81.685 ;
      RECT 0 81.515 1.84 81.685 ;
      RECT 72.68 78.795 73.6 78.965 ;
      RECT 0 78.795 1.84 78.965 ;
      RECT 72.68 76.075 73.6 76.245 ;
      RECT 0 76.075 3.68 76.245 ;
      RECT 72.68 73.355 73.6 73.525 ;
      RECT 0 73.355 3.68 73.525 ;
      RECT 72.68 70.635 73.6 70.805 ;
      RECT 0 70.635 1.84 70.805 ;
      RECT 72.68 67.915 73.6 68.085 ;
      RECT 0 67.915 1.84 68.085 ;
      RECT 72.68 65.195 73.6 65.365 ;
      RECT 0 65.195 1.84 65.365 ;
      RECT 72.68 62.475 73.6 62.645 ;
      RECT 0 62.475 1.84 62.645 ;
      RECT 72.68 59.755 73.6 59.925 ;
      RECT 0 59.755 1.84 59.925 ;
      RECT 72.68 57.035 73.6 57.205 ;
      RECT 0 57.035 1.84 57.205 ;
      RECT 72.68 54.315 73.6 54.485 ;
      RECT 0 54.315 3.68 54.485 ;
      RECT 72.68 51.595 73.6 51.765 ;
      RECT 0 51.595 3.68 51.765 ;
      RECT 72.68 48.875 73.6 49.045 ;
      RECT 0 48.875 1.84 49.045 ;
      RECT 72.68 46.155 73.6 46.325 ;
      RECT 0 46.155 1.84 46.325 ;
      RECT 72.68 43.435 73.6 43.605 ;
      RECT 0 43.435 1.84 43.605 ;
      RECT 72.68 40.715 73.6 40.885 ;
      RECT 0 40.715 1.84 40.885 ;
      RECT 72.68 37.995 73.6 38.165 ;
      RECT 0 37.995 1.84 38.165 ;
      RECT 72.68 35.275 73.6 35.445 ;
      RECT 0 35.275 1.84 35.445 ;
      RECT 72.68 32.555 73.6 32.725 ;
      RECT 0 32.555 1.84 32.725 ;
      RECT 72.68 29.835 73.6 30.005 ;
      RECT 0 29.835 1.84 30.005 ;
      RECT 69.92 27.115 73.6 27.285 ;
      RECT 0 27.115 1.84 27.285 ;
      RECT 69.92 24.395 73.6 24.565 ;
      RECT 0 24.395 1.84 24.565 ;
      RECT 72.68 21.675 73.6 21.845 ;
      RECT 0 21.675 1.84 21.845 ;
      RECT 72.68 18.955 73.6 19.125 ;
      RECT 0 18.955 1.84 19.125 ;
      RECT 72.68 16.235 73.6 16.405 ;
      RECT 0 16.235 1.84 16.405 ;
      RECT 72.68 13.515 73.6 13.685 ;
      RECT 0 13.515 1.84 13.685 ;
      RECT 72.68 10.795 73.6 10.965 ;
      RECT 0 10.795 1.84 10.965 ;
      RECT 72.68 8.075 73.6 8.245 ;
      RECT 0 8.075 1.84 8.245 ;
      RECT 72.68 5.355 73.6 5.525 ;
      RECT 0 5.355 1.84 5.525 ;
      RECT 72.68 2.635 73.6 2.805 ;
      RECT 0 2.635 3.68 2.805 ;
      POLYGON 46.14 0.905 46.14 0.085 47.395 0.085 47.395 0.885 47.725 0.885 47.725 0.085 48.235 0.085 48.235 0.565 48.565 0.565 48.565 0.085 49.075 0.085 49.075 0.565 49.405 0.565 49.405 0.085 49.915 0.085 49.915 0.565 50.245 0.565 50.245 0.085 50.755 0.085 50.755 0.565 51.085 0.565 51.085 0.085 51.595 0.085 51.595 0.565 51.925 0.565 51.925 0.085 52.915 0.085 52.915 0.885 53.245 0.885 53.245 0.085 53.755 0.085 53.755 0.565 54.085 0.565 54.085 0.085 54.595 0.085 54.595 0.565 54.925 0.565 54.925 0.085 55.435 0.085 55.435 0.565 55.765 0.565 55.765 0.085 56.275 0.085 56.275 0.565 56.605 0.565 56.605 0.085 57.115 0.085 57.115 0.565 57.445 0.565 57.445 0.085 58.935 0.085 58.935 0.595 59.35 0.595 59.35 0.085 60.765 0.085 60.765 0.485 61.095 0.485 61.095 0.085 61.605 0.085 61.605 0.485 61.935 0.485 61.935 0.085 67.325 0.085 67.325 0.485 67.655 0.485 67.655 0.085 68.165 0.085 68.165 0.485 68.495 0.485 68.495 0.085 69.91 0.085 69.91 0.595 70.325 0.595 70.325 0.085 73.6 0.085 73.6 -0.085 0 -0.085 0 0.085 4.235 0.085 4.235 0.885 4.565 0.885 4.565 0.085 5.075 0.085 5.075 0.565 5.405 0.565 5.405 0.085 5.915 0.085 5.915 0.565 6.245 0.565 6.245 0.085 6.835 0.085 6.835 0.565 7.005 0.565 7.005 0.085 7.675 0.085 7.675 0.565 7.845 0.565 7.845 0.085 8.935 0.085 8.935 0.545 9.205 0.545 9.205 0.085 10.995 0.085 10.995 0.545 11.32 0.545 11.32 0.085 12.395 0.085 12.395 0.565 12.565 0.565 12.565 0.085 13.235 0.085 13.235 0.565 13.405 0.565 13.405 0.085 13.995 0.085 13.995 0.565 14.325 0.565 14.325 0.085 14.835 0.085 14.835 0.565 15.165 0.565 15.165 0.085 15.675 0.085 15.675 0.885 16.005 0.885 16.005 0.085 17.075 0.085 17.075 0.565 17.405 0.565 17.405 0.085 17.915 0.085 17.915 0.565 18.245 0.565 18.245 0.085 18.755 0.085 18.755 0.565 19.085 0.565 19.085 0.085 19.595 0.085 19.595 0.565 19.925 0.565 19.925 0.085 20.435 0.085 20.435 0.565 20.765 0.565 20.765 0.085 21.275 0.085 21.275 0.885 21.605 0.885 21.605 0.085 22.595 0.085 22.595 0.565 22.925 0.565 22.925 0.085 23.435 0.085 23.435 0.565 23.765 0.565 23.765 0.085 24.275 0.085 24.275 0.565 24.605 0.565 24.605 0.085 25.115 0.085 25.115 0.565 25.445 0.565 25.445 0.085 25.955 0.085 25.955 0.565 26.285 0.565 26.285 0.085 26.795 0.085 26.795 0.885 27.125 0.885 27.125 0.085 29.035 0.085 29.035 0.565 29.365 0.565 29.365 0.085 29.875 0.085 29.875 0.565 30.205 0.565 30.205 0.085 30.715 0.085 30.715 0.565 31.045 0.565 31.045 0.085 31.555 0.085 31.555 0.565 31.885 0.565 31.885 0.085 32.395 0.085 32.395 0.565 32.725 0.565 32.725 0.085 33.235 0.085 33.235 0.885 33.565 0.885 33.565 0.085 35.475 0.085 35.475 0.565 35.805 0.565 35.805 0.085 36.315 0.085 36.315 0.565 36.645 0.565 36.645 0.085 37.155 0.085 37.155 0.565 37.485 0.565 37.485 0.085 37.995 0.085 37.995 0.565 38.325 0.565 38.325 0.085 38.835 0.085 38.835 0.565 39.165 0.565 39.165 0.085 39.675 0.085 39.675 0.885 40.005 0.885 40.005 0.085 41.195 0.085 41.195 0.545 41.45 0.545 41.45 0.085 42.12 0.085 42.12 0.545 42.29 0.545 42.29 0.085 42.96 0.085 42.96 0.545 43.13 0.545 43.13 0.085 43.8 0.085 43.8 0.545 43.97 0.545 43.97 0.085 44.64 0.085 44.64 0.545 44.945 0.545 44.945 0.085 45.91 0.085 45.91 0.905 ;
      RECT 0.17 0.17 73.43 119.51 ;
    LAYER met3 ;
      POLYGON 59.045 119.725 59.045 119.72 59.26 119.72 59.26 119.4 59.045 119.4 59.045 119.395 58.715 119.395 58.715 119.4 58.5 119.4 58.5 119.72 58.715 119.72 58.715 119.725 ;
      POLYGON 29.605 119.725 29.605 119.72 29.82 119.72 29.82 119.4 29.605 119.4 29.605 119.395 29.275 119.395 29.275 119.4 29.06 119.4 29.06 119.72 29.275 119.72 29.275 119.725 ;
      POLYGON 34.895 119.505 34.895 119.49 36.15 119.49 36.15 119.5 36.53 119.5 36.53 119.18 36.15 119.18 36.15 119.19 34.895 119.19 34.895 119.175 34.565 119.175 34.565 119.505 ;
      POLYGON 21.095 119.505 21.095 119.49 26.03 119.49 26.03 119.5 26.41 119.5 26.41 119.18 26.03 119.18 26.03 119.19 21.095 119.19 21.095 119.175 20.765 119.175 20.765 119.505 ;
      POLYGON 31.01 119.5 31.01 119.18 30.97 119.18 30.97 117.83 30.67 117.83 30.67 119.18 30.63 119.18 30.63 119.5 ;
      POLYGON 7.05 1.85 7.05 0.5 7.09 0.5 7.09 0.18 6.71 0.18 6.71 0.5 6.75 0.5 6.75 1.85 ;
      POLYGON 59.045 0.285 59.045 0.28 59.26 0.28 59.26 -0.04 59.045 -0.04 59.045 -0.045 58.715 -0.045 58.715 -0.04 58.5 -0.04 58.5 0.28 58.715 0.28 58.715 0.285 ;
      POLYGON 29.605 0.285 29.605 0.28 29.82 0.28 29.82 -0.04 29.605 -0.04 29.605 -0.045 29.275 -0.045 29.275 -0.04 29.06 -0.04 29.06 0.28 29.275 0.28 29.275 0.285 ;
      RECT 0.4 0.4 73.2 119.28 ;
    LAYER via ;
      RECT 58.805 119.485 58.955 119.635 ;
      RECT 29.365 119.485 29.515 119.635 ;
      RECT 55.355 119.095 55.505 119.245 ;
      RECT 8.435 0.435 8.585 0.585 ;
      RECT 58.805 0.045 58.955 0.195 ;
      RECT 29.365 0.045 29.515 0.195 ;
    LAYER via2 ;
      RECT 58.78 119.46 58.98 119.66 ;
      RECT 29.34 119.46 29.54 119.66 ;
      RECT 34.63 119.24 34.83 119.44 ;
      RECT 20.83 119.24 21.03 119.44 ;
      RECT 58.78 0.02 58.98 0.22 ;
      RECT 29.34 0.02 29.54 0.22 ;
    LAYER via3 ;
      RECT 58.78 119.46 58.98 119.66 ;
      RECT 29.34 119.46 29.54 119.66 ;
      RECT 36.24 119.24 36.44 119.44 ;
      RECT 30.72 119.24 30.92 119.44 ;
      RECT 26.12 119.24 26.32 119.44 ;
      RECT 38.08 0.92 38.28 1.12 ;
      RECT 6.8 0.24 7 0.44 ;
      RECT 58.78 0.02 58.98 0.22 ;
      RECT 29.34 0.02 29.54 0.22 ;
    LAYER OVERLAP ;
      POLYGON 0 0 0 119.68 73.6 119.68 73.6 0 ;
  END
END cby_2__1_

END LIBRARY
