VERSION 5.7 ;
BUSBITCHARS "[]" ;

UNITS
  DATABASE MICRONS 1000 ;
END UNITS

MANUFACTURINGGRID 0.005 ;

LAYER li1
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.46 ;
  WIDTH 0.17 ;
END li1

LAYER mcon
  TYPE CUT ;
END mcon

LAYER met1
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.34 ;
  WIDTH 0.14 ;
END met1

LAYER via
  TYPE CUT ;
END via

LAYER met2
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.46 ;
  WIDTH 0.14 ;
END met2

LAYER via2
  TYPE CUT ;
END via2

LAYER met3
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.68 ;
  WIDTH 0.3 ;
END met3

LAYER via3
  TYPE CUT ;
END via3

LAYER met4
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.92 ;
  WIDTH 0.3 ;
END met4

LAYER via4
  TYPE CUT ;
END via4

LAYER met5
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 3.4 ;
  WIDTH 1.6 ;
END met5

LAYER nwell
  TYPE MASTERSLICE ;
END nwell

LAYER pwell
  TYPE MASTERSLICE ;
END pwell

LAYER OVERLAP
  TYPE OVERLAP ;
END OVERLAP

VIA L1M1_PR
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.145 -0.115 0.145 0.115 ;
END L1M1_PR

VIA L1M1_PR_R
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.115 -0.145 0.115 0.145 ;
END L1M1_PR_R

VIA L1M1_PR_M
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.115 -0.145 0.115 0.145 ;
END L1M1_PR_M

VIA L1M1_PR_MR
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.145 -0.115 0.145 0.115 ;
END L1M1_PR_MR

VIA L1M1_PR_C
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.145 -0.145 0.145 0.145 ;
END L1M1_PR_C

VIA M1M2_PR
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR

VIA M1M2_PR_Enc
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_Enc

VIA M1M2_PR_R
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_R

VIA M1M2_PR_R_Enc
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR_R_Enc

VIA M1M2_PR_M
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_M

VIA M1M2_PR_M_Enc
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR_M_Enc

VIA M1M2_PR_MR
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR_MR

VIA M1M2_PR_MR_Enc
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_MR_Enc

VIA M1M2_PR_C
  LAYER met1 ;
    RECT -0.16 -0.16 0.16 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.16 0.16 0.16 ;
END M1M2_PR_C

VIA M2M3_PR
  LAYER met2 ;
    RECT -0.14 -0.185 0.14 0.185 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR

VIA M2M3_PR_R
  LAYER met2 ;
    RECT -0.185 -0.14 0.185 0.14 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_R

VIA M2M3_PR_M
  LAYER met2 ;
    RECT -0.14 -0.185 0.14 0.185 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_M

VIA M2M3_PR_MR
  LAYER met2 ;
    RECT -0.185 -0.14 0.185 0.14 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_MR

VIA M2M3_PR_C
  LAYER met2 ;
    RECT -0.185 -0.185 0.185 0.185 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_C

VIA M3M4_PR
  LAYER met3 ;
    RECT -0.19 -0.16 0.19 0.16 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR

VIA M3M4_PR_R
  LAYER met3 ;
    RECT -0.16 -0.19 0.16 0.19 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_R

VIA M3M4_PR_M
  LAYER met3 ;
    RECT -0.19 -0.16 0.19 0.16 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_M

VIA M3M4_PR_MR
  LAYER met3 ;
    RECT -0.16 -0.19 0.16 0.19 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_MR

VIA M3M4_PR_C
  LAYER met3 ;
    RECT -0.19 -0.19 0.19 0.19 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_C

VIA M4M5_PR
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR

VIA M4M5_PR_R
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_R

VIA M4M5_PR_M
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_M

VIA M4M5_PR_MR
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_MR

VIA M4M5_PR_C
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_C

SITE unit
  CLASS CORE ;
  SYMMETRY Y ;
  SIZE 0.46 BY 2.72 ;
END unit

SITE unithddbl
  CLASS CORE ;
  SIZE 0.46 BY 5.44 ;
END unithddbl

MACRO cby_1__1_
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  SIZE 73.6 BY 119.68 ;
  SYMMETRY X Y ;
  PIN pReset[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 64.02 0.595 64.16 ;
    END
  END pReset[0]
  PIN chany_bottom_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.16 0 46.3 0.485 ;
    END
  END chany_bottom_in[0]
  PIN chany_bottom_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.88 0 15.02 0.485 ;
    END
  END chany_bottom_in[1]
  PIN chany_bottom_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.74 0 10.88 0.485 ;
    END
  END chany_bottom_in[2]
  PIN chany_bottom_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.92 0 49.06 0.485 ;
    END
  END chany_bottom_in[3]
  PIN chany_bottom_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.64 0 17.78 0.485 ;
    END
  END chany_bottom_in[4]
  PIN chany_bottom_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.44 0 31.58 0.485 ;
    END
  END chany_bottom_in[5]
  PIN chany_bottom_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.24 0 45.38 0.485 ;
    END
  END chany_bottom_in[6]
  PIN chany_bottom_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.32 0 44.46 0.485 ;
    END
  END chany_bottom_in[7]
  PIN chany_bottom_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.28 0 33.42 0.485 ;
    END
  END chany_bottom_in[8]
  PIN chany_bottom_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.8 0 38.94 0.485 ;
    END
  END chany_bottom_in[9]
  PIN chany_bottom_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.88 0 38.02 0.485 ;
    END
  END chany_bottom_in[10]
  PIN chany_bottom_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.04 0 36.18 0.485 ;
    END
  END chany_bottom_in[11]
  PIN chany_bottom_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.36 0 32.5 0.485 ;
    END
  END chany_bottom_in[12]
  PIN chany_bottom_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.48 0 19.62 0.485 ;
    END
  END chany_bottom_in[13]
  PIN chany_bottom_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.52 0 30.66 0.485 ;
    END
  END chany_bottom_in[14]
  PIN chany_bottom_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.72 0 39.86 0.485 ;
    END
  END chany_bottom_in[15]
  PIN chany_bottom_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.8 0 15.94 0.485 ;
    END
  END chany_bottom_in[16]
  PIN chany_bottom_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.2 0 34.34 0.485 ;
    END
  END chany_bottom_in[17]
  PIN chany_bottom_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.56 0 41.7 0.485 ;
    END
  END chany_bottom_in[18]
  PIN chany_bottom_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.56 0 18.7 0.485 ;
    END
  END chany_bottom_in[19]
  PIN chany_bottom_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 61.95 0 62.25 0.8 ;
    END
  END chany_bottom_in[20]
  PIN chany_bottom_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.08 0 47.22 0.485 ;
    END
  END chany_bottom_in[21]
  PIN chany_bottom_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.72 0 16.86 0.485 ;
    END
  END chany_bottom_in[22]
  PIN chany_bottom_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.06 0 7.2 0.485 ;
    END
  END chany_bottom_in[23]
  PIN chany_bottom_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.56 0 64.7 0.485 ;
    END
  END chany_bottom_in[24]
  PIN chany_bottom_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.96 0 14.1 0.485 ;
    END
  END chany_bottom_in[25]
  PIN chany_bottom_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.12 0 35.26 0.485 ;
    END
  END chany_bottom_in[26]
  PIN chany_bottom_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.44 0 8.58 0.485 ;
    END
  END chany_bottom_in[27]
  PIN chany_bottom_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.96 0 37.1 0.485 ;
    END
  END chany_bottom_in[28]
  PIN chany_bottom_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.04 0 13.18 0.485 ;
    END
  END chany_bottom_in[29]
  PIN chany_top_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.82 119.195 55.96 119.68 ;
    END
  END chany_top_in[0]
  PIN chany_top_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.96 119.195 14.1 119.68 ;
    END
  END chany_top_in[1]
  PIN chany_top_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.12 119.195 12.26 119.68 ;
    END
  END chany_top_in[2]
  PIN chany_top_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.18 119.195 63.32 119.68 ;
    END
  END chany_top_in[3]
  PIN chany_top_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.76 119.195 50.9 119.68 ;
    END
  END chany_top_in[4]
  PIN chany_top_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.8 119.195 15.94 119.68 ;
    END
  END chany_top_in[5]
  PIN chany_top_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.1 119.195 41.24 119.68 ;
    END
  END chany_top_in[6]
  PIN chany_top_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.64 119.195 17.78 119.68 ;
    END
  END chany_top_in[7]
  PIN chany_top_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.72 119.195 16.86 119.68 ;
    END
  END chany_top_in[8]
  PIN chany_top_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.96 119.195 37.1 119.68 ;
    END
  END chany_top_in[9]
  PIN chany_top_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.04 119.195 36.18 119.68 ;
    END
  END chany_top_in[10]
  PIN chany_top_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.34 119.195 61.48 119.68 ;
    END
  END chany_top_in[11]
  PIN chany_top_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.66 119.195 57.8 119.68 ;
    END
  END chany_top_in[12]
  PIN chany_top_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.92 119.195 49.06 119.68 ;
    END
  END chany_top_in[13]
  PIN chany_top_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.2 119.195 34.34 119.68 ;
    END
  END chany_top_in[14]
  PIN chany_top_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.34 119.195 38.48 119.68 ;
    END
  END chany_top_in[15]
  PIN chany_top_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.18 119.195 40.32 119.68 ;
    END
  END chany_top_in[16]
  PIN chany_top_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.12 119.195 35.26 119.68 ;
    END
  END chany_top_in[17]
  PIN chany_top_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48 119.195 48.14 119.68 ;
    END
  END chany_top_in[18]
  PIN chany_top_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.08 119.195 47.22 119.68 ;
    END
  END chany_top_in[19]
  PIN chany_top_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.5 119.195 59.64 119.68 ;
    END
  END chany_top_in[20]
  PIN chany_top_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.44 119.195 31.58 119.68 ;
    END
  END chany_top_in[21]
  PIN chany_top_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.04 119.195 13.18 119.68 ;
    END
  END chany_top_in[22]
  PIN chany_top_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.52 119.195 30.66 119.68 ;
    END
  END chany_top_in[23]
  PIN chany_top_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.74 119.195 56.88 119.68 ;
    END
  END chany_top_in[24]
  PIN chany_top_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.36 119.195 32.5 119.68 ;
    END
  END chany_top_in[25]
  PIN chany_top_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.28 119.195 33.42 119.68 ;
    END
  END chany_top_in[26]
  PIN chany_top_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.56 119.195 18.7 119.68 ;
    END
  END chany_top_in[27]
  PIN chany_top_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.26 119.195 39.4 119.68 ;
    END
  END chany_top_in[28]
  PIN chany_top_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.88 119.195 15.02 119.68 ;
    END
  END chany_top_in[29]
  PIN ccff_head[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 17.44 0.595 17.58 ;
    END
  END ccff_head[0]
  PIN chany_bottom_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 45.39 0 45.69 0.8 ;
    END
  END chany_bottom_out[0]
  PIN chany_bottom_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 49.07 0 49.37 0.8 ;
    END
  END chany_bottom_out[1]
  PIN chany_bottom_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.74 0 56.88 0.485 ;
    END
  END chany_bottom_out[2]
  PIN chany_bottom_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 56.43 0 56.73 0.8 ;
    END
  END chany_bottom_out[3]
  PIN chany_bottom_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 33.43 0 33.73 0.8 ;
    END
  END chany_bottom_out[4]
  PIN chany_bottom_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.64 0 40.78 0.485 ;
    END
  END chany_bottom_out[5]
  PIN chany_bottom_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.26 0 62.4 0.485 ;
    END
  END chany_bottom_out[6]
  PIN chany_bottom_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 47.23 0 47.53 0.8 ;
    END
  END chany_bottom_out[7]
  PIN chany_bottom_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 39.87 0 40.17 0.8 ;
    END
  END chany_bottom_out[8]
  PIN chany_bottom_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.3 0 4.44 0.485 ;
    END
  END chany_bottom_out[9]
  PIN chany_bottom_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.22 0 5.36 0.485 ;
    END
  END chany_bottom_out[10]
  PIN chany_bottom_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.48 0 65.62 0.485 ;
    END
  END chany_bottom_out[11]
  PIN chany_bottom_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.22 0 51.36 0.485 ;
    END
  END chany_bottom_out[12]
  PIN chany_bottom_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48 0 48.14 0.485 ;
    END
  END chany_bottom_out[13]
  PIN chany_bottom_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 31.59 0 31.89 0.8 ;
    END
  END chany_bottom_out[14]
  PIN chany_bottom_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 41.71 0 42.01 0.8 ;
    END
  END chany_bottom_out[15]
  PIN chany_bottom_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.82 0 55.96 0.485 ;
    END
  END chany_bottom_out[16]
  PIN chany_bottom_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.64 0 63.78 0.485 ;
    END
  END chany_bottom_out[17]
  PIN chany_bottom_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 52.75 0 53.05 0.8 ;
    END
  END chany_bottom_out[18]
  PIN chany_bottom_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.84 0 49.98 0.485 ;
    END
  END chany_bottom_out[19]
  PIN chany_bottom_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.66 0 11.8 0.485 ;
    END
  END chany_bottom_out[20]
  PIN chany_bottom_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 35.27 0 35.57 0.8 ;
    END
  END chany_bottom_out[21]
  PIN chany_bottom_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 38.03 0 38.33 0.8 ;
    END
  END chany_bottom_out[22]
  PIN chany_bottom_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.06 0 53.2 0.485 ;
    END
  END chany_bottom_out[23]
  PIN chany_bottom_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 50.91 0 51.21 0.8 ;
    END
  END chany_bottom_out[24]
  PIN chany_bottom_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 54.59 0 54.89 0.8 ;
    END
  END chany_bottom_out[25]
  PIN chany_bottom_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.66 0 57.8 0.485 ;
    END
  END chany_bottom_out[26]
  PIN chany_bottom_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.5 0 59.64 0.485 ;
    END
  END chany_bottom_out[27]
  PIN chany_bottom_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.34 0 61.48 0.485 ;
    END
  END chany_bottom_out[28]
  PIN chany_bottom_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.14 0 52.28 0.485 ;
    END
  END chany_bottom_out[29]
  PIN chany_top_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 39.87 118.88 40.17 119.68 ;
    END
  END chany_top_out[0]
  PIN chany_top_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 60.11 118.88 60.41 119.68 ;
    END
  END chany_top_out[1]
  PIN chany_top_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 36.19 118.88 36.49 119.68 ;
    END
  END chany_top_out[2]
  PIN chany_top_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 61.95 118.88 62.25 119.68 ;
    END
  END chany_top_out[3]
  PIN chany_top_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 56.43 118.88 56.73 119.68 ;
    END
  END chany_top_out[4]
  PIN chany_top_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 32.51 118.88 32.81 119.68 ;
    END
  END chany_top_out[5]
  PIN chany_top_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 53.67 118.88 53.97 119.68 ;
    END
  END chany_top_out[6]
  PIN chany_top_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.36 119.195 9.5 119.68 ;
    END
  END chany_top_out[7]
  PIN chany_top_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.26 119.195 62.4 119.68 ;
    END
  END chany_top_out[8]
  PIN chany_top_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.24 119.195 45.38 119.68 ;
    END
  END chany_top_out[9]
  PIN chany_top_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 45.39 118.88 45.69 119.68 ;
    END
  END chany_top_out[10]
  PIN chany_top_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 41.71 118.88 42.01 119.68 ;
    END
  END chany_top_out[11]
  PIN chany_top_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 65.63 118.88 65.93 119.68 ;
    END
  END chany_top_out[12]
  PIN chany_top_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.86 119.195 67 119.68 ;
    END
  END chany_top_out[13]
  PIN chany_top_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.1 119.195 64.24 119.68 ;
    END
  END chany_top_out[14]
  PIN chany_top_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.16 119.195 46.3 119.68 ;
    END
  END chany_top_out[15]
  PIN chany_top_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 34.35 118.88 34.65 119.68 ;
    END
  END chany_top_out[16]
  PIN chany_top_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 30.67 118.88 30.97 119.68 ;
    END
  END chany_top_out[17]
  PIN chany_top_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 63.79 118.88 64.09 119.68 ;
    END
  END chany_top_out[18]
  PIN chany_top_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 50.91 118.88 51.21 119.68 ;
    END
  END chany_top_out[19]
  PIN chany_top_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.94 119.195 66.08 119.68 ;
    END
  END chany_top_out[20]
  PIN chany_top_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.02 119.195 65.16 119.68 ;
    END
  END chany_top_out[21]
  PIN chany_top_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.28 119.195 10.42 119.68 ;
    END
  END chany_top_out[22]
  PIN chany_top_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.32 119.195 44.46 119.68 ;
    END
  END chany_top_out[23]
  PIN chany_top_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 67.47 118.88 67.77 119.68 ;
    END
  END chany_top_out[24]
  PIN chany_top_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.84 119.195 49.98 119.68 ;
    END
  END chany_top_out[25]
  PIN chany_top_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 38.03 118.88 38.33 119.68 ;
    END
  END chany_top_out[26]
  PIN chany_top_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.42 119.195 60.56 119.68 ;
    END
  END chany_top_out[27]
  PIN chany_top_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 47.23 118.88 47.53 119.68 ;
    END
  END chany_top_out[28]
  PIN chany_top_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 49.07 118.88 49.37 119.68 ;
    END
  END chany_top_out[29]
  PIN left_grid_pin_16_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 63.34 0.595 63.48 ;
    END
  END left_grid_pin_16_[0]
  PIN left_grid_pin_17_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 105.16 0.595 105.3 ;
    END
  END left_grid_pin_17_[0]
  PIN left_grid_pin_18_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 83.4 0.595 83.54 ;
    END
  END left_grid_pin_18_[0]
  PIN left_grid_pin_19_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 85.1 0.595 85.24 ;
    END
  END left_grid_pin_19_[0]
  PIN left_grid_pin_20_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 41.58 0.595 41.72 ;
    END
  END left_grid_pin_20_[0]
  PIN left_grid_pin_21_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 39.88 0.595 40.02 ;
    END
  END left_grid_pin_21_[0]
  PIN left_grid_pin_22_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 42.26 0.595 42.4 ;
    END
  END left_grid_pin_22_[0]
  PIN left_grid_pin_23_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 61.64 0.595 61.78 ;
    END
  END left_grid_pin_23_[0]
  PIN left_grid_pin_24_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 37.16 0.595 37.3 ;
    END
  END left_grid_pin_24_[0]
  PIN left_grid_pin_25_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 60.96 0.595 61.1 ;
    END
  END left_grid_pin_25_[0]
  PIN left_grid_pin_26_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 19.82 0.595 19.96 ;
    END
  END left_grid_pin_26_[0]
  PIN left_grid_pin_27_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 39.2 0.595 39.34 ;
    END
  END left_grid_pin_27_[0]
  PIN left_grid_pin_28_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 4.52 0.595 4.66 ;
    END
  END left_grid_pin_28_[0]
  PIN left_grid_pin_29_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 3.84 0.595 3.98 ;
    END
  END left_grid_pin_29_[0]
  PIN left_grid_pin_30_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 18.12 0.595 18.26 ;
    END
  END left_grid_pin_30_[0]
  PIN left_grid_pin_31_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 20.5 0.595 20.64 ;
    END
  END left_grid_pin_31_[0]
  PIN ccff_tail[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 73.005 105.16 73.6 105.3 ;
    END
  END ccff_tail[0]
  PIN Test_en_S_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.98 0 54.12 0.485 ;
    END
  END Test_en_S_in
  PIN Test_en_E_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 73.005 77.62 73.6 77.76 ;
    END
  END Test_en_E_in
  PIN Test_en_W_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 80.68 0.595 80.82 ;
    END
  END Test_en_W_in
  PIN Test_en_N_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.14 119.195 52.28 119.68 ;
    END
  END Test_en_N_out
  PIN Test_en_W_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 69.8 0.595 69.94 ;
    END
  END Test_en_W_out
  PIN Test_en_E_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 73.005 71.5 73.6 71.64 ;
    END
  END Test_en_E_out
  PIN pReset_S_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.36 0 9.5 0.485 ;
    END
  END pReset_S_in
  PIN pReset_N_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.2 119.195 11.34 119.68 ;
    END
  END pReset_N_out
  PIN Reset_S_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.9 0 55.04 0.485 ;
    END
  END Reset_S_in
  PIN Reset_E_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 73.005 68.78 73.6 68.92 ;
    END
  END Reset_E_in
  PIN Reset_W_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 77.96 0.595 78.1 ;
    END
  END Reset_W_in
  PIN Reset_N_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.06 119.195 53.2 119.68 ;
    END
  END Reset_N_out
  PIN Reset_W_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 71.5 0.595 71.64 ;
    END
  END Reset_W_out
  PIN Reset_E_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 73.005 63.68 73.6 63.82 ;
    END
  END Reset_E_out
  PIN prog_clk_0_W_in
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER met1 ;
        RECT 0 1.8 0.595 1.94 ;
    END
  END prog_clk_0_W_in
  PIN prog_clk_0_S_out
    DIRECTION OUTPUT ;
    USE CLOCK ;
    PORT
      LAYER met2 ;
        RECT 6.14 0 6.28 0.485 ;
    END
  END prog_clk_0_S_out
  PIN prog_clk_0_N_out
    DIRECTION OUTPUT ;
    USE CLOCK ;
    PORT
      LAYER met2 ;
        RECT 6.14 119.195 6.28 119.68 ;
    END
  END prog_clk_0_N_out
  PIN prog_clk_2_N_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.78 119.195 67.92 119.68 ;
    END
  END prog_clk_2_N_in
  PIN prog_clk_2_S_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.86 0 67 0.485 ;
    END
  END prog_clk_2_S_in
  PIN prog_clk_2_S_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.4 0 43.54 0.485 ;
    END
  END prog_clk_2_S_out
  PIN prog_clk_2_N_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.4 119.195 43.54 119.68 ;
    END
  END prog_clk_2_N_out
  PIN prog_clk_3_S_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.78 0 67.92 0.485 ;
    END
  END prog_clk_3_S_in
  PIN prog_clk_3_N_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.7 119.195 68.84 119.68 ;
    END
  END prog_clk_3_N_in
  PIN prog_clk_3_N_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.98 119.195 54.12 119.68 ;
    END
  END prog_clk_3_N_out
  PIN prog_clk_3_S_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.7 0 68.84 0.485 ;
    END
  END prog_clk_3_S_out
  PIN clk_2_N_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.62 119.195 69.76 119.68 ;
    END
  END clk_2_N_in
  PIN clk_2_S_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.62 0 69.76 0.485 ;
    END
  END clk_2_S_in
  PIN clk_2_S_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.48 0 42.62 0.485 ;
    END
  END clk_2_S_out
  PIN clk_2_N_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.48 119.195 42.62 119.68 ;
    END
  END clk_2_N_out
  PIN clk_3_S_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71 0 71.14 0.485 ;
    END
  END clk_3_S_in
  PIN clk_3_N_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71 119.195 71.14 119.68 ;
    END
  END clk_3_N_in
  PIN clk_3_N_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.9 119.195 55.04 119.68 ;
    END
  END clk_3_N_out
  PIN clk_3_S_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.42 0 60.56 0.485 ;
    END
  END clk_3_S_out
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0 7.24 3.2 10.44 ;
        RECT 70.4 7.24 73.6 10.44 ;
        RECT 0 48.04 3.2 51.24 ;
        RECT 70.4 48.04 73.6 51.24 ;
        RECT 0 88.84 3.2 92.04 ;
        RECT 70.4 88.84 73.6 92.04 ;
      LAYER met4 ;
        RECT 14.42 0 15.02 0.6 ;
        RECT 43.86 0 44.46 0.6 ;
        RECT 14.42 119.08 15.02 119.68 ;
        RECT 43.86 119.08 44.46 119.68 ;
      LAYER met1 ;
        RECT 0 2.48 0.48 2.96 ;
        RECT 73.12 2.48 73.6 2.96 ;
        RECT 0 7.92 0.48 8.4 ;
        RECT 73.12 7.92 73.6 8.4 ;
        RECT 0 13.36 0.48 13.84 ;
        RECT 73.12 13.36 73.6 13.84 ;
        RECT 0 18.8 0.48 19.28 ;
        RECT 73.12 18.8 73.6 19.28 ;
        RECT 0 24.24 0.48 24.72 ;
        RECT 73.12 24.24 73.6 24.72 ;
        RECT 0 29.68 0.48 30.16 ;
        RECT 73.12 29.68 73.6 30.16 ;
        RECT 0 35.12 0.48 35.6 ;
        RECT 73.12 35.12 73.6 35.6 ;
        RECT 0 40.56 0.48 41.04 ;
        RECT 73.12 40.56 73.6 41.04 ;
        RECT 0 46 0.48 46.48 ;
        RECT 73.12 46 73.6 46.48 ;
        RECT 0 51.44 0.48 51.92 ;
        RECT 73.12 51.44 73.6 51.92 ;
        RECT 0 56.88 0.48 57.36 ;
        RECT 73.12 56.88 73.6 57.36 ;
        RECT 0 62.32 0.48 62.8 ;
        RECT 73.12 62.32 73.6 62.8 ;
        RECT 0 67.76 0.48 68.24 ;
        RECT 73.12 67.76 73.6 68.24 ;
        RECT 0 73.2 0.48 73.68 ;
        RECT 73.12 73.2 73.6 73.68 ;
        RECT 0 78.64 0.48 79.12 ;
        RECT 73.12 78.64 73.6 79.12 ;
        RECT 0 84.08 0.48 84.56 ;
        RECT 73.12 84.08 73.6 84.56 ;
        RECT 0 89.52 0.48 90 ;
        RECT 73.12 89.52 73.6 90 ;
        RECT 0 94.96 0.48 95.44 ;
        RECT 73.12 94.96 73.6 95.44 ;
        RECT 0 100.4 0.48 100.88 ;
        RECT 73.12 100.4 73.6 100.88 ;
        RECT 0 105.84 0.48 106.32 ;
        RECT 73.12 105.84 73.6 106.32 ;
        RECT 0 111.28 0.48 111.76 ;
        RECT 73.12 111.28 73.6 111.76 ;
        RECT 0 116.72 0.48 117.2 ;
        RECT 73.12 116.72 73.6 117.2 ;
    END
  END VDD
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0 27.64 3.2 30.84 ;
        RECT 70.4 27.64 73.6 30.84 ;
        RECT 0 68.44 3.2 71.64 ;
        RECT 70.4 68.44 73.6 71.64 ;
        RECT 0 109.24 3.2 112.44 ;
        RECT 70.4 109.24 73.6 112.44 ;
      LAYER met4 ;
        RECT 29.14 0 29.74 0.6 ;
        RECT 58.58 0 59.18 0.6 ;
        RECT 29.14 119.08 29.74 119.68 ;
        RECT 58.58 119.08 59.18 119.68 ;
      LAYER met1 ;
        RECT 0 -0.24 0.48 0.24 ;
        RECT 73.12 -0.24 73.6 0.24 ;
        RECT 0 5.2 0.48 5.68 ;
        RECT 73.12 5.2 73.6 5.68 ;
        RECT 0 10.64 0.48 11.12 ;
        RECT 73.12 10.64 73.6 11.12 ;
        RECT 0 16.08 0.48 16.56 ;
        RECT 73.12 16.08 73.6 16.56 ;
        RECT 0 21.52 0.48 22 ;
        RECT 73.12 21.52 73.6 22 ;
        RECT 0 26.96 0.48 27.44 ;
        RECT 73.12 26.96 73.6 27.44 ;
        RECT 0 32.4 0.48 32.88 ;
        RECT 73.12 32.4 73.6 32.88 ;
        RECT 0 37.84 0.48 38.32 ;
        RECT 73.12 37.84 73.6 38.32 ;
        RECT 0 43.28 0.48 43.76 ;
        RECT 73.12 43.28 73.6 43.76 ;
        RECT 0 48.72 0.48 49.2 ;
        RECT 73.12 48.72 73.6 49.2 ;
        RECT 0 54.16 0.48 54.64 ;
        RECT 73.12 54.16 73.6 54.64 ;
        RECT 0 59.6 0.48 60.08 ;
        RECT 73.12 59.6 73.6 60.08 ;
        RECT 0 65.04 0.48 65.52 ;
        RECT 73.12 65.04 73.6 65.52 ;
        RECT 0 70.48 0.48 70.96 ;
        RECT 73.12 70.48 73.6 70.96 ;
        RECT 0 75.92 0.48 76.4 ;
        RECT 73.12 75.92 73.6 76.4 ;
        RECT 0 81.36 0.48 81.84 ;
        RECT 73.12 81.36 73.6 81.84 ;
        RECT 0 86.8 0.48 87.28 ;
        RECT 73.12 86.8 73.6 87.28 ;
        RECT 0 92.24 0.48 92.72 ;
        RECT 73.12 92.24 73.6 92.72 ;
        RECT 0 97.68 0.48 98.16 ;
        RECT 73.12 97.68 73.6 98.16 ;
        RECT 0 103.12 0.48 103.6 ;
        RECT 73.12 103.12 73.6 103.6 ;
        RECT 0 108.56 0.48 109.04 ;
        RECT 73.12 108.56 73.6 109.04 ;
        RECT 0 114 0.48 114.48 ;
        RECT 73.12 114 73.6 114.48 ;
        RECT 0 119.44 0.48 119.92 ;
        RECT 73.12 119.44 73.6 119.92 ;
    END
  END VSS
  OBS
    LAYER met1 ;
      POLYGON 72.84 119.92 72.84 119.44 59.04 119.44 59.04 119.43 58.72 119.43 58.72 119.44 29.6 119.44 29.6 119.43 29.28 119.43 29.28 119.44 0.76 119.44 0.76 119.92 ;
      POLYGON 59.04 0.25 59.04 0.24 72.84 0.24 72.84 -0.24 0.76 -0.24 0.76 0.24 29.28 0.24 29.28 0.25 29.6 0.25 29.6 0.24 58.72 0.24 58.72 0.25 ;
      POLYGON 72.84 119.4 72.84 119.16 73.32 119.16 73.32 117.48 72.84 117.48 72.84 116.44 73.32 116.44 73.32 114.76 72.84 114.76 72.84 113.72 73.32 113.72 73.32 112.04 72.84 112.04 72.84 111 73.32 111 73.32 109.32 72.84 109.32 72.84 108.28 73.32 108.28 73.32 106.6 72.84 106.6 72.84 105.58 72.725 105.58 72.725 104.88 73.32 104.88 73.32 103.88 72.84 103.88 72.84 102.84 73.32 102.84 73.32 101.16 72.84 101.16 72.84 100.12 73.32 100.12 73.32 98.44 72.84 98.44 72.84 97.4 73.32 97.4 73.32 95.72 72.84 95.72 72.84 94.68 73.32 94.68 73.32 93 72.84 93 72.84 91.96 73.32 91.96 73.32 90.28 72.84 90.28 72.84 89.24 73.32 89.24 73.32 87.56 72.84 87.56 72.84 86.52 73.32 86.52 73.32 84.84 72.84 84.84 72.84 83.8 73.32 83.8 73.32 82.12 72.84 82.12 72.84 81.08 73.32 81.08 73.32 79.4 72.84 79.4 72.84 78.36 73.32 78.36 73.32 78.04 72.725 78.04 72.725 77.34 73.32 77.34 73.32 76.68 72.84 76.68 72.84 75.64 73.32 75.64 73.32 73.96 72.84 73.96 72.84 72.92 73.32 72.92 73.32 71.92 72.725 71.92 72.725 71.22 72.84 71.22 72.84 70.2 73.32 70.2 73.32 69.2 72.725 69.2 72.725 68.5 72.84 68.5 72.84 67.48 73.32 67.48 73.32 65.8 72.84 65.8 72.84 64.76 73.32 64.76 73.32 64.1 72.725 64.1 72.725 63.4 73.32 63.4 73.32 63.08 72.84 63.08 72.84 62.04 73.32 62.04 73.32 60.36 72.84 60.36 72.84 59.32 73.32 59.32 73.32 57.64 72.84 57.64 72.84 56.6 73.32 56.6 73.32 54.92 72.84 54.92 72.84 53.88 73.32 53.88 73.32 52.2 72.84 52.2 72.84 51.16 73.32 51.16 73.32 49.48 72.84 49.48 72.84 48.44 73.32 48.44 73.32 46.76 72.84 46.76 72.84 45.72 73.32 45.72 73.32 44.04 72.84 44.04 72.84 43 73.32 43 73.32 41.32 72.84 41.32 72.84 40.28 73.32 40.28 73.32 38.6 72.84 38.6 72.84 37.56 73.32 37.56 73.32 35.88 72.84 35.88 72.84 34.84 73.32 34.84 73.32 33.16 72.84 33.16 72.84 32.12 73.32 32.12 73.32 30.44 72.84 30.44 72.84 29.4 73.32 29.4 73.32 27.72 72.84 27.72 72.84 26.68 73.32 26.68 73.32 25 72.84 25 72.84 23.96 73.32 23.96 73.32 22.28 72.84 22.28 72.84 21.24 73.32 21.24 73.32 19.56 72.84 19.56 72.84 18.52 73.32 18.52 73.32 16.84 72.84 16.84 72.84 15.8 73.32 15.8 73.32 14.12 72.84 14.12 72.84 13.08 73.32 13.08 73.32 11.4 72.84 11.4 72.84 10.36 73.32 10.36 73.32 8.68 72.84 8.68 72.84 7.64 73.32 7.64 73.32 5.96 72.84 5.96 72.84 4.92 73.32 4.92 73.32 3.24 72.84 3.24 72.84 2.2 73.32 2.2 73.32 0.52 72.84 0.52 72.84 0.28 0.76 0.28 0.76 0.52 0.28 0.52 0.28 1.52 0.875 1.52 0.875 2.22 0.76 2.22 0.76 3.24 0.28 3.24 0.28 3.56 0.875 3.56 0.875 4.94 0.76 4.94 0.76 5.96 0.28 5.96 0.28 7.64 0.76 7.64 0.76 8.68 0.28 8.68 0.28 10.36 0.76 10.36 0.76 11.4 0.28 11.4 0.28 13.08 0.76 13.08 0.76 14.12 0.28 14.12 0.28 15.8 0.76 15.8 0.76 16.84 0.28 16.84 0.28 17.16 0.875 17.16 0.875 18.54 0.76 18.54 0.76 19.54 0.875 19.54 0.875 20.92 0.28 20.92 0.28 21.24 0.76 21.24 0.76 22.28 0.28 22.28 0.28 23.96 0.76 23.96 0.76 25 0.28 25 0.28 26.68 0.76 26.68 0.76 27.72 0.28 27.72 0.28 29.4 0.76 29.4 0.76 30.44 0.28 30.44 0.28 32.12 0.76 32.12 0.76 33.16 0.28 33.16 0.28 34.84 0.76 34.84 0.76 35.88 0.28 35.88 0.28 36.88 0.875 36.88 0.875 37.58 0.76 37.58 0.76 38.6 0.28 38.6 0.28 38.92 0.875 38.92 0.875 40.3 0.76 40.3 0.76 41.3 0.875 41.3 0.875 42.68 0.28 42.68 0.28 43 0.76 43 0.76 44.04 0.28 44.04 0.28 45.72 0.76 45.72 0.76 46.76 0.28 46.76 0.28 48.44 0.76 48.44 0.76 49.48 0.28 49.48 0.28 51.16 0.76 51.16 0.76 52.2 0.28 52.2 0.28 53.88 0.76 53.88 0.76 54.92 0.28 54.92 0.28 56.6 0.76 56.6 0.76 57.64 0.28 57.64 0.28 59.32 0.76 59.32 0.76 60.36 0.28 60.36 0.28 60.68 0.875 60.68 0.875 62.06 0.76 62.06 0.76 63.06 0.875 63.06 0.875 64.44 0.28 64.44 0.28 64.76 0.76 64.76 0.76 65.8 0.28 65.8 0.28 67.48 0.76 67.48 0.76 68.52 0.28 68.52 0.28 69.52 0.875 69.52 0.875 70.22 0.76 70.22 0.76 71.22 0.875 71.22 0.875 71.92 0.28 71.92 0.28 72.92 0.76 72.92 0.76 73.96 0.28 73.96 0.28 75.64 0.76 75.64 0.76 76.68 0.28 76.68 0.28 77.68 0.875 77.68 0.875 78.38 0.76 78.38 0.76 79.4 0.28 79.4 0.28 80.4 0.875 80.4 0.875 81.1 0.76 81.1 0.76 82.12 0.28 82.12 0.28 83.12 0.875 83.12 0.875 83.82 0.76 83.82 0.76 84.82 0.875 84.82 0.875 85.52 0.28 85.52 0.28 86.52 0.76 86.52 0.76 87.56 0.28 87.56 0.28 89.24 0.76 89.24 0.76 90.28 0.28 90.28 0.28 91.96 0.76 91.96 0.76 93 0.28 93 0.28 94.68 0.76 94.68 0.76 95.72 0.28 95.72 0.28 97.4 0.76 97.4 0.76 98.44 0.28 98.44 0.28 100.12 0.76 100.12 0.76 101.16 0.28 101.16 0.28 102.84 0.76 102.84 0.76 103.88 0.28 103.88 0.28 104.88 0.875 104.88 0.875 105.58 0.76 105.58 0.76 106.6 0.28 106.6 0.28 108.28 0.76 108.28 0.76 109.32 0.28 109.32 0.28 111 0.76 111 0.76 112.04 0.28 112.04 0.28 113.72 0.76 113.72 0.76 114.76 0.28 114.76 0.28 116.44 0.76 116.44 0.76 117.48 0.28 117.48 0.28 119.16 0.76 119.16 0.76 119.4 ;
    LAYER met2 ;
      RECT 58.74 119.375 59.02 119.745 ;
      RECT 29.3 119.375 29.58 119.745 ;
      POLYGON 50.48 119.58 50.48 119.44 50.44 119.44 50.44 112.98 50.3 112.98 50.3 119.58 ;
      POLYGON 31.12 119.58 31.12 112.98 30.98 112.98 30.98 119.44 30.94 119.44 30.94 119.58 ;
      RECT 39.66 119.01 39.92 119.33 ;
      POLYGON 9.96 12.48 9.96 0.1 9.78 0.1 9.78 0.24 9.82 0.24 9.82 12.48 ;
      POLYGON 3.06 11.97 3.06 0.24 4.02 0.24 4.02 0.1 2.92 0.1 2.92 11.97 ;
      POLYGON 44.92 7.04 44.92 0.1 44.74 0.1 44.74 0.24 44.78 0.24 44.78 7.04 ;
      POLYGON 15.48 4.32 15.48 0.1 15.3 0.1 15.3 0.24 15.34 0.24 15.34 4.32 ;
      POLYGON 11.34 1.26 11.34 0.525 11.41 0.525 11.41 0.155 11.13 0.155 11.13 0.525 11.2 0.525 11.2 1.26 ;
      RECT 58.74 -0.065 59.02 0.305 ;
      RECT 29.3 -0.065 29.58 0.305 ;
      POLYGON 73.32 119.4 73.32 0.28 71.42 0.28 71.42 0.765 70.72 0.765 70.72 0.28 70.04 0.28 70.04 0.765 69.34 0.765 69.34 0.28 69.12 0.28 69.12 0.765 68.42 0.765 68.42 0.28 68.2 0.28 68.2 0.765 67.5 0.765 67.5 0.28 67.28 0.28 67.28 0.765 66.58 0.765 66.58 0.28 65.9 0.28 65.9 0.765 65.2 0.765 65.2 0.28 64.98 0.28 64.98 0.765 64.28 0.765 64.28 0.28 64.06 0.28 64.06 0.765 63.36 0.765 63.36 0.28 62.68 0.28 62.68 0.765 61.98 0.765 61.98 0.28 61.76 0.28 61.76 0.765 61.06 0.765 61.06 0.28 60.84 0.28 60.84 0.765 60.14 0.765 60.14 0.28 59.92 0.28 59.92 0.765 59.22 0.765 59.22 0.28 58.08 0.28 58.08 0.765 57.38 0.765 57.38 0.28 57.16 0.28 57.16 0.765 56.46 0.765 56.46 0.28 56.24 0.28 56.24 0.765 55.54 0.765 55.54 0.28 55.32 0.28 55.32 0.765 54.62 0.765 54.62 0.28 54.4 0.28 54.4 0.765 53.7 0.765 53.7 0.28 53.48 0.28 53.48 0.765 52.78 0.765 52.78 0.28 52.56 0.28 52.56 0.765 51.86 0.765 51.86 0.28 51.64 0.28 51.64 0.765 50.94 0.765 50.94 0.28 50.26 0.28 50.26 0.765 49.56 0.765 49.56 0.28 49.34 0.28 49.34 0.765 48.64 0.765 48.64 0.28 48.42 0.28 48.42 0.765 47.72 0.765 47.72 0.28 47.5 0.28 47.5 0.765 46.8 0.765 46.8 0.28 46.58 0.28 46.58 0.765 45.88 0.765 45.88 0.28 45.66 0.28 45.66 0.765 44.96 0.765 44.96 0.28 44.74 0.28 44.74 0.765 44.04 0.765 44.04 0.28 43.82 0.28 43.82 0.765 43.12 0.765 43.12 0.28 42.9 0.28 42.9 0.765 42.2 0.765 42.2 0.28 41.98 0.28 41.98 0.765 41.28 0.765 41.28 0.28 41.06 0.28 41.06 0.765 40.36 0.765 40.36 0.28 40.14 0.28 40.14 0.765 39.44 0.765 39.44 0.28 39.22 0.28 39.22 0.765 38.52 0.765 38.52 0.28 38.3 0.28 38.3 0.765 37.6 0.765 37.6 0.28 37.38 0.28 37.38 0.765 36.68 0.765 36.68 0.28 36.46 0.28 36.46 0.765 35.76 0.765 35.76 0.28 35.54 0.28 35.54 0.765 34.84 0.765 34.84 0.28 34.62 0.28 34.62 0.765 33.92 0.765 33.92 0.28 33.7 0.28 33.7 0.765 33 0.765 33 0.28 32.78 0.28 32.78 0.765 32.08 0.765 32.08 0.28 31.86 0.28 31.86 0.765 31.16 0.765 31.16 0.28 30.94 0.28 30.94 0.765 30.24 0.765 30.24 0.28 19.9 0.28 19.9 0.765 19.2 0.765 19.2 0.28 18.98 0.28 18.98 0.765 18.28 0.765 18.28 0.28 18.06 0.28 18.06 0.765 17.36 0.765 17.36 0.28 17.14 0.28 17.14 0.765 16.44 0.765 16.44 0.28 16.22 0.28 16.22 0.765 15.52 0.765 15.52 0.28 15.3 0.28 15.3 0.765 14.6 0.765 14.6 0.28 14.38 0.28 14.38 0.765 13.68 0.765 13.68 0.28 13.46 0.28 13.46 0.765 12.76 0.765 12.76 0.28 12.08 0.28 12.08 0.765 11.38 0.765 11.38 0.28 11.16 0.28 11.16 0.765 10.46 0.765 10.46 0.28 9.78 0.28 9.78 0.765 9.08 0.765 9.08 0.28 8.86 0.28 8.86 0.765 8.16 0.765 8.16 0.28 7.48 0.28 7.48 0.765 6.78 0.765 6.78 0.28 6.56 0.28 6.56 0.765 5.86 0.765 5.86 0.28 5.64 0.28 5.64 0.765 4.94 0.765 4.94 0.28 4.72 0.28 4.72 0.765 4.02 0.765 4.02 0.28 0.28 0.28 0.28 119.4 5.86 119.4 5.86 118.915 6.56 118.915 6.56 119.4 9.08 119.4 9.08 118.915 9.78 118.915 9.78 119.4 10 119.4 10 118.915 10.7 118.915 10.7 119.4 10.92 119.4 10.92 118.915 11.62 118.915 11.62 119.4 11.84 119.4 11.84 118.915 12.54 118.915 12.54 119.4 12.76 119.4 12.76 118.915 13.46 118.915 13.46 119.4 13.68 119.4 13.68 118.915 14.38 118.915 14.38 119.4 14.6 119.4 14.6 118.915 15.3 118.915 15.3 119.4 15.52 119.4 15.52 118.915 16.22 118.915 16.22 119.4 16.44 119.4 16.44 118.915 17.14 118.915 17.14 119.4 17.36 119.4 17.36 118.915 18.06 118.915 18.06 119.4 18.28 119.4 18.28 118.915 18.98 118.915 18.98 119.4 30.24 119.4 30.24 118.915 30.94 118.915 30.94 119.4 31.16 119.4 31.16 118.915 31.86 118.915 31.86 119.4 32.08 119.4 32.08 118.915 32.78 118.915 32.78 119.4 33 119.4 33 118.915 33.7 118.915 33.7 119.4 33.92 119.4 33.92 118.915 34.62 118.915 34.62 119.4 34.84 119.4 34.84 118.915 35.54 118.915 35.54 119.4 35.76 119.4 35.76 118.915 36.46 118.915 36.46 119.4 36.68 119.4 36.68 118.915 37.38 118.915 37.38 119.4 38.06 119.4 38.06 118.915 38.76 118.915 38.76 119.4 38.98 119.4 38.98 118.915 39.68 118.915 39.68 119.4 39.9 119.4 39.9 118.915 40.6 118.915 40.6 119.4 40.82 119.4 40.82 118.915 41.52 118.915 41.52 119.4 42.2 119.4 42.2 118.915 42.9 118.915 42.9 119.4 43.12 119.4 43.12 118.915 43.82 118.915 43.82 119.4 44.04 119.4 44.04 118.915 44.74 118.915 44.74 119.4 44.96 119.4 44.96 118.915 45.66 118.915 45.66 119.4 45.88 119.4 45.88 118.915 46.58 118.915 46.58 119.4 46.8 119.4 46.8 118.915 47.5 118.915 47.5 119.4 47.72 119.4 47.72 118.915 48.42 118.915 48.42 119.4 48.64 119.4 48.64 118.915 49.34 118.915 49.34 119.4 49.56 119.4 49.56 118.915 50.26 118.915 50.26 119.4 50.48 119.4 50.48 118.915 51.18 118.915 51.18 119.4 51.86 119.4 51.86 118.915 52.56 118.915 52.56 119.4 52.78 119.4 52.78 118.915 53.48 118.915 53.48 119.4 53.7 119.4 53.7 118.915 54.4 118.915 54.4 119.4 54.62 119.4 54.62 118.915 55.32 118.915 55.32 119.4 55.54 119.4 55.54 118.915 56.24 118.915 56.24 119.4 56.46 119.4 56.46 118.915 57.16 118.915 57.16 119.4 57.38 119.4 57.38 118.915 58.08 118.915 58.08 119.4 59.22 119.4 59.22 118.915 59.92 118.915 59.92 119.4 60.14 119.4 60.14 118.915 60.84 118.915 60.84 119.4 61.06 119.4 61.06 118.915 61.76 118.915 61.76 119.4 61.98 119.4 61.98 118.915 62.68 118.915 62.68 119.4 62.9 119.4 62.9 118.915 63.6 118.915 63.6 119.4 63.82 119.4 63.82 118.915 64.52 118.915 64.52 119.4 64.74 119.4 64.74 118.915 65.44 118.915 65.44 119.4 65.66 119.4 65.66 118.915 66.36 118.915 66.36 119.4 66.58 119.4 66.58 118.915 67.28 118.915 67.28 119.4 67.5 119.4 67.5 118.915 68.2 118.915 68.2 119.4 68.42 119.4 68.42 118.915 69.12 118.915 69.12 119.4 69.34 119.4 69.34 118.915 70.04 118.915 70.04 119.4 70.72 119.4 70.72 118.915 71.42 118.915 71.42 119.4 ;
    LAYER met4 ;
      POLYGON 53.27 119.49 53.27 119.19 53.05 119.19 53.05 58.67 52.75 58.67 52.75 119.49 ;
      POLYGON 48.45 119.49 48.45 102.87 48.15 102.87 48.15 119.19 47.93 119.19 47.93 119.49 ;
      POLYGON 5.21 14.77 5.21 0.505 5.225 0.505 5.225 0.175 4.895 0.175 4.895 0.505 4.91 0.505 4.91 14.77 ;
      POLYGON 73.2 119.28 73.2 0.4 62.65 0.4 62.65 1.2 61.55 1.2 61.55 0.4 59.58 0.4 59.58 1 58.18 1 58.18 0.4 57.13 0.4 57.13 1.2 56.03 1.2 56.03 0.4 55.29 0.4 55.29 1.2 54.19 1.2 54.19 0.4 53.45 0.4 53.45 1.2 52.35 1.2 52.35 0.4 51.61 0.4 51.61 1.2 50.51 1.2 50.51 0.4 49.77 0.4 49.77 1.2 48.67 1.2 48.67 0.4 47.93 0.4 47.93 1.2 46.83 1.2 46.83 0.4 46.09 0.4 46.09 1.2 44.99 1.2 44.99 0.4 44.86 0.4 44.86 1 43.46 1 43.46 0.4 42.41 0.4 42.41 1.2 41.31 1.2 41.31 0.4 40.57 0.4 40.57 1.2 39.47 1.2 39.47 0.4 38.73 0.4 38.73 1.2 37.63 1.2 37.63 0.4 35.97 0.4 35.97 1.2 34.87 1.2 34.87 0.4 34.13 0.4 34.13 1.2 33.03 1.2 33.03 0.4 32.29 0.4 32.29 1.2 31.19 1.2 31.19 0.4 30.14 0.4 30.14 1 28.74 1 28.74 0.4 15.42 0.4 15.42 1 14.02 1 14.02 0.4 0.4 0.4 0.4 119.28 14.02 119.28 14.02 118.68 15.42 118.68 15.42 119.28 28.74 119.28 28.74 118.68 30.14 118.68 30.14 119.28 30.27 119.28 30.27 118.48 31.37 118.48 31.37 119.28 32.11 119.28 32.11 118.48 33.21 118.48 33.21 119.28 33.95 119.28 33.95 118.48 35.05 118.48 35.05 119.28 35.79 119.28 35.79 118.48 36.89 118.48 36.89 119.28 37.63 119.28 37.63 118.48 38.73 118.48 38.73 119.28 39.47 119.28 39.47 118.48 40.57 118.48 40.57 119.28 41.31 119.28 41.31 118.48 42.41 118.48 42.41 119.28 43.46 119.28 43.46 118.68 44.86 118.68 44.86 119.28 44.99 119.28 44.99 118.48 46.09 118.48 46.09 119.28 46.83 119.28 46.83 118.48 47.93 118.48 47.93 119.28 48.67 119.28 48.67 118.48 49.77 118.48 49.77 119.28 50.51 119.28 50.51 118.48 51.61 118.48 51.61 119.28 53.27 119.28 53.27 118.48 54.37 118.48 54.37 119.28 56.03 119.28 56.03 118.48 57.13 118.48 57.13 119.28 58.18 119.28 58.18 118.68 59.58 118.68 59.58 119.28 59.71 119.28 59.71 118.48 60.81 118.48 60.81 119.28 61.55 119.28 61.55 118.48 62.65 118.48 62.65 119.28 63.39 119.28 63.39 118.48 64.49 118.48 64.49 119.28 65.23 119.28 65.23 118.48 66.33 118.48 66.33 119.28 67.07 119.28 67.07 118.48 68.17 118.48 68.17 119.28 ;
    LAYER met5 ;
      POLYGON 72 118.08 72 114.04 68.8 114.04 68.8 107.64 72 107.64 72 93.64 68.8 93.64 68.8 87.24 72 87.24 72 73.24 68.8 73.24 68.8 66.84 72 66.84 72 52.84 68.8 52.84 68.8 46.44 72 46.44 72 32.44 68.8 32.44 68.8 26.04 72 26.04 72 12.04 68.8 12.04 68.8 5.64 72 5.64 72 1.6 1.6 1.6 1.6 5.64 4.8 5.64 4.8 12.04 1.6 12.04 1.6 26.04 4.8 26.04 4.8 32.44 1.6 32.44 1.6 46.44 4.8 46.44 4.8 52.84 1.6 52.84 1.6 66.84 4.8 66.84 4.8 73.24 1.6 73.24 1.6 87.24 4.8 87.24 4.8 93.64 1.6 93.64 1.6 107.64 4.8 107.64 4.8 114.04 1.6 114.04 1.6 118.08 ;
    LAYER li1 ;
      POLYGON 73.6 119.765 73.6 119.595 69.905 119.595 69.905 118.795 69.575 118.795 69.575 119.595 69.065 119.595 69.065 119.115 68.735 119.115 68.735 119.595 68.225 119.595 68.225 119.115 67.895 119.115 67.895 119.595 67.385 119.595 67.385 119.115 67.055 119.115 67.055 119.595 66.545 119.595 66.545 119.115 66.215 119.115 66.215 119.595 65.705 119.595 65.705 119.115 65.375 119.115 65.375 119.595 64.385 119.595 64.385 118.795 64.055 118.795 64.055 119.595 63.545 119.595 63.545 119.115 63.215 119.115 63.215 119.595 62.705 119.595 62.705 119.115 62.375 119.115 62.375 119.595 61.865 119.595 61.865 119.115 61.535 119.115 61.535 119.595 61.025 119.595 61.025 119.115 60.695 119.115 60.695 119.595 60.185 119.595 60.185 119.115 59.855 119.115 59.855 119.595 58.405 119.595 58.405 118.795 58.075 118.795 58.075 119.595 57.565 119.595 57.565 119.115 57.235 119.115 57.235 119.595 56.725 119.595 56.725 119.115 56.395 119.115 56.395 119.595 55.885 119.595 55.885 119.115 55.555 119.115 55.555 119.595 55.045 119.595 55.045 119.115 54.715 119.115 54.715 119.595 54.205 119.595 54.205 119.115 53.875 119.115 53.875 119.595 52.385 119.595 52.385 119.115 52.055 119.115 52.055 119.595 51.545 119.595 51.545 119.115 51.215 119.115 51.215 119.595 50.705 119.595 50.705 119.115 50.375 119.115 50.375 119.595 49.865 119.595 49.865 119.115 49.535 119.115 49.535 119.595 49.025 119.595 49.025 119.115 48.695 119.115 48.695 119.595 48.185 119.595 48.185 118.795 47.855 118.795 47.855 119.595 46.485 119.595 46.485 119.115 46.315 119.115 46.315 119.595 45.645 119.595 45.645 119.115 45.475 119.115 45.475 119.595 44.885 119.595 44.885 119.115 44.555 119.115 44.555 119.595 44.045 119.595 44.045 119.115 43.715 119.115 43.715 119.595 43.205 119.595 43.205 118.795 42.875 118.795 42.875 119.595 41.845 119.595 41.845 118.795 41.515 118.795 41.515 119.595 41.005 119.595 41.005 119.115 40.675 119.115 40.675 119.595 40.165 119.595 40.165 119.115 39.835 119.115 39.835 119.595 39.325 119.595 39.325 119.115 38.995 119.115 38.995 119.595 38.485 119.595 38.485 119.115 38.155 119.115 38.155 119.595 37.645 119.595 37.645 119.115 37.315 119.115 37.315 119.595 35.865 119.595 35.865 118.795 35.535 118.795 35.535 119.595 35.025 119.595 35.025 119.115 34.695 119.115 34.695 119.595 34.185 119.595 34.185 119.115 33.855 119.115 33.855 119.595 33.345 119.595 33.345 119.115 33.015 119.115 33.015 119.595 32.505 119.595 32.505 119.115 32.175 119.115 32.175 119.595 31.665 119.595 31.665 119.115 31.335 119.115 31.335 119.595 29.885 119.595 29.885 118.795 29.555 118.795 29.555 119.595 29.045 119.595 29.045 119.115 28.715 119.115 28.715 119.595 28.205 119.595 28.205 119.115 27.875 119.115 27.875 119.595 27.365 119.595 27.365 119.115 27.035 119.115 27.035 119.595 26.525 119.595 26.525 119.115 26.195 119.115 26.195 119.595 25.685 119.595 25.685 119.115 25.355 119.115 25.355 119.595 23.905 119.595 23.905 118.795 23.575 118.795 23.575 119.595 23.065 119.595 23.065 119.115 22.735 119.115 22.735 119.595 22.225 119.595 22.225 119.115 21.895 119.115 21.895 119.595 21.385 119.595 21.385 119.115 21.055 119.115 21.055 119.595 20.545 119.595 20.545 119.115 20.215 119.115 20.215 119.595 19.705 119.595 19.705 119.115 19.375 119.115 19.375 119.595 17.925 119.595 17.925 118.795 17.595 118.795 17.595 119.595 17.085 119.595 17.085 119.115 16.755 119.115 16.755 119.595 16.245 119.595 16.245 119.115 15.915 119.115 15.915 119.595 15.405 119.595 15.405 119.115 15.075 119.115 15.075 119.595 14.565 119.595 14.565 119.115 14.235 119.115 14.235 119.595 13.725 119.595 13.725 119.115 13.395 119.115 13.395 119.595 11.905 119.595 11.905 119.115 11.575 119.115 11.575 119.595 11.065 119.595 11.065 119.115 10.735 119.115 10.735 119.595 10.225 119.595 10.225 119.115 9.895 119.115 9.895 119.595 9.385 119.595 9.385 119.115 9.055 119.115 9.055 119.595 8.545 119.595 8.545 119.115 8.215 119.115 8.215 119.595 7.705 119.595 7.705 118.795 7.375 118.795 7.375 119.595 4.995 119.595 4.995 119.215 4.665 119.215 4.665 119.595 0 119.595 0 119.765 ;
      RECT 69.92 116.875 73.6 117.045 ;
      RECT 0 116.875 3.68 117.045 ;
      RECT 69.92 114.155 73.6 114.325 ;
      RECT 0 114.155 1.84 114.325 ;
      RECT 72.68 111.435 73.6 111.605 ;
      RECT 0 111.435 1.84 111.605 ;
      RECT 72.68 108.715 73.6 108.885 ;
      RECT 0 108.715 1.84 108.885 ;
      RECT 72.68 105.995 73.6 106.165 ;
      RECT 0 105.995 1.84 106.165 ;
      RECT 72.68 103.275 73.6 103.445 ;
      RECT 0 103.275 1.84 103.445 ;
      RECT 72.68 100.555 73.6 100.725 ;
      RECT 0 100.555 3.68 100.725 ;
      RECT 72.68 97.835 73.6 98.005 ;
      RECT 0 97.835 3.68 98.005 ;
      RECT 72.68 95.115 73.6 95.285 ;
      RECT 0 95.115 1.84 95.285 ;
      RECT 72.68 92.395 73.6 92.565 ;
      RECT 0 92.395 1.84 92.565 ;
      RECT 72.68 89.675 73.6 89.845 ;
      RECT 0 89.675 1.84 89.845 ;
      RECT 72.68 86.955 73.6 87.125 ;
      RECT 0 86.955 1.84 87.125 ;
      RECT 72.68 84.235 73.6 84.405 ;
      RECT 0 84.235 1.84 84.405 ;
      RECT 72.68 81.515 73.6 81.685 ;
      RECT 0 81.515 1.84 81.685 ;
      RECT 72.68 78.795 73.6 78.965 ;
      RECT 0 78.795 1.84 78.965 ;
      RECT 72.68 76.075 73.6 76.245 ;
      RECT 0 76.075 1.84 76.245 ;
      RECT 72.68 73.355 73.6 73.525 ;
      RECT 0 73.355 1.84 73.525 ;
      RECT 72.68 70.635 73.6 70.805 ;
      RECT 0 70.635 1.84 70.805 ;
      RECT 72.68 67.915 73.6 68.085 ;
      RECT 0 67.915 1.84 68.085 ;
      RECT 72.68 65.195 73.6 65.365 ;
      RECT 0 65.195 1.84 65.365 ;
      RECT 72.68 62.475 73.6 62.645 ;
      RECT 0 62.475 3.68 62.645 ;
      RECT 72.68 59.755 73.6 59.925 ;
      RECT 0 59.755 3.68 59.925 ;
      RECT 72.68 57.035 73.6 57.205 ;
      RECT 0 57.035 1.84 57.205 ;
      RECT 72.68 54.315 73.6 54.485 ;
      RECT 0 54.315 1.84 54.485 ;
      RECT 72.68 51.595 73.6 51.765 ;
      RECT 0 51.595 3.68 51.765 ;
      RECT 72.68 48.875 73.6 49.045 ;
      RECT 0 48.875 3.68 49.045 ;
      RECT 69.92 46.155 73.6 46.325 ;
      RECT 0 46.155 1.84 46.325 ;
      RECT 69.92 43.435 73.6 43.605 ;
      RECT 0 43.435 1.84 43.605 ;
      RECT 72.68 40.715 73.6 40.885 ;
      RECT 0 40.715 3.68 40.885 ;
      RECT 72.68 37.995 73.6 38.165 ;
      RECT 0 37.995 3.68 38.165 ;
      RECT 72.68 35.275 73.6 35.445 ;
      RECT 0 35.275 1.84 35.445 ;
      RECT 69.92 32.555 73.6 32.725 ;
      RECT 0 32.555 1.84 32.725 ;
      RECT 69.92 29.835 73.6 30.005 ;
      RECT 0 29.835 1.84 30.005 ;
      RECT 72.68 27.115 73.6 27.285 ;
      RECT 0 27.115 1.84 27.285 ;
      RECT 72.68 24.395 73.6 24.565 ;
      RECT 0 24.395 1.84 24.565 ;
      RECT 72.68 21.675 73.6 21.845 ;
      RECT 0 21.675 1.84 21.845 ;
      RECT 72.68 18.955 73.6 19.125 ;
      RECT 0 18.955 1.84 19.125 ;
      RECT 72.68 16.235 73.6 16.405 ;
      RECT 0 16.235 3.68 16.405 ;
      RECT 72.68 13.515 73.6 13.685 ;
      RECT 0 13.515 3.68 13.685 ;
      RECT 72.68 10.795 73.6 10.965 ;
      RECT 0 10.795 1.84 10.965 ;
      RECT 72.68 8.075 73.6 8.245 ;
      RECT 0 8.075 3.68 8.245 ;
      RECT 72.68 5.355 73.6 5.525 ;
      RECT 0 5.355 3.68 5.525 ;
      RECT 72.68 2.635 73.6 2.805 ;
      RECT 0 2.635 3.68 2.805 ;
      POLYGON 70.665 0.905 70.665 0.085 73.6 0.085 73.6 -0.085 0 -0.085 0 0.085 4.665 0.085 4.665 0.465 4.995 0.465 4.995 0.085 5.995 0.085 5.995 0.885 6.325 0.885 6.325 0.085 6.835 0.085 6.835 0.565 7.165 0.565 7.165 0.085 7.675 0.085 7.675 0.565 8.005 0.565 8.005 0.085 8.515 0.085 8.515 0.565 8.845 0.565 8.845 0.085 9.355 0.085 9.355 0.565 9.685 0.565 9.685 0.085 10.195 0.085 10.195 0.565 10.525 0.565 10.525 0.085 11.555 0.085 11.555 0.565 11.885 0.565 11.885 0.085 12.395 0.085 12.395 0.565 12.725 0.565 12.725 0.085 13.235 0.085 13.235 0.565 13.565 0.565 13.565 0.085 14.075 0.085 14.075 0.565 14.405 0.565 14.405 0.085 14.915 0.085 14.915 0.565 15.245 0.565 15.245 0.085 15.755 0.085 15.755 0.885 16.085 0.885 16.085 0.085 17.075 0.085 17.075 0.565 17.405 0.565 17.405 0.085 17.915 0.085 17.915 0.565 18.245 0.565 18.245 0.085 18.755 0.085 18.755 0.565 19.085 0.565 19.085 0.085 19.595 0.085 19.595 0.565 19.925 0.565 19.925 0.085 20.435 0.085 20.435 0.565 20.765 0.565 20.765 0.085 21.275 0.085 21.275 0.885 21.605 0.885 21.605 0.085 22.595 0.085 22.595 0.565 22.925 0.565 22.925 0.085 23.435 0.085 23.435 0.565 23.765 0.565 23.765 0.085 24.275 0.085 24.275 0.565 24.605 0.565 24.605 0.085 25.115 0.085 25.115 0.565 25.445 0.565 25.445 0.085 25.955 0.085 25.955 0.565 26.285 0.565 26.285 0.085 26.795 0.085 26.795 0.885 27.125 0.885 27.125 0.085 28.075 0.085 28.075 0.885 28.405 0.885 28.405 0.085 28.915 0.085 28.915 0.565 29.245 0.565 29.245 0.085 29.755 0.085 29.755 0.565 30.085 0.565 30.085 0.085 30.595 0.085 30.595 0.565 30.925 0.565 30.925 0.085 31.435 0.085 31.435 0.565 31.765 0.565 31.765 0.085 32.275 0.085 32.275 0.565 32.605 0.565 32.605 0.085 33.595 0.085 33.595 0.885 33.925 0.885 33.925 0.085 34.435 0.085 34.435 0.565 34.765 0.565 34.765 0.085 35.275 0.085 35.275 0.565 35.605 0.565 35.605 0.085 36.115 0.085 36.115 0.565 36.445 0.565 36.445 0.085 36.955 0.085 36.955 0.565 37.285 0.565 37.285 0.085 37.795 0.085 37.795 0.565 38.125 0.565 38.125 0.085 39.615 0.085 39.615 0.565 39.945 0.565 39.945 0.085 40.455 0.085 40.455 0.565 40.785 0.565 40.785 0.085 41.295 0.085 41.295 0.565 41.625 0.565 41.625 0.085 42.135 0.085 42.135 0.565 42.465 0.565 42.465 0.085 42.975 0.085 42.975 0.565 43.305 0.565 43.305 0.085 43.815 0.085 43.815 0.885 44.145 0.885 44.145 0.085 44.715 0.085 44.715 0.885 45.045 0.885 45.045 0.085 45.555 0.085 45.555 0.565 45.885 0.565 45.885 0.085 46.395 0.085 46.395 0.565 46.725 0.565 46.725 0.085 47.315 0.085 47.315 0.565 47.485 0.565 47.485 0.085 48.155 0.085 48.155 0.565 48.325 0.565 48.325 0.085 50.665 0.085 50.665 0.465 50.995 0.465 50.995 0.085 53.875 0.085 53.875 0.565 54.205 0.565 54.205 0.085 54.715 0.085 54.715 0.565 55.045 0.565 55.045 0.085 55.555 0.085 55.555 0.565 55.885 0.565 55.885 0.085 56.395 0.085 56.395 0.565 56.725 0.565 56.725 0.085 57.235 0.085 57.235 0.565 57.565 0.565 57.565 0.085 58.075 0.085 58.075 0.885 58.405 0.885 58.405 0.085 59.055 0.085 59.055 0.565 59.225 0.565 59.225 0.085 59.895 0.085 59.895 0.565 60.065 0.565 60.065 0.085 60.735 0.085 60.735 0.565 60.905 0.565 60.905 0.085 61.575 0.085 61.575 0.565 61.745 0.565 61.745 0.085 62.415 0.085 62.415 0.565 62.585 0.565 62.585 0.085 63.255 0.085 63.255 0.565 63.425 0.565 63.425 0.085 64.095 0.085 64.095 0.565 64.265 0.565 64.265 0.085 64.935 0.085 64.935 0.565 65.105 0.565 65.105 0.085 65.775 0.085 65.775 0.565 65.945 0.565 65.945 0.085 66.615 0.085 66.615 0.565 66.785 0.565 66.785 0.085 67.455 0.085 67.455 0.565 67.625 0.565 67.625 0.085 68.295 0.085 68.295 0.565 68.465 0.565 68.465 0.085 69.135 0.085 69.135 0.565 69.305 0.565 69.305 0.085 70.495 0.085 70.495 0.905 ;
      RECT 0.17 0.17 73.43 119.51 ;
    LAYER met3 ;
      POLYGON 59.045 119.725 59.045 119.72 59.26 119.72 59.26 119.4 59.045 119.4 59.045 119.395 58.715 119.395 58.715 119.4 58.5 119.4 58.5 119.72 58.715 119.72 58.715 119.725 ;
      POLYGON 29.605 119.725 29.605 119.72 29.82 119.72 29.82 119.4 29.605 119.4 29.605 119.395 29.275 119.395 29.275 119.4 29.06 119.4 29.06 119.72 29.275 119.72 29.275 119.725 ;
      POLYGON 45.69 2.53 45.69 0.5 45.73 0.5 45.73 0.18 45.35 0.18 45.35 0.5 45.39 0.5 45.39 2.53 ;
      POLYGON 11.435 0.505 11.435 0.175 11.105 0.175 11.105 0.19 8.675 0.19 8.675 0.175 8.345 0.175 8.345 0.505 8.675 0.505 8.675 0.49 11.105 0.49 11.105 0.505 ;
      RECT 4.725 0.175 5.455 0.505 ;
      POLYGON 59.045 0.285 59.045 0.28 59.26 0.28 59.26 -0.04 59.045 -0.04 59.045 -0.045 58.715 -0.045 58.715 -0.04 58.5 -0.04 58.5 0.28 58.715 0.28 58.715 0.285 ;
      POLYGON 29.605 0.285 29.605 0.28 29.82 0.28 29.82 -0.04 29.605 -0.04 29.605 -0.045 29.275 -0.045 29.275 -0.04 29.06 -0.04 29.06 0.28 29.275 0.28 29.275 0.285 ;
      RECT 0.4 0.4 73.2 119.28 ;
    LAYER via ;
      RECT 58.805 119.485 58.955 119.635 ;
      RECT 29.365 119.485 29.515 119.635 ;
      RECT 59.495 119.095 59.645 119.245 ;
      RECT 49.835 119.095 49.985 119.245 ;
      RECT 7.055 0.435 7.205 0.585 ;
      RECT 58.805 0.045 58.955 0.195 ;
      RECT 29.365 0.045 29.515 0.195 ;
    LAYER via2 ;
      RECT 58.78 119.46 58.98 119.66 ;
      RECT 29.34 119.46 29.54 119.66 ;
      RECT 11.17 0.24 11.37 0.44 ;
      RECT 8.41 0.24 8.61 0.44 ;
      RECT 5.19 0.24 5.39 0.44 ;
      RECT 58.78 0.02 58.98 0.22 ;
      RECT 29.34 0.02 29.54 0.22 ;
    LAYER via3 ;
      RECT 58.78 119.46 58.98 119.66 ;
      RECT 29.34 119.46 29.54 119.66 ;
      RECT 33.48 0.92 33.68 1.12 ;
      RECT 45.44 0.24 45.64 0.44 ;
      RECT 4.96 0.24 5.16 0.44 ;
      RECT 58.78 0.02 58.98 0.22 ;
      RECT 29.34 0.02 29.54 0.22 ;
    LAYER OVERLAP ;
      POLYGON 0 0 0 119.68 73.6 119.68 73.6 0 ;
  END
END cby_1__1_

END LIBRARY
