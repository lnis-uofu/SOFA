VERSION 5.7 ;
BUSBITCHARS "[]" ;

UNITS
  DATABASE MICRONS 1000 ;
END UNITS

MANUFACTURINGGRID 0.005 ;

LAYER li1
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.46 ;
  WIDTH 0.17 ;
END li1

LAYER mcon
  TYPE CUT ;
END mcon

LAYER met1
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.34 ;
  WIDTH 0.14 ;
END met1

LAYER via
  TYPE CUT ;
END via

LAYER met2
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.46 ;
  WIDTH 0.14 ;
END met2

LAYER via2
  TYPE CUT ;
END via2

LAYER met3
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.68 ;
  WIDTH 0.3 ;
END met3

LAYER via3
  TYPE CUT ;
END via3

LAYER met4
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.92 ;
  WIDTH 0.3 ;
END met4

LAYER via4
  TYPE CUT ;
END via4

LAYER met5
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 3.4 ;
  WIDTH 1.6 ;
END met5

LAYER nwell
  TYPE MASTERSLICE ;
END nwell

LAYER pwell
  TYPE MASTERSLICE ;
END pwell

LAYER OVERLAP
  TYPE OVERLAP ;
END OVERLAP

VIA L1M1_PR
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.145 -0.115 0.145 0.115 ;
END L1M1_PR

VIA L1M1_PR_R
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.115 -0.145 0.115 0.145 ;
END L1M1_PR_R

VIA L1M1_PR_M
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.115 -0.145 0.115 0.145 ;
END L1M1_PR_M

VIA L1M1_PR_MR
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.145 -0.115 0.145 0.115 ;
END L1M1_PR_MR

VIA L1M1_PR_C
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.145 -0.145 0.145 0.145 ;
END L1M1_PR_C

VIA M1M2_PR
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR

VIA M1M2_PR_Enc
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_Enc

VIA M1M2_PR_R
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_R

VIA M1M2_PR_R_Enc
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR_R_Enc

VIA M1M2_PR_M
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_M

VIA M1M2_PR_M_Enc
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR_M_Enc

VIA M1M2_PR_MR
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR_MR

VIA M1M2_PR_MR_Enc
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_MR_Enc

VIA M1M2_PR_C
  LAYER met1 ;
    RECT -0.16 -0.16 0.16 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.16 0.16 0.16 ;
END M1M2_PR_C

VIA M2M3_PR
  LAYER met2 ;
    RECT -0.14 -0.185 0.14 0.185 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR

VIA M2M3_PR_R
  LAYER met2 ;
    RECT -0.185 -0.14 0.185 0.14 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_R

VIA M2M3_PR_M
  LAYER met2 ;
    RECT -0.14 -0.185 0.14 0.185 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_M

VIA M2M3_PR_MR
  LAYER met2 ;
    RECT -0.185 -0.14 0.185 0.14 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_MR

VIA M2M3_PR_C
  LAYER met2 ;
    RECT -0.185 -0.185 0.185 0.185 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_C

VIA M3M4_PR
  LAYER met3 ;
    RECT -0.19 -0.16 0.19 0.16 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR

VIA M3M4_PR_R
  LAYER met3 ;
    RECT -0.16 -0.19 0.16 0.19 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_R

VIA M3M4_PR_M
  LAYER met3 ;
    RECT -0.19 -0.16 0.19 0.16 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_M

VIA M3M4_PR_MR
  LAYER met3 ;
    RECT -0.16 -0.19 0.16 0.19 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_MR

VIA M3M4_PR_C
  LAYER met3 ;
    RECT -0.19 -0.19 0.19 0.19 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_C

VIA M4M5_PR
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR

VIA M4M5_PR_R
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_R

VIA M4M5_PR_M
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_M

VIA M4M5_PR_MR
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_MR

VIA M4M5_PR_C
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_C

SITE unit
  CLASS CORE ;
  SYMMETRY Y ;
  SIZE 0.46 BY 2.72 ;
END unit

SITE unithddbl
  CLASS CORE ;
  SIZE 0.46 BY 5.44 ;
END unithddbl

MACRO cbx_1__0_
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  SIZE 66.24 BY 87.04 ;
  SYMMETRY X Y ;
  PIN prog_clk[0]
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER met3 ;
        RECT 64.86 13.45 66.24 13.75 ;
    END
  END prog_clk[0]
  PIN chanx_left_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 56.97 1.38 57.27 ;
    END
  END chanx_left_in[0]
  PIN chanx_left_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 67.85 1.38 68.15 ;
    END
  END chanx_left_in[1]
  PIN chanx_left_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 43.37 1.38 43.67 ;
    END
  END chanx_left_in[2]
  PIN chanx_left_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 80.09 1.38 80.39 ;
    END
  END chanx_left_in[3]
  PIN chanx_left_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 33.85 1.38 34.15 ;
    END
  END chanx_left_in[4]
  PIN chanx_left_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 82.13 1.38 82.43 ;
    END
  END chanx_left_in[5]
  PIN chanx_left_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 39.29 1.38 39.59 ;
    END
  END chanx_left_in[6]
  PIN chanx_left_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 53.57 1.38 53.87 ;
    END
  END chanx_left_in[7]
  PIN chanx_left_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 47.45 1.38 47.75 ;
    END
  END chanx_left_in[8]
  PIN chanx_left_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 78.73 1.38 79.03 ;
    END
  END chanx_left_in[9]
  PIN chanx_left_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 46.09 1.38 46.39 ;
    END
  END chanx_left_in[10]
  PIN chanx_left_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 69.21 1.38 69.51 ;
    END
  END chanx_left_in[11]
  PIN chanx_left_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 40.65 1.38 40.95 ;
    END
  END chanx_left_in[12]
  PIN chanx_left_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 37.93 1.38 38.23 ;
    END
  END chanx_left_in[13]
  PIN chanx_left_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 29.77 1.38 30.07 ;
    END
  END chanx_left_in[14]
  PIN chanx_left_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 52.21 1.38 52.51 ;
    END
  END chanx_left_in[15]
  PIN chanx_left_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 58.33 1.38 58.63 ;
    END
  END chanx_left_in[16]
  PIN chanx_left_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 63.09 1.38 63.39 ;
    END
  END chanx_left_in[17]
  PIN chanx_left_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 70.57 1.38 70.87 ;
    END
  END chanx_left_in[18]
  PIN chanx_left_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 65.13 1.38 65.43 ;
    END
  END chanx_left_in[19]
  PIN chanx_right_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 64.86 59.69 66.24 59.99 ;
    END
  END chanx_right_in[0]
  PIN chanx_right_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 64.86 56.29 66.24 56.59 ;
    END
  END chanx_right_in[1]
  PIN chanx_right_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 64.86 77.37 66.24 77.67 ;
    END
  END chanx_right_in[2]
  PIN chanx_right_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 64.86 80.09 66.24 80.39 ;
    END
  END chanx_right_in[3]
  PIN chanx_right_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 64.86 48.13 66.24 48.43 ;
    END
  END chanx_right_in[4]
  PIN chanx_right_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 64.86 82.13 66.24 82.43 ;
    END
  END chanx_right_in[5]
  PIN chanx_right_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 64.86 73.29 66.24 73.59 ;
    END
  END chanx_right_in[6]
  PIN chanx_right_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 64.86 58.33 66.24 58.63 ;
    END
  END chanx_right_in[7]
  PIN chanx_right_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 64.86 19.57 66.24 19.87 ;
    END
  END chanx_right_in[8]
  PIN chanx_right_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 64.86 44.73 66.24 45.03 ;
    END
  END chanx_right_in[9]
  PIN chanx_right_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 64.86 71.93 66.24 72.23 ;
    END
  END chanx_right_in[10]
  PIN chanx_right_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 64.86 70.57 66.24 70.87 ;
    END
  END chanx_right_in[11]
  PIN chanx_right_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 64.86 74.65 66.24 74.95 ;
    END
  END chanx_right_in[12]
  PIN chanx_right_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 64.86 65.13 66.24 65.43 ;
    END
  END chanx_right_in[13]
  PIN chanx_right_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 64.86 27.73 66.24 28.03 ;
    END
  END chanx_right_in[14]
  PIN chanx_right_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 64.86 49.49 66.24 49.79 ;
    END
  END chanx_right_in[15]
  PIN chanx_right_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 64.86 40.65 66.24 40.95 ;
    END
  END chanx_right_in[16]
  PIN chanx_right_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 64.86 8.69 66.24 8.99 ;
    END
  END chanx_right_in[17]
  PIN chanx_right_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 64.86 50.85 66.24 51.15 ;
    END
  END chanx_right_in[18]
  PIN chanx_right_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 64.86 52.21 66.24 52.51 ;
    END
  END chanx_right_in[19]
  PIN ccff_head[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 64.86 16.85 66.24 17.15 ;
    END
  END ccff_head[0]
  PIN chanx_left_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 73.29 1.38 73.59 ;
    END
  END chanx_left_out[0]
  PIN chanx_left_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 71.93 1.38 72.23 ;
    END
  END chanx_left_out[1]
  PIN chanx_left_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 9.37 1.38 9.67 ;
    END
  END chanx_left_out[2]
  PIN chanx_left_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 21.61 1.38 21.91 ;
    END
  END chanx_left_out[3]
  PIN chanx_left_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 76.01 1.38 76.31 ;
    END
  END chanx_left_out[4]
  PIN chanx_left_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 22.97 1.38 23.27 ;
    END
  END chanx_left_out[5]
  PIN chanx_left_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 42.01 1.38 42.31 ;
    END
  END chanx_left_out[6]
  PIN chanx_left_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 36.57 1.38 36.87 ;
    END
  END chanx_left_out[7]
  PIN chanx_left_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 24.33 1.38 24.63 ;
    END
  END chanx_left_out[8]
  PIN chanx_left_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 44.73 1.38 45.03 ;
    END
  END chanx_left_out[9]
  PIN chanx_left_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 54.93 1.38 55.23 ;
    END
  END chanx_left_out[10]
  PIN chanx_left_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 31.13 1.38 31.43 ;
    END
  END chanx_left_out[11]
  PIN chanx_left_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 12.09 1.38 12.39 ;
    END
  END chanx_left_out[12]
  PIN chanx_left_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 83.49 1.38 83.79 ;
    END
  END chanx_left_out[13]
  PIN chanx_left_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 77.37 1.38 77.67 ;
    END
  END chanx_left_out[14]
  PIN chanx_left_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 26.37 1.38 26.67 ;
    END
  END chanx_left_out[15]
  PIN chanx_left_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 32.49 1.38 32.79 ;
    END
  END chanx_left_out[16]
  PIN chanx_left_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 10.73 1.38 11.03 ;
    END
  END chanx_left_out[17]
  PIN chanx_left_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 35.21 1.38 35.51 ;
    END
  END chanx_left_out[18]
  PIN chanx_left_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 28.41 1.38 28.71 ;
    END
  END chanx_left_out[19]
  PIN chanx_right_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 64.86 11.41 66.24 11.71 ;
    END
  END chanx_right_out[0]
  PIN chanx_right_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 64.86 66.49 66.24 66.79 ;
    END
  END chanx_right_out[1]
  PIN chanx_right_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 64.86 10.05 66.24 10.35 ;
    END
  END chanx_right_out[2]
  PIN chanx_right_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 64.86 21.61 66.24 21.91 ;
    END
  END chanx_right_out[3]
  PIN chanx_right_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 64.86 78.73 66.24 79.03 ;
    END
  END chanx_right_out[4]
  PIN chanx_right_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 64.86 15.49 66.24 15.79 ;
    END
  END chanx_right_out[5]
  PIN chanx_right_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 64.86 33.17 66.24 33.47 ;
    END
  END chanx_right_out[6]
  PIN chanx_right_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 64.86 83.49 66.24 83.79 ;
    END
  END chanx_right_out[7]
  PIN chanx_right_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 64.86 25.69 66.24 25.99 ;
    END
  END chanx_right_out[8]
  PIN chanx_right_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 64.86 34.53 66.24 34.83 ;
    END
  END chanx_right_out[9]
  PIN chanx_right_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 64.86 39.29 66.24 39.59 ;
    END
  END chanx_right_out[10]
  PIN chanx_right_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 64.86 18.21 66.24 18.51 ;
    END
  END chanx_right_out[11]
  PIN chanx_right_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 64.86 76.01 66.24 76.31 ;
    END
  END chanx_right_out[12]
  PIN chanx_right_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 64.86 69.21 66.24 69.51 ;
    END
  END chanx_right_out[13]
  PIN chanx_right_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 64.86 42.01 66.24 42.31 ;
    END
  END chanx_right_out[14]
  PIN chanx_right_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 64.86 46.09 66.24 46.39 ;
    END
  END chanx_right_out[15]
  PIN chanx_right_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 64.86 29.77 66.24 30.07 ;
    END
  END chanx_right_out[16]
  PIN chanx_right_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 64.86 24.33 66.24 24.63 ;
    END
  END chanx_right_out[17]
  PIN chanx_right_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 64.86 22.97 66.24 23.27 ;
    END
  END chanx_right_out[18]
  PIN chanx_right_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 64.86 67.85 66.24 68.15 ;
    END
  END chanx_right_out[19]
  PIN bottom_grid_pin_0_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 16.17 1.38 16.47 ;
    END
  END bottom_grid_pin_0_[0]
  PIN bottom_grid_pin_2_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.43 85.68 11.57 87.04 ;
    END
  END bottom_grid_pin_2_[0]
  PIN bottom_grid_pin_4_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 18.89 1.38 19.19 ;
    END
  END bottom_grid_pin_4_[0]
  PIN bottom_grid_pin_6_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 64.86 5.97 66.24 6.27 ;
    END
  END bottom_grid_pin_6_[0]
  PIN bottom_grid_pin_8_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.09 0 44.23 1.36 ;
    END
  END bottom_grid_pin_8_[0]
  PIN bottom_grid_pin_10_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.91 0 29.05 1.36 ;
    END
  END bottom_grid_pin_10_[0]
  PIN ccff_tail[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 13.45 1.38 13.75 ;
    END
  END ccff_tail[0]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.49 0 39.63 1.36 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[0]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.63 0 20.77 1.36 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[1]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.87 0 41.01 1.36 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[2]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.51 0 33.65 1.36 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[3]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.61 0 26.75 1.36 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[4]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.11 0 61.25 1.36 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[5]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.43 0 34.57 1.36 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[0]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.07 0 4.21 1.36 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[1]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.19 0 14.33 1.36 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[2]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.25 0 42.39 1.36 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[3]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.05 0 56.19 1.36 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[4]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.85 0 23.99 1.36 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[5]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.21 0 31.35 1.36 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[0]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.99 0 28.13 1.36 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[1]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.77 0 24.91 1.36 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[2]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.81 0 12.95 1.36 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[3]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.67 0 8.81 1.36 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[4]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.75 0 7.89 1.36 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[5]
  PIN top_width_0_height_0__pin_0_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 17.53 1.38 17.83 ;
    END
  END top_width_0_height_0__pin_0_[0]
  PIN top_width_0_height_0__pin_2_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.35 85.68 12.49 87.04 ;
    END
  END top_width_0_height_0__pin_2_[0]
  PIN top_width_0_height_0__pin_4_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 20.25 1.38 20.55 ;
    END
  END top_width_0_height_0__pin_4_[0]
  PIN top_width_0_height_0__pin_6_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 64.86 7.33 66.24 7.63 ;
    END
  END top_width_0_height_0__pin_6_[0]
  PIN top_width_0_height_0__pin_8_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.17 0 43.31 1.36 ;
    END
  END top_width_0_height_0__pin_8_[0]
  PIN top_width_0_height_0__pin_10_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.83 0 29.97 1.36 ;
    END
  END top_width_0_height_0__pin_10_[0]
  PIN top_width_0_height_0__pin_1_upper[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 74.65 1.38 74.95 ;
    END
  END top_width_0_height_0__pin_1_upper[0]
  PIN top_width_0_height_0__pin_1_lower[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 64.86 63.77 66.24 64.07 ;
    END
  END top_width_0_height_0__pin_1_lower[0]
  PIN top_width_0_height_0__pin_3_upper[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 59.69 1.38 59.99 ;
    END
  END top_width_0_height_0__pin_3_upper[0]
  PIN top_width_0_height_0__pin_3_lower[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 64.86 31.13 66.24 31.43 ;
    END
  END top_width_0_height_0__pin_3_lower[0]
  PIN top_width_0_height_0__pin_5_upper[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 66.49 1.38 66.79 ;
    END
  END top_width_0_height_0__pin_5_upper[0]
  PIN top_width_0_height_0__pin_5_lower[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 64.86 43.37 66.24 43.67 ;
    END
  END top_width_0_height_0__pin_5_lower[0]
  PIN top_width_0_height_0__pin_7_upper[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 50.17 1.38 50.47 ;
    END
  END top_width_0_height_0__pin_7_upper[0]
  PIN top_width_0_height_0__pin_7_lower[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 64.86 54.25 66.24 54.55 ;
    END
  END top_width_0_height_0__pin_7_lower[0]
  PIN top_width_0_height_0__pin_9_upper[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 61.73 1.38 62.03 ;
    END
  END top_width_0_height_0__pin_9_upper[0]
  PIN top_width_0_height_0__pin_9_lower[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 64.86 61.73 66.24 62.03 ;
    END
  END top_width_0_height_0__pin_9_lower[0]
  PIN top_width_0_height_0__pin_11_upper[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 48.81 1.38 49.11 ;
    END
  END top_width_0_height_0__pin_11_upper[0]
  PIN top_width_0_height_0__pin_11_lower[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 64.86 37.25 66.24 37.55 ;
    END
  END top_width_0_height_0__pin_11_lower[0]
  PIN SC_IN_TOP
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.87 85.68 64.01 87.04 ;
    END
  END SC_IN_TOP
  PIN SC_IN_BOT
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 14.81 1.38 15.11 ;
    END
  END SC_IN_BOT
  PIN SC_OUT_TOP
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.19 85.68 14.33 87.04 ;
    END
  END SC_OUT_TOP
  PIN SC_OUT_BOT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 64.86 35.89 66.24 36.19 ;
    END
  END SC_OUT_BOT
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0 11.32 3.2 14.52 ;
        RECT 63.04 11.32 66.24 14.52 ;
        RECT 0 52.12 3.2 55.32 ;
        RECT 63.04 52.12 66.24 55.32 ;
      LAYER met4 ;
        RECT 10.74 0 11.34 0.6 ;
        RECT 40.18 0 40.78 0.6 ;
        RECT 10.74 86.44 11.34 87.04 ;
        RECT 40.18 86.44 40.78 87.04 ;
      LAYER met1 ;
        RECT 0 2.48 0.48 2.96 ;
        RECT 65.76 2.48 66.24 2.96 ;
        RECT 0 7.92 0.48 8.4 ;
        RECT 65.76 7.92 66.24 8.4 ;
        RECT 0 13.36 0.48 13.84 ;
        RECT 65.76 13.36 66.24 13.84 ;
        RECT 0 18.8 0.48 19.28 ;
        RECT 65.76 18.8 66.24 19.28 ;
        RECT 0 24.24 0.48 24.72 ;
        RECT 65.76 24.24 66.24 24.72 ;
        RECT 0 29.68 0.48 30.16 ;
        RECT 65.76 29.68 66.24 30.16 ;
        RECT 0 35.12 0.48 35.6 ;
        RECT 65.76 35.12 66.24 35.6 ;
        RECT 0 40.56 0.48 41.04 ;
        RECT 65.76 40.56 66.24 41.04 ;
        RECT 0 46 0.48 46.48 ;
        RECT 65.76 46 66.24 46.48 ;
        RECT 0 51.44 0.48 51.92 ;
        RECT 65.76 51.44 66.24 51.92 ;
        RECT 0 56.88 0.48 57.36 ;
        RECT 65.76 56.88 66.24 57.36 ;
        RECT 0 62.32 0.48 62.8 ;
        RECT 65.76 62.32 66.24 62.8 ;
        RECT 0 67.76 0.48 68.24 ;
        RECT 65.76 67.76 66.24 68.24 ;
        RECT 0 73.2 0.48 73.68 ;
        RECT 65.76 73.2 66.24 73.68 ;
        RECT 0 78.64 0.48 79.12 ;
        RECT 65.76 78.64 66.24 79.12 ;
        RECT 0 84.08 0.48 84.56 ;
        RECT 65.76 84.08 66.24 84.56 ;
    END
  END VDD
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0 31.72 3.2 34.92 ;
        RECT 63.04 31.72 66.24 34.92 ;
        RECT 0 72.52 3.2 75.72 ;
        RECT 63.04 72.52 66.24 75.72 ;
      LAYER met4 ;
        RECT 25.46 0 26.06 0.6 ;
        RECT 54.9 0 55.5 0.6 ;
        RECT 25.46 86.44 26.06 87.04 ;
        RECT 54.9 86.44 55.5 87.04 ;
      LAYER met1 ;
        RECT 0 0 66.24 0.24 ;
        RECT 0 5.2 0.48 5.68 ;
        RECT 65.76 5.2 66.24 5.68 ;
        RECT 0 10.64 0.48 11.12 ;
        RECT 65.76 10.64 66.24 11.12 ;
        RECT 0 16.08 0.48 16.56 ;
        RECT 65.76 16.08 66.24 16.56 ;
        RECT 0 21.52 0.48 22 ;
        RECT 65.76 21.52 66.24 22 ;
        RECT 0 26.96 0.48 27.44 ;
        RECT 65.76 26.96 66.24 27.44 ;
        RECT 0 32.4 0.48 32.88 ;
        RECT 65.76 32.4 66.24 32.88 ;
        RECT 0 37.84 0.48 38.32 ;
        RECT 65.76 37.84 66.24 38.32 ;
        RECT 0 43.28 0.48 43.76 ;
        RECT 65.76 43.28 66.24 43.76 ;
        RECT 0 48.72 0.48 49.2 ;
        RECT 65.76 48.72 66.24 49.2 ;
        RECT 0 54.16 0.48 54.64 ;
        RECT 65.76 54.16 66.24 54.64 ;
        RECT 0 59.6 0.48 60.08 ;
        RECT 65.76 59.6 66.24 60.08 ;
        RECT 0 65.04 0.48 65.52 ;
        RECT 65.76 65.04 66.24 65.52 ;
        RECT 0 70.48 0.48 70.96 ;
        RECT 65.76 70.48 66.24 70.96 ;
        RECT 0 75.92 0.48 76.4 ;
        RECT 65.76 75.92 66.24 76.4 ;
        RECT 0 81.36 0.48 81.84 ;
        RECT 65.76 81.36 66.24 81.84 ;
        RECT 0 86.8 66.24 87.04 ;
    END
  END VSS
  PIN prog_clk__FEEDTHRU_1[0]
    DIRECTION OUTPUT ;
    USE CLOCK ;
    PORT
      LAYER met2 ;
        RECT 6.37 85.68 6.51 87.04 ;
    END
  END prog_clk__FEEDTHRU_1[0]
  OBS
    LAYER li1 ;
      RECT 0 86.955 66.24 87.125 ;
      RECT 65.32 84.235 66.24 84.405 ;
      RECT 0 84.235 3.68 84.405 ;
      RECT 65.32 81.515 66.24 81.685 ;
      RECT 0 81.515 1.84 81.685 ;
      RECT 65.32 78.795 66.24 78.965 ;
      RECT 0 78.795 1.84 78.965 ;
      RECT 65.32 76.075 66.24 76.245 ;
      RECT 0 76.075 1.84 76.245 ;
      RECT 65.32 73.355 66.24 73.525 ;
      RECT 0 73.355 1.84 73.525 ;
      RECT 65.32 70.635 66.24 70.805 ;
      RECT 0 70.635 1.84 70.805 ;
      RECT 65.32 67.915 66.24 68.085 ;
      RECT 0 67.915 1.84 68.085 ;
      RECT 65.32 65.195 66.24 65.365 ;
      RECT 0 65.195 1.84 65.365 ;
      RECT 65.32 62.475 66.24 62.645 ;
      RECT 0 62.475 3.68 62.645 ;
      RECT 65.32 59.755 66.24 59.925 ;
      RECT 0 59.755 3.68 59.925 ;
      RECT 65.32 57.035 66.24 57.205 ;
      RECT 0 57.035 1.84 57.205 ;
      RECT 65.32 54.315 66.24 54.485 ;
      RECT 0 54.315 1.84 54.485 ;
      RECT 65.32 51.595 66.24 51.765 ;
      RECT 0 51.595 1.84 51.765 ;
      RECT 65.32 48.875 66.24 49.045 ;
      RECT 0 48.875 1.84 49.045 ;
      RECT 65.32 46.155 66.24 46.325 ;
      RECT 0 46.155 1.84 46.325 ;
      RECT 65.32 43.435 66.24 43.605 ;
      RECT 0 43.435 1.84 43.605 ;
      RECT 65.32 40.715 66.24 40.885 ;
      RECT 0 40.715 1.84 40.885 ;
      RECT 62.56 37.995 66.24 38.165 ;
      RECT 0 37.995 1.84 38.165 ;
      RECT 62.56 35.275 66.24 35.445 ;
      RECT 0 35.275 1.84 35.445 ;
      RECT 65.32 32.555 66.24 32.725 ;
      RECT 0 32.555 1.84 32.725 ;
      RECT 65.32 29.835 66.24 30.005 ;
      RECT 0 29.835 1.84 30.005 ;
      RECT 65.32 27.115 66.24 27.285 ;
      RECT 0 27.115 1.84 27.285 ;
      RECT 65.32 24.395 66.24 24.565 ;
      RECT 0 24.395 1.84 24.565 ;
      RECT 65.32 21.675 66.24 21.845 ;
      RECT 0 21.675 1.84 21.845 ;
      RECT 65.32 18.955 66.24 19.125 ;
      RECT 0 18.955 1.84 19.125 ;
      RECT 64.4 16.235 66.24 16.405 ;
      RECT 0 16.235 1.84 16.405 ;
      RECT 64.4 13.515 66.24 13.685 ;
      RECT 0 13.515 1.84 13.685 ;
      RECT 65.32 10.795 66.24 10.965 ;
      RECT 0 10.795 1.84 10.965 ;
      RECT 65.32 8.075 66.24 8.245 ;
      RECT 0 8.075 1.84 8.245 ;
      RECT 65.78 5.355 66.24 5.525 ;
      RECT 0 5.355 3.68 5.525 ;
      RECT 65.78 2.635 66.24 2.805 ;
      RECT 0 2.635 3.68 2.805 ;
      RECT 0 -0.085 66.24 0.085 ;
    LAYER met3 ;
      POLYGON 55.365 87.205 55.365 87.2 55.58 87.2 55.58 86.88 55.365 86.88 55.365 86.875 55.035 86.875 55.035 86.88 54.82 86.88 54.82 87.2 55.035 87.2 55.035 87.205 ;
      POLYGON 25.925 87.205 25.925 87.2 26.14 87.2 26.14 86.88 25.925 86.88 25.925 86.875 25.595 86.875 25.595 86.88 25.38 86.88 25.38 87.2 25.595 87.2 25.595 87.205 ;
      POLYGON 14.41 71.55 14.41 71.25 1.23 71.25 1.23 71.53 1.78 71.53 1.78 71.55 ;
      POLYGON 1.99 45.03 1.99 44.35 4.29 44.35 4.29 44.05 1.69 44.05 1.69 44.33 1.78 44.33 1.78 45.03 ;
      POLYGON 6.59 37.55 6.59 37.25 1.99 37.25 1.99 36.57 1.78 36.57 1.78 37.27 1.69 37.27 1.69 37.55 ;
      POLYGON 55.365 0.165 55.365 0.16 55.58 0.16 55.58 -0.16 55.365 -0.16 55.365 -0.165 55.035 -0.165 55.035 -0.16 54.82 -0.16 54.82 0.16 55.035 0.16 55.035 0.165 ;
      POLYGON 25.925 0.165 25.925 0.16 26.14 0.16 26.14 -0.16 25.925 -0.16 25.925 -0.165 25.595 -0.165 25.595 -0.16 25.38 -0.16 25.38 0.16 25.595 0.16 25.595 0.165 ;
      POLYGON 65.84 86.64 65.84 84.19 64.46 84.19 64.46 83.09 65.84 83.09 65.84 82.83 64.46 82.83 64.46 81.73 65.84 81.73 65.84 80.79 64.46 80.79 64.46 79.69 65.84 79.69 65.84 79.43 64.46 79.43 64.46 78.33 65.84 78.33 65.84 78.07 64.46 78.07 64.46 76.97 65.84 76.97 65.84 76.71 64.46 76.71 64.46 75.61 65.84 75.61 65.84 75.35 64.46 75.35 64.46 74.25 65.84 74.25 65.84 73.99 64.46 73.99 64.46 72.89 65.84 72.89 65.84 72.63 64.46 72.63 64.46 71.53 65.84 71.53 65.84 71.27 64.46 71.27 64.46 70.17 65.84 70.17 65.84 69.91 64.46 69.91 64.46 68.81 65.84 68.81 65.84 68.55 64.46 68.55 64.46 67.45 65.84 67.45 65.84 67.19 64.46 67.19 64.46 66.09 65.84 66.09 65.84 65.83 64.46 65.83 64.46 64.73 65.84 64.73 65.84 64.47 64.46 64.47 64.46 63.37 65.84 63.37 65.84 62.43 64.46 62.43 64.46 61.33 65.84 61.33 65.84 60.39 64.46 60.39 64.46 59.29 65.84 59.29 65.84 59.03 64.46 59.03 64.46 57.93 65.84 57.93 65.84 56.99 64.46 56.99 64.46 55.89 65.84 55.89 65.84 54.95 64.46 54.95 64.46 53.85 65.84 53.85 65.84 52.91 64.46 52.91 64.46 51.81 65.84 51.81 65.84 51.55 64.46 51.55 64.46 50.45 65.84 50.45 65.84 50.19 64.46 50.19 64.46 49.09 65.84 49.09 65.84 48.83 64.46 48.83 64.46 47.73 65.84 47.73 65.84 46.79 64.46 46.79 64.46 45.69 65.84 45.69 65.84 45.43 64.46 45.43 64.46 44.33 65.84 44.33 65.84 44.07 64.46 44.07 64.46 42.97 65.84 42.97 65.84 42.71 64.46 42.71 64.46 41.61 65.84 41.61 65.84 41.35 64.46 41.35 64.46 40.25 65.84 40.25 65.84 39.99 64.46 39.99 64.46 38.89 65.84 38.89 65.84 37.95 64.46 37.95 64.46 36.85 65.84 36.85 65.84 36.59 64.46 36.59 64.46 35.49 65.84 35.49 65.84 35.23 64.46 35.23 64.46 34.13 65.84 34.13 65.84 33.87 64.46 33.87 64.46 32.77 65.84 32.77 65.84 31.83 64.46 31.83 64.46 30.73 65.84 30.73 65.84 30.47 64.46 30.47 64.46 29.37 65.84 29.37 65.84 28.43 64.46 28.43 64.46 27.33 65.84 27.33 65.84 26.39 64.46 26.39 64.46 25.29 65.84 25.29 65.84 25.03 64.46 25.03 64.46 23.93 65.84 23.93 65.84 23.67 64.46 23.67 64.46 22.57 65.84 22.57 65.84 22.31 64.46 22.31 64.46 21.21 65.84 21.21 65.84 20.27 64.46 20.27 64.46 19.17 65.84 19.17 65.84 18.91 64.46 18.91 64.46 17.81 65.84 17.81 65.84 17.55 64.46 17.55 64.46 16.45 65.84 16.45 65.84 16.19 64.46 16.19 64.46 15.09 65.84 15.09 65.84 14.15 64.46 14.15 64.46 13.05 65.84 13.05 65.84 12.11 64.46 12.11 64.46 11.01 65.84 11.01 65.84 10.75 64.46 10.75 64.46 9.65 65.84 9.65 65.84 9.39 64.46 9.39 64.46 8.29 65.84 8.29 65.84 8.03 64.46 8.03 64.46 6.93 65.84 6.93 65.84 6.67 64.46 6.67 64.46 5.57 65.84 5.57 65.84 0.4 0.4 0.4 0.4 8.97 1.78 8.97 1.78 10.07 0.4 10.07 0.4 10.33 1.78 10.33 1.78 11.43 0.4 11.43 0.4 11.69 1.78 11.69 1.78 12.79 0.4 12.79 0.4 13.05 1.78 13.05 1.78 14.15 0.4 14.15 0.4 14.41 1.78 14.41 1.78 15.51 0.4 15.51 0.4 15.77 1.78 15.77 1.78 16.87 0.4 16.87 0.4 17.13 1.78 17.13 1.78 18.23 0.4 18.23 0.4 18.49 1.78 18.49 1.78 19.59 0.4 19.59 0.4 19.85 1.78 19.85 1.78 20.95 0.4 20.95 0.4 21.21 1.78 21.21 1.78 22.31 0.4 22.31 0.4 22.57 1.78 22.57 1.78 23.67 0.4 23.67 0.4 23.93 1.78 23.93 1.78 25.03 0.4 25.03 0.4 25.97 1.78 25.97 1.78 27.07 0.4 27.07 0.4 28.01 1.78 28.01 1.78 29.11 0.4 29.11 0.4 29.37 1.78 29.37 1.78 30.47 0.4 30.47 0.4 30.73 1.78 30.73 1.78 31.83 0.4 31.83 0.4 32.09 1.78 32.09 1.78 33.19 0.4 33.19 0.4 33.45 1.78 33.45 1.78 34.55 0.4 34.55 0.4 34.81 1.78 34.81 1.78 35.91 0.4 35.91 0.4 36.17 1.78 36.17 1.78 37.27 0.4 37.27 0.4 37.53 1.78 37.53 1.78 38.63 0.4 38.63 0.4 38.89 1.78 38.89 1.78 39.99 0.4 39.99 0.4 40.25 1.78 40.25 1.78 41.35 0.4 41.35 0.4 41.61 1.78 41.61 1.78 42.71 0.4 42.71 0.4 42.97 1.78 42.97 1.78 44.07 0.4 44.07 0.4 44.33 1.78 44.33 1.78 45.43 0.4 45.43 0.4 45.69 1.78 45.69 1.78 46.79 0.4 46.79 0.4 47.05 1.78 47.05 1.78 48.15 0.4 48.15 0.4 48.41 1.78 48.41 1.78 49.51 0.4 49.51 0.4 49.77 1.78 49.77 1.78 50.87 0.4 50.87 0.4 51.81 1.78 51.81 1.78 52.91 0.4 52.91 0.4 53.17 1.78 53.17 1.78 54.27 0.4 54.27 0.4 54.53 1.78 54.53 1.78 55.63 0.4 55.63 0.4 56.57 1.78 56.57 1.78 57.67 0.4 57.67 0.4 57.93 1.78 57.93 1.78 59.03 0.4 59.03 0.4 59.29 1.78 59.29 1.78 60.39 0.4 60.39 0.4 61.33 1.78 61.33 1.78 62.43 0.4 62.43 0.4 62.69 1.78 62.69 1.78 63.79 0.4 63.79 0.4 64.73 1.78 64.73 1.78 65.83 0.4 65.83 0.4 66.09 1.78 66.09 1.78 67.19 0.4 67.19 0.4 67.45 1.78 67.45 1.78 68.55 0.4 68.55 0.4 68.81 1.78 68.81 1.78 69.91 0.4 69.91 0.4 70.17 1.78 70.17 1.78 71.27 0.4 71.27 0.4 71.53 1.78 71.53 1.78 72.63 0.4 72.63 0.4 72.89 1.78 72.89 1.78 73.99 0.4 73.99 0.4 74.25 1.78 74.25 1.78 75.35 0.4 75.35 0.4 75.61 1.78 75.61 1.78 76.71 0.4 76.71 0.4 76.97 1.78 76.97 1.78 78.07 0.4 78.07 0.4 78.33 1.78 78.33 1.78 79.43 0.4 79.43 0.4 79.69 1.78 79.69 1.78 80.79 0.4 80.79 0.4 81.73 1.78 81.73 1.78 82.83 0.4 82.83 0.4 83.09 1.78 83.09 1.78 84.19 0.4 84.19 0.4 86.64 ;
    LAYER met2 ;
      RECT 55.06 86.855 55.34 87.225 ;
      RECT 25.62 86.855 25.9 87.225 ;
      RECT 55.06 -0.185 55.34 0.185 ;
      RECT 25.62 -0.185 25.9 0.185 ;
      POLYGON 65.96 86.76 65.96 0.28 61.53 0.28 61.53 1.64 60.83 1.64 60.83 0.28 56.47 0.28 56.47 1.64 55.77 1.64 55.77 0.28 44.51 0.28 44.51 1.64 43.81 1.64 43.81 0.28 43.59 0.28 43.59 1.64 42.89 1.64 42.89 0.28 42.67 0.28 42.67 1.64 41.97 1.64 41.97 0.28 41.29 0.28 41.29 1.64 40.59 1.64 40.59 0.28 39.91 0.28 39.91 1.64 39.21 1.64 39.21 0.28 34.85 0.28 34.85 1.64 34.15 1.64 34.15 0.28 33.93 0.28 33.93 1.64 33.23 1.64 33.23 0.28 31.63 0.28 31.63 1.64 30.93 1.64 30.93 0.28 30.25 0.28 30.25 1.64 29.55 1.64 29.55 0.28 29.33 0.28 29.33 1.64 28.63 1.64 28.63 0.28 28.41 0.28 28.41 1.64 27.71 1.64 27.71 0.28 27.03 0.28 27.03 1.64 26.33 1.64 26.33 0.28 25.19 0.28 25.19 1.64 24.49 1.64 24.49 0.28 24.27 0.28 24.27 1.64 23.57 1.64 23.57 0.28 21.05 0.28 21.05 1.64 20.35 1.64 20.35 0.28 14.61 0.28 14.61 1.64 13.91 1.64 13.91 0.28 13.23 0.28 13.23 1.64 12.53 1.64 12.53 0.28 9.09 0.28 9.09 1.64 8.39 1.64 8.39 0.28 8.17 0.28 8.17 1.64 7.47 1.64 7.47 0.28 4.49 0.28 4.49 1.64 3.79 1.64 3.79 0.28 0.28 0.28 0.28 86.76 6.09 86.76 6.09 85.4 6.79 85.4 6.79 86.76 11.15 86.76 11.15 85.4 11.85 85.4 11.85 86.76 12.07 86.76 12.07 85.4 12.77 85.4 12.77 86.76 13.91 86.76 13.91 85.4 14.61 85.4 14.61 86.76 63.59 86.76 63.59 85.4 64.29 85.4 64.29 86.76 ;
    LAYER met1 ;
      POLYGON 65.96 86.52 65.96 84.84 65.48 84.84 65.48 83.8 65.96 83.8 65.96 82.12 65.48 82.12 65.48 81.08 65.96 81.08 65.96 79.4 65.48 79.4 65.48 78.36 65.96 78.36 65.96 76.68 65.48 76.68 65.48 75.64 65.96 75.64 65.96 73.96 65.48 73.96 65.48 72.92 65.96 72.92 65.96 71.24 65.48 71.24 65.48 70.2 65.96 70.2 65.96 68.52 65.48 68.52 65.48 67.48 65.96 67.48 65.96 65.8 65.48 65.8 65.48 64.76 65.96 64.76 65.96 63.08 65.48 63.08 65.48 62.04 65.96 62.04 65.96 60.36 65.48 60.36 65.48 59.32 65.96 59.32 65.96 57.64 65.48 57.64 65.48 56.6 65.96 56.6 65.96 54.92 65.48 54.92 65.48 53.88 65.96 53.88 65.96 52.2 65.48 52.2 65.48 51.16 65.96 51.16 65.96 49.48 65.48 49.48 65.48 48.44 65.96 48.44 65.96 46.76 65.48 46.76 65.48 45.72 65.96 45.72 65.96 44.04 65.48 44.04 65.48 43 65.96 43 65.96 41.32 65.48 41.32 65.48 40.28 65.96 40.28 65.96 38.6 65.48 38.6 65.48 37.56 65.96 37.56 65.96 35.88 65.48 35.88 65.48 34.84 65.96 34.84 65.96 33.16 65.48 33.16 65.48 32.12 65.96 32.12 65.96 30.44 65.48 30.44 65.48 29.4 65.96 29.4 65.96 27.72 65.48 27.72 65.48 26.68 65.96 26.68 65.96 25 65.48 25 65.48 23.96 65.96 23.96 65.96 22.28 65.48 22.28 65.48 21.24 65.96 21.24 65.96 19.56 65.48 19.56 65.48 18.52 65.96 18.52 65.96 16.84 65.48 16.84 65.48 15.8 65.96 15.8 65.96 14.12 65.48 14.12 65.48 13.08 65.96 13.08 65.96 11.4 65.48 11.4 65.48 10.36 65.96 10.36 65.96 8.68 65.48 8.68 65.48 7.64 65.96 7.64 65.96 5.96 65.48 5.96 65.48 4.92 65.96 4.92 65.96 3.24 65.48 3.24 65.48 2.2 65.96 2.2 65.96 0.52 0.28 0.52 0.28 2.2 0.76 2.2 0.76 3.24 0.28 3.24 0.28 4.92 0.76 4.92 0.76 5.96 0.28 5.96 0.28 7.64 0.76 7.64 0.76 8.68 0.28 8.68 0.28 10.36 0.76 10.36 0.76 11.4 0.28 11.4 0.28 13.08 0.76 13.08 0.76 14.12 0.28 14.12 0.28 15.8 0.76 15.8 0.76 16.84 0.28 16.84 0.28 18.52 0.76 18.52 0.76 19.56 0.28 19.56 0.28 21.24 0.76 21.24 0.76 22.28 0.28 22.28 0.28 23.96 0.76 23.96 0.76 25 0.28 25 0.28 26.68 0.76 26.68 0.76 27.72 0.28 27.72 0.28 29.4 0.76 29.4 0.76 30.44 0.28 30.44 0.28 32.12 0.76 32.12 0.76 33.16 0.28 33.16 0.28 34.84 0.76 34.84 0.76 35.88 0.28 35.88 0.28 37.56 0.76 37.56 0.76 38.6 0.28 38.6 0.28 40.28 0.76 40.28 0.76 41.32 0.28 41.32 0.28 43 0.76 43 0.76 44.04 0.28 44.04 0.28 45.72 0.76 45.72 0.76 46.76 0.28 46.76 0.28 48.44 0.76 48.44 0.76 49.48 0.28 49.48 0.28 51.16 0.76 51.16 0.76 52.2 0.28 52.2 0.28 53.88 0.76 53.88 0.76 54.92 0.28 54.92 0.28 56.6 0.76 56.6 0.76 57.64 0.28 57.64 0.28 59.32 0.76 59.32 0.76 60.36 0.28 60.36 0.28 62.04 0.76 62.04 0.76 63.08 0.28 63.08 0.28 64.76 0.76 64.76 0.76 65.8 0.28 65.8 0.28 67.48 0.76 67.48 0.76 68.52 0.28 68.52 0.28 70.2 0.76 70.2 0.76 71.24 0.28 71.24 0.28 72.92 0.76 72.92 0.76 73.96 0.28 73.96 0.28 75.64 0.76 75.64 0.76 76.68 0.28 76.68 0.28 78.36 0.76 78.36 0.76 79.4 0.28 79.4 0.28 81.08 0.76 81.08 0.76 82.12 0.28 82.12 0.28 83.8 0.76 83.8 0.76 84.84 0.28 84.84 0.28 86.52 ;
    LAYER met4 ;
      POLYGON 65.84 86.64 65.84 0.4 55.9 0.4 55.9 1 54.5 1 54.5 0.4 41.18 0.4 41.18 1 39.78 1 39.78 0.4 26.46 0.4 26.46 1 25.06 1 25.06 0.4 11.74 0.4 11.74 1 10.34 1 10.34 0.4 0.4 0.4 0.4 86.64 10.34 86.64 10.34 86.04 11.74 86.04 11.74 86.64 25.06 86.64 25.06 86.04 26.46 86.04 26.46 86.64 39.78 86.64 39.78 86.04 41.18 86.04 41.18 86.64 54.5 86.64 54.5 86.04 55.9 86.04 55.9 86.64 ;
    LAYER met5 ;
      POLYGON 64.64 85.44 64.64 77.32 61.44 77.32 61.44 70.92 64.64 70.92 64.64 56.92 61.44 56.92 61.44 50.52 64.64 50.52 64.64 36.52 61.44 36.52 61.44 30.12 64.64 30.12 64.64 16.12 61.44 16.12 61.44 9.72 64.64 9.72 64.64 1.6 1.6 1.6 1.6 9.72 4.8 9.72 4.8 16.12 1.6 16.12 1.6 30.12 4.8 30.12 4.8 36.52 1.6 36.52 1.6 50.52 4.8 50.52 4.8 56.92 1.6 56.92 1.6 70.92 4.8 70.92 4.8 77.32 1.6 77.32 1.6 85.44 ;
    LAYER li1 ;
      RECT 0.17 0.17 66.07 86.87 ;
    LAYER mcon ;
      RECT 65.925 86.955 66.095 87.125 ;
      RECT 65.465 86.955 65.635 87.125 ;
      RECT 65.005 86.955 65.175 87.125 ;
      RECT 64.545 86.955 64.715 87.125 ;
      RECT 64.085 86.955 64.255 87.125 ;
      RECT 63.625 86.955 63.795 87.125 ;
      RECT 63.165 86.955 63.335 87.125 ;
      RECT 62.705 86.955 62.875 87.125 ;
      RECT 62.245 86.955 62.415 87.125 ;
      RECT 61.785 86.955 61.955 87.125 ;
      RECT 61.325 86.955 61.495 87.125 ;
      RECT 60.865 86.955 61.035 87.125 ;
      RECT 60.405 86.955 60.575 87.125 ;
      RECT 59.945 86.955 60.115 87.125 ;
      RECT 59.485 86.955 59.655 87.125 ;
      RECT 59.025 86.955 59.195 87.125 ;
      RECT 58.565 86.955 58.735 87.125 ;
      RECT 58.105 86.955 58.275 87.125 ;
      RECT 57.645 86.955 57.815 87.125 ;
      RECT 57.185 86.955 57.355 87.125 ;
      RECT 56.725 86.955 56.895 87.125 ;
      RECT 56.265 86.955 56.435 87.125 ;
      RECT 55.805 86.955 55.975 87.125 ;
      RECT 55.345 86.955 55.515 87.125 ;
      RECT 54.885 86.955 55.055 87.125 ;
      RECT 54.425 86.955 54.595 87.125 ;
      RECT 53.965 86.955 54.135 87.125 ;
      RECT 53.505 86.955 53.675 87.125 ;
      RECT 53.045 86.955 53.215 87.125 ;
      RECT 52.585 86.955 52.755 87.125 ;
      RECT 52.125 86.955 52.295 87.125 ;
      RECT 51.665 86.955 51.835 87.125 ;
      RECT 51.205 86.955 51.375 87.125 ;
      RECT 50.745 86.955 50.915 87.125 ;
      RECT 50.285 86.955 50.455 87.125 ;
      RECT 49.825 86.955 49.995 87.125 ;
      RECT 49.365 86.955 49.535 87.125 ;
      RECT 48.905 86.955 49.075 87.125 ;
      RECT 48.445 86.955 48.615 87.125 ;
      RECT 47.985 86.955 48.155 87.125 ;
      RECT 47.525 86.955 47.695 87.125 ;
      RECT 47.065 86.955 47.235 87.125 ;
      RECT 46.605 86.955 46.775 87.125 ;
      RECT 46.145 86.955 46.315 87.125 ;
      RECT 45.685 86.955 45.855 87.125 ;
      RECT 45.225 86.955 45.395 87.125 ;
      RECT 44.765 86.955 44.935 87.125 ;
      RECT 44.305 86.955 44.475 87.125 ;
      RECT 43.845 86.955 44.015 87.125 ;
      RECT 43.385 86.955 43.555 87.125 ;
      RECT 42.925 86.955 43.095 87.125 ;
      RECT 42.465 86.955 42.635 87.125 ;
      RECT 42.005 86.955 42.175 87.125 ;
      RECT 41.545 86.955 41.715 87.125 ;
      RECT 41.085 86.955 41.255 87.125 ;
      RECT 40.625 86.955 40.795 87.125 ;
      RECT 40.165 86.955 40.335 87.125 ;
      RECT 39.705 86.955 39.875 87.125 ;
      RECT 39.245 86.955 39.415 87.125 ;
      RECT 38.785 86.955 38.955 87.125 ;
      RECT 38.325 86.955 38.495 87.125 ;
      RECT 37.865 86.955 38.035 87.125 ;
      RECT 37.405 86.955 37.575 87.125 ;
      RECT 36.945 86.955 37.115 87.125 ;
      RECT 36.485 86.955 36.655 87.125 ;
      RECT 36.025 86.955 36.195 87.125 ;
      RECT 35.565 86.955 35.735 87.125 ;
      RECT 35.105 86.955 35.275 87.125 ;
      RECT 34.645 86.955 34.815 87.125 ;
      RECT 34.185 86.955 34.355 87.125 ;
      RECT 33.725 86.955 33.895 87.125 ;
      RECT 33.265 86.955 33.435 87.125 ;
      RECT 32.805 86.955 32.975 87.125 ;
      RECT 32.345 86.955 32.515 87.125 ;
      RECT 31.885 86.955 32.055 87.125 ;
      RECT 31.425 86.955 31.595 87.125 ;
      RECT 30.965 86.955 31.135 87.125 ;
      RECT 30.505 86.955 30.675 87.125 ;
      RECT 30.045 86.955 30.215 87.125 ;
      RECT 29.585 86.955 29.755 87.125 ;
      RECT 29.125 86.955 29.295 87.125 ;
      RECT 28.665 86.955 28.835 87.125 ;
      RECT 28.205 86.955 28.375 87.125 ;
      RECT 27.745 86.955 27.915 87.125 ;
      RECT 27.285 86.955 27.455 87.125 ;
      RECT 26.825 86.955 26.995 87.125 ;
      RECT 26.365 86.955 26.535 87.125 ;
      RECT 25.905 86.955 26.075 87.125 ;
      RECT 25.445 86.955 25.615 87.125 ;
      RECT 24.985 86.955 25.155 87.125 ;
      RECT 24.525 86.955 24.695 87.125 ;
      RECT 24.065 86.955 24.235 87.125 ;
      RECT 23.605 86.955 23.775 87.125 ;
      RECT 23.145 86.955 23.315 87.125 ;
      RECT 22.685 86.955 22.855 87.125 ;
      RECT 22.225 86.955 22.395 87.125 ;
      RECT 21.765 86.955 21.935 87.125 ;
      RECT 21.305 86.955 21.475 87.125 ;
      RECT 20.845 86.955 21.015 87.125 ;
      RECT 20.385 86.955 20.555 87.125 ;
      RECT 19.925 86.955 20.095 87.125 ;
      RECT 19.465 86.955 19.635 87.125 ;
      RECT 19.005 86.955 19.175 87.125 ;
      RECT 18.545 86.955 18.715 87.125 ;
      RECT 18.085 86.955 18.255 87.125 ;
      RECT 17.625 86.955 17.795 87.125 ;
      RECT 17.165 86.955 17.335 87.125 ;
      RECT 16.705 86.955 16.875 87.125 ;
      RECT 16.245 86.955 16.415 87.125 ;
      RECT 15.785 86.955 15.955 87.125 ;
      RECT 15.325 86.955 15.495 87.125 ;
      RECT 14.865 86.955 15.035 87.125 ;
      RECT 14.405 86.955 14.575 87.125 ;
      RECT 13.945 86.955 14.115 87.125 ;
      RECT 13.485 86.955 13.655 87.125 ;
      RECT 13.025 86.955 13.195 87.125 ;
      RECT 12.565 86.955 12.735 87.125 ;
      RECT 12.105 86.955 12.275 87.125 ;
      RECT 11.645 86.955 11.815 87.125 ;
      RECT 11.185 86.955 11.355 87.125 ;
      RECT 10.725 86.955 10.895 87.125 ;
      RECT 10.265 86.955 10.435 87.125 ;
      RECT 9.805 86.955 9.975 87.125 ;
      RECT 9.345 86.955 9.515 87.125 ;
      RECT 8.885 86.955 9.055 87.125 ;
      RECT 8.425 86.955 8.595 87.125 ;
      RECT 7.965 86.955 8.135 87.125 ;
      RECT 7.505 86.955 7.675 87.125 ;
      RECT 7.045 86.955 7.215 87.125 ;
      RECT 6.585 86.955 6.755 87.125 ;
      RECT 6.125 86.955 6.295 87.125 ;
      RECT 5.665 86.955 5.835 87.125 ;
      RECT 5.205 86.955 5.375 87.125 ;
      RECT 4.745 86.955 4.915 87.125 ;
      RECT 4.285 86.955 4.455 87.125 ;
      RECT 3.825 86.955 3.995 87.125 ;
      RECT 3.365 86.955 3.535 87.125 ;
      RECT 2.905 86.955 3.075 87.125 ;
      RECT 2.445 86.955 2.615 87.125 ;
      RECT 1.985 86.955 2.155 87.125 ;
      RECT 1.525 86.955 1.695 87.125 ;
      RECT 1.065 86.955 1.235 87.125 ;
      RECT 0.605 86.955 0.775 87.125 ;
      RECT 0.145 86.955 0.315 87.125 ;
      RECT 65.925 84.235 66.095 84.405 ;
      RECT 65.465 84.235 65.635 84.405 ;
      RECT 0.605 84.235 0.775 84.405 ;
      RECT 0.145 84.235 0.315 84.405 ;
      RECT 65.925 81.515 66.095 81.685 ;
      RECT 65.465 81.515 65.635 81.685 ;
      RECT 0.605 81.515 0.775 81.685 ;
      RECT 0.145 81.515 0.315 81.685 ;
      RECT 65.925 78.795 66.095 78.965 ;
      RECT 65.465 78.795 65.635 78.965 ;
      RECT 0.605 78.795 0.775 78.965 ;
      RECT 0.145 78.795 0.315 78.965 ;
      RECT 65.925 76.075 66.095 76.245 ;
      RECT 65.465 76.075 65.635 76.245 ;
      RECT 0.605 76.075 0.775 76.245 ;
      RECT 0.145 76.075 0.315 76.245 ;
      RECT 65.925 73.355 66.095 73.525 ;
      RECT 65.465 73.355 65.635 73.525 ;
      RECT 0.605 73.355 0.775 73.525 ;
      RECT 0.145 73.355 0.315 73.525 ;
      RECT 65.925 70.635 66.095 70.805 ;
      RECT 65.465 70.635 65.635 70.805 ;
      RECT 0.605 70.635 0.775 70.805 ;
      RECT 0.145 70.635 0.315 70.805 ;
      RECT 65.925 67.915 66.095 68.085 ;
      RECT 65.465 67.915 65.635 68.085 ;
      RECT 0.605 67.915 0.775 68.085 ;
      RECT 0.145 67.915 0.315 68.085 ;
      RECT 65.925 65.195 66.095 65.365 ;
      RECT 65.465 65.195 65.635 65.365 ;
      RECT 0.605 65.195 0.775 65.365 ;
      RECT 0.145 65.195 0.315 65.365 ;
      RECT 65.925 62.475 66.095 62.645 ;
      RECT 65.465 62.475 65.635 62.645 ;
      RECT 0.605 62.475 0.775 62.645 ;
      RECT 0.145 62.475 0.315 62.645 ;
      RECT 65.925 59.755 66.095 59.925 ;
      RECT 65.465 59.755 65.635 59.925 ;
      RECT 0.605 59.755 0.775 59.925 ;
      RECT 0.145 59.755 0.315 59.925 ;
      RECT 65.925 57.035 66.095 57.205 ;
      RECT 65.465 57.035 65.635 57.205 ;
      RECT 0.605 57.035 0.775 57.205 ;
      RECT 0.145 57.035 0.315 57.205 ;
      RECT 65.925 54.315 66.095 54.485 ;
      RECT 65.465 54.315 65.635 54.485 ;
      RECT 0.605 54.315 0.775 54.485 ;
      RECT 0.145 54.315 0.315 54.485 ;
      RECT 65.925 51.595 66.095 51.765 ;
      RECT 65.465 51.595 65.635 51.765 ;
      RECT 0.605 51.595 0.775 51.765 ;
      RECT 0.145 51.595 0.315 51.765 ;
      RECT 65.925 48.875 66.095 49.045 ;
      RECT 65.465 48.875 65.635 49.045 ;
      RECT 0.605 48.875 0.775 49.045 ;
      RECT 0.145 48.875 0.315 49.045 ;
      RECT 65.925 46.155 66.095 46.325 ;
      RECT 65.465 46.155 65.635 46.325 ;
      RECT 0.605 46.155 0.775 46.325 ;
      RECT 0.145 46.155 0.315 46.325 ;
      RECT 65.925 43.435 66.095 43.605 ;
      RECT 65.465 43.435 65.635 43.605 ;
      RECT 0.605 43.435 0.775 43.605 ;
      RECT 0.145 43.435 0.315 43.605 ;
      RECT 65.925 40.715 66.095 40.885 ;
      RECT 65.465 40.715 65.635 40.885 ;
      RECT 0.605 40.715 0.775 40.885 ;
      RECT 0.145 40.715 0.315 40.885 ;
      RECT 65.925 37.995 66.095 38.165 ;
      RECT 65.465 37.995 65.635 38.165 ;
      RECT 0.605 37.995 0.775 38.165 ;
      RECT 0.145 37.995 0.315 38.165 ;
      RECT 65.925 35.275 66.095 35.445 ;
      RECT 65.465 35.275 65.635 35.445 ;
      RECT 0.605 35.275 0.775 35.445 ;
      RECT 0.145 35.275 0.315 35.445 ;
      RECT 65.925 32.555 66.095 32.725 ;
      RECT 65.465 32.555 65.635 32.725 ;
      RECT 0.605 32.555 0.775 32.725 ;
      RECT 0.145 32.555 0.315 32.725 ;
      RECT 65.925 29.835 66.095 30.005 ;
      RECT 65.465 29.835 65.635 30.005 ;
      RECT 0.605 29.835 0.775 30.005 ;
      RECT 0.145 29.835 0.315 30.005 ;
      RECT 65.925 27.115 66.095 27.285 ;
      RECT 65.465 27.115 65.635 27.285 ;
      RECT 0.605 27.115 0.775 27.285 ;
      RECT 0.145 27.115 0.315 27.285 ;
      RECT 65.925 24.395 66.095 24.565 ;
      RECT 65.465 24.395 65.635 24.565 ;
      RECT 0.605 24.395 0.775 24.565 ;
      RECT 0.145 24.395 0.315 24.565 ;
      RECT 65.925 21.675 66.095 21.845 ;
      RECT 65.465 21.675 65.635 21.845 ;
      RECT 0.605 21.675 0.775 21.845 ;
      RECT 0.145 21.675 0.315 21.845 ;
      RECT 65.925 18.955 66.095 19.125 ;
      RECT 65.465 18.955 65.635 19.125 ;
      RECT 0.605 18.955 0.775 19.125 ;
      RECT 0.145 18.955 0.315 19.125 ;
      RECT 65.925 16.235 66.095 16.405 ;
      RECT 65.465 16.235 65.635 16.405 ;
      RECT 0.605 16.235 0.775 16.405 ;
      RECT 0.145 16.235 0.315 16.405 ;
      RECT 65.925 13.515 66.095 13.685 ;
      RECT 65.465 13.515 65.635 13.685 ;
      RECT 0.605 13.515 0.775 13.685 ;
      RECT 0.145 13.515 0.315 13.685 ;
      RECT 65.925 10.795 66.095 10.965 ;
      RECT 65.465 10.795 65.635 10.965 ;
      RECT 0.605 10.795 0.775 10.965 ;
      RECT 0.145 10.795 0.315 10.965 ;
      RECT 65.925 8.075 66.095 8.245 ;
      RECT 65.465 8.075 65.635 8.245 ;
      RECT 0.605 8.075 0.775 8.245 ;
      RECT 0.145 8.075 0.315 8.245 ;
      RECT 65.925 5.355 66.095 5.525 ;
      RECT 65.465 5.355 65.635 5.525 ;
      RECT 0.605 5.355 0.775 5.525 ;
      RECT 0.145 5.355 0.315 5.525 ;
      RECT 65.925 2.635 66.095 2.805 ;
      RECT 65.465 2.635 65.635 2.805 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 65.925 -0.085 66.095 0.085 ;
      RECT 65.465 -0.085 65.635 0.085 ;
      RECT 65.005 -0.085 65.175 0.085 ;
      RECT 64.545 -0.085 64.715 0.085 ;
      RECT 64.085 -0.085 64.255 0.085 ;
      RECT 63.625 -0.085 63.795 0.085 ;
      RECT 63.165 -0.085 63.335 0.085 ;
      RECT 62.705 -0.085 62.875 0.085 ;
      RECT 62.245 -0.085 62.415 0.085 ;
      RECT 61.785 -0.085 61.955 0.085 ;
      RECT 61.325 -0.085 61.495 0.085 ;
      RECT 60.865 -0.085 61.035 0.085 ;
      RECT 60.405 -0.085 60.575 0.085 ;
      RECT 59.945 -0.085 60.115 0.085 ;
      RECT 59.485 -0.085 59.655 0.085 ;
      RECT 59.025 -0.085 59.195 0.085 ;
      RECT 58.565 -0.085 58.735 0.085 ;
      RECT 58.105 -0.085 58.275 0.085 ;
      RECT 57.645 -0.085 57.815 0.085 ;
      RECT 57.185 -0.085 57.355 0.085 ;
      RECT 56.725 -0.085 56.895 0.085 ;
      RECT 56.265 -0.085 56.435 0.085 ;
      RECT 55.805 -0.085 55.975 0.085 ;
      RECT 55.345 -0.085 55.515 0.085 ;
      RECT 54.885 -0.085 55.055 0.085 ;
      RECT 54.425 -0.085 54.595 0.085 ;
      RECT 53.965 -0.085 54.135 0.085 ;
      RECT 53.505 -0.085 53.675 0.085 ;
      RECT 53.045 -0.085 53.215 0.085 ;
      RECT 52.585 -0.085 52.755 0.085 ;
      RECT 52.125 -0.085 52.295 0.085 ;
      RECT 51.665 -0.085 51.835 0.085 ;
      RECT 51.205 -0.085 51.375 0.085 ;
      RECT 50.745 -0.085 50.915 0.085 ;
      RECT 50.285 -0.085 50.455 0.085 ;
      RECT 49.825 -0.085 49.995 0.085 ;
      RECT 49.365 -0.085 49.535 0.085 ;
      RECT 48.905 -0.085 49.075 0.085 ;
      RECT 48.445 -0.085 48.615 0.085 ;
      RECT 47.985 -0.085 48.155 0.085 ;
      RECT 47.525 -0.085 47.695 0.085 ;
      RECT 47.065 -0.085 47.235 0.085 ;
      RECT 46.605 -0.085 46.775 0.085 ;
      RECT 46.145 -0.085 46.315 0.085 ;
      RECT 45.685 -0.085 45.855 0.085 ;
      RECT 45.225 -0.085 45.395 0.085 ;
      RECT 44.765 -0.085 44.935 0.085 ;
      RECT 44.305 -0.085 44.475 0.085 ;
      RECT 43.845 -0.085 44.015 0.085 ;
      RECT 43.385 -0.085 43.555 0.085 ;
      RECT 42.925 -0.085 43.095 0.085 ;
      RECT 42.465 -0.085 42.635 0.085 ;
      RECT 42.005 -0.085 42.175 0.085 ;
      RECT 41.545 -0.085 41.715 0.085 ;
      RECT 41.085 -0.085 41.255 0.085 ;
      RECT 40.625 -0.085 40.795 0.085 ;
      RECT 40.165 -0.085 40.335 0.085 ;
      RECT 39.705 -0.085 39.875 0.085 ;
      RECT 39.245 -0.085 39.415 0.085 ;
      RECT 38.785 -0.085 38.955 0.085 ;
      RECT 38.325 -0.085 38.495 0.085 ;
      RECT 37.865 -0.085 38.035 0.085 ;
      RECT 37.405 -0.085 37.575 0.085 ;
      RECT 36.945 -0.085 37.115 0.085 ;
      RECT 36.485 -0.085 36.655 0.085 ;
      RECT 36.025 -0.085 36.195 0.085 ;
      RECT 35.565 -0.085 35.735 0.085 ;
      RECT 35.105 -0.085 35.275 0.085 ;
      RECT 34.645 -0.085 34.815 0.085 ;
      RECT 34.185 -0.085 34.355 0.085 ;
      RECT 33.725 -0.085 33.895 0.085 ;
      RECT 33.265 -0.085 33.435 0.085 ;
      RECT 32.805 -0.085 32.975 0.085 ;
      RECT 32.345 -0.085 32.515 0.085 ;
      RECT 31.885 -0.085 32.055 0.085 ;
      RECT 31.425 -0.085 31.595 0.085 ;
      RECT 30.965 -0.085 31.135 0.085 ;
      RECT 30.505 -0.085 30.675 0.085 ;
      RECT 30.045 -0.085 30.215 0.085 ;
      RECT 29.585 -0.085 29.755 0.085 ;
      RECT 29.125 -0.085 29.295 0.085 ;
      RECT 28.665 -0.085 28.835 0.085 ;
      RECT 28.205 -0.085 28.375 0.085 ;
      RECT 27.745 -0.085 27.915 0.085 ;
      RECT 27.285 -0.085 27.455 0.085 ;
      RECT 26.825 -0.085 26.995 0.085 ;
      RECT 26.365 -0.085 26.535 0.085 ;
      RECT 25.905 -0.085 26.075 0.085 ;
      RECT 25.445 -0.085 25.615 0.085 ;
      RECT 24.985 -0.085 25.155 0.085 ;
      RECT 24.525 -0.085 24.695 0.085 ;
      RECT 24.065 -0.085 24.235 0.085 ;
      RECT 23.605 -0.085 23.775 0.085 ;
      RECT 23.145 -0.085 23.315 0.085 ;
      RECT 22.685 -0.085 22.855 0.085 ;
      RECT 22.225 -0.085 22.395 0.085 ;
      RECT 21.765 -0.085 21.935 0.085 ;
      RECT 21.305 -0.085 21.475 0.085 ;
      RECT 20.845 -0.085 21.015 0.085 ;
      RECT 20.385 -0.085 20.555 0.085 ;
      RECT 19.925 -0.085 20.095 0.085 ;
      RECT 19.465 -0.085 19.635 0.085 ;
      RECT 19.005 -0.085 19.175 0.085 ;
      RECT 18.545 -0.085 18.715 0.085 ;
      RECT 18.085 -0.085 18.255 0.085 ;
      RECT 17.625 -0.085 17.795 0.085 ;
      RECT 17.165 -0.085 17.335 0.085 ;
      RECT 16.705 -0.085 16.875 0.085 ;
      RECT 16.245 -0.085 16.415 0.085 ;
      RECT 15.785 -0.085 15.955 0.085 ;
      RECT 15.325 -0.085 15.495 0.085 ;
      RECT 14.865 -0.085 15.035 0.085 ;
      RECT 14.405 -0.085 14.575 0.085 ;
      RECT 13.945 -0.085 14.115 0.085 ;
      RECT 13.485 -0.085 13.655 0.085 ;
      RECT 13.025 -0.085 13.195 0.085 ;
      RECT 12.565 -0.085 12.735 0.085 ;
      RECT 12.105 -0.085 12.275 0.085 ;
      RECT 11.645 -0.085 11.815 0.085 ;
      RECT 11.185 -0.085 11.355 0.085 ;
      RECT 10.725 -0.085 10.895 0.085 ;
      RECT 10.265 -0.085 10.435 0.085 ;
      RECT 9.805 -0.085 9.975 0.085 ;
      RECT 9.345 -0.085 9.515 0.085 ;
      RECT 8.885 -0.085 9.055 0.085 ;
      RECT 8.425 -0.085 8.595 0.085 ;
      RECT 7.965 -0.085 8.135 0.085 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.145 -0.085 0.315 0.085 ;
    LAYER via ;
      RECT 55.125 86.965 55.275 87.115 ;
      RECT 25.685 86.965 25.835 87.115 ;
      RECT 56.045 1.625 56.195 1.775 ;
      RECT 43.165 1.625 43.315 1.775 ;
      RECT 29.825 1.625 29.975 1.775 ;
      RECT 23.845 1.625 23.995 1.775 ;
      RECT 55.125 -0.075 55.275 0.075 ;
      RECT 25.685 -0.075 25.835 0.075 ;
    LAYER via2 ;
      RECT 55.1 86.94 55.3 87.14 ;
      RECT 25.66 86.94 25.86 87.14 ;
      RECT 64.76 67.9 64.96 68.1 ;
      RECT 1.74 66.54 1.94 66.74 ;
      RECT 64.76 63.82 64.96 64.02 ;
      RECT 1.28 61.78 1.48 61.98 ;
      RECT 1.74 23.02 1.94 23.22 ;
      RECT 64.76 15.54 64.96 15.74 ;
      RECT 1.74 13.5 1.94 13.7 ;
      RECT 55.1 -0.1 55.3 0.1 ;
      RECT 25.66 -0.1 25.86 0.1 ;
    LAYER via3 ;
      RECT 55.1 86.94 55.3 87.14 ;
      RECT 25.66 86.94 25.86 87.14 ;
      RECT 55.1 -0.1 55.3 0.1 ;
      RECT 25.66 -0.1 25.86 0.1 ;
    LAYER OVERLAP ;
      POLYGON 0 0 0 87.04 66.24 87.04 66.24 0 ;
  END
END cbx_1__0_

END LIBRARY
