VERSION 5.7 ;
BUSBITCHARS "[]" ;

UNITS
  DATABASE MICRONS 1000 ;
END UNITS

MANUFACTURINGGRID 0.005 ;

LAYER nwell
  TYPE MASTERSLICE ;
END nwell

LAYER pwell
  TYPE MASTERSLICE ;
END pwell

LAYER fieldpoly
  TYPE MASTERSLICE ;
END fieldpoly

LAYER li1
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.46 ;
  WIDTH 0.17 ;
END li1

LAYER mcon
  TYPE CUT ;
END mcon

LAYER met1
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.34 ;
  WIDTH 0.14 ;
END met1

LAYER via
  TYPE CUT ;
END via

LAYER met2
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.46 ;
  WIDTH 0.14 ;
END met2

LAYER via2
  TYPE CUT ;
END via2

LAYER met3
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.68 ;
  WIDTH 0.3 ;
END met3

LAYER via3
  TYPE CUT ;
END via3

LAYER met4
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.92 ;
  WIDTH 0.3 ;
END met4

LAYER via4
  TYPE CUT ;
END via4

LAYER met5
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 3.4 ;
  WIDTH 1.6 ;
END met5

LAYER diff
  TYPE MASTERSLICE ;
END diff

LAYER licon1
  TYPE MASTERSLICE ;
END licon1

LAYER OVERLAP
  TYPE OVERLAP ;
END OVERLAP

VIA L1M1_PR
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.145 -0.115 0.145 0.115 ;
END L1M1_PR

VIA L1M1_PR_R
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.115 -0.145 0.115 0.145 ;
END L1M1_PR_R

VIA L1M1_PR_M
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.115 -0.145 0.115 0.145 ;
END L1M1_PR_M

VIA L1M1_PR_MR
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.145 -0.115 0.145 0.115 ;
END L1M1_PR_MR

VIA L1M1_PR_C
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.145 -0.145 0.145 0.145 ;
END L1M1_PR_C

VIA M1M2_PR
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR

VIA M1M2_PR_Enc
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_Enc

VIA M1M2_PR_R
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_R

VIA M1M2_PR_R_Enc
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR_R_Enc

VIA M1M2_PR_M
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_M

VIA M1M2_PR_M_Enc
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR_M_Enc

VIA M1M2_PR_MR
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR_MR

VIA M1M2_PR_MR_Enc
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_MR_Enc

VIA M1M2_PR_C
  LAYER met1 ;
    RECT -0.16 -0.16 0.16 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.16 0.16 0.16 ;
END M1M2_PR_C

VIA M2M3_PR
  LAYER met2 ;
    RECT -0.14 -0.185 0.14 0.185 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR

VIA M2M3_PR_R
  LAYER met2 ;
    RECT -0.185 -0.14 0.185 0.14 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_R

VIA M2M3_PR_M
  LAYER met2 ;
    RECT -0.14 -0.185 0.14 0.185 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_M

VIA M2M3_PR_MR
  LAYER met2 ;
    RECT -0.185 -0.14 0.185 0.14 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_MR

VIA M2M3_PR_C
  LAYER met2 ;
    RECT -0.185 -0.185 0.185 0.185 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_C

VIA M3M4_PR
  LAYER met3 ;
    RECT -0.19 -0.16 0.19 0.16 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR

VIA M3M4_PR_R
  LAYER met3 ;
    RECT -0.16 -0.19 0.16 0.19 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_R

VIA M3M4_PR_M
  LAYER met3 ;
    RECT -0.19 -0.16 0.19 0.16 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_M

VIA M3M4_PR_MR
  LAYER met3 ;
    RECT -0.16 -0.19 0.16 0.19 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_MR

VIA M3M4_PR_C
  LAYER met3 ;
    RECT -0.19 -0.19 0.19 0.19 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_C

VIA M4M5_PR
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR

VIA M4M5_PR_R
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_R

VIA M4M5_PR_M
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_M

VIA M4M5_PR_MR
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_MR

VIA M4M5_PR_C
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_C

SITE unit
  CLASS CORE ;
  SYMMETRY Y ;
  SIZE 0.46 BY 2.72 ;
END unit

SITE unithddbl
  CLASS CORE ;
  SIZE 0.46 BY 5.44 ;
END unithddbl

MACRO sb_0__2_
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  SIZE 113.16 BY 103.36 ;
  SYMMETRY X Y ;
  PIN prog_clk[0]
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER met2 ;
        RECT 36.27 0 36.41 1.36 ;
    END
  END prog_clk[0]
  PIN chanx_right_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.78 86.89 113.16 87.19 ;
    END
  END chanx_right_in[0]
  PIN chanx_right_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.78 56.97 113.16 57.27 ;
    END
  END chanx_right_in[1]
  PIN chanx_right_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.78 99.13 113.16 99.43 ;
    END
  END chanx_right_in[2]
  PIN chanx_right_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.78 96.41 113.16 96.71 ;
    END
  END chanx_right_in[3]
  PIN chanx_right_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.78 33.85 113.16 34.15 ;
    END
  END chanx_right_in[4]
  PIN chanx_right_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.78 62.41 113.16 62.71 ;
    END
  END chanx_right_in[5]
  PIN chanx_right_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.78 31.13 113.16 31.43 ;
    END
  END chanx_right_in[6]
  PIN chanx_right_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.78 50.17 113.16 50.47 ;
    END
  END chanx_right_in[7]
  PIN chanx_right_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.78 77.37 113.16 77.67 ;
    END
  END chanx_right_in[8]
  PIN chanx_right_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.78 35.21 113.16 35.51 ;
    END
  END chanx_right_in[9]
  PIN chanx_right_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.78 80.09 113.16 80.39 ;
    END
  END chanx_right_in[10]
  PIN chanx_right_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.78 58.33 113.16 58.63 ;
    END
  END chanx_right_in[11]
  PIN chanx_right_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.78 74.65 113.16 74.95 ;
    END
  END chanx_right_in[12]
  PIN chanx_right_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.78 36.57 113.16 36.87 ;
    END
  END chanx_right_in[13]
  PIN chanx_right_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.78 43.37 113.16 43.67 ;
    END
  END chanx_right_in[14]
  PIN chanx_right_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.78 55.61 113.16 55.91 ;
    END
  END chanx_right_in[15]
  PIN chanx_right_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.78 40.65 113.16 40.95 ;
    END
  END chanx_right_in[16]
  PIN chanx_right_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.78 61.05 113.16 61.35 ;
    END
  END chanx_right_in[17]
  PIN chanx_right_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.78 39.29 113.16 39.59 ;
    END
  END chanx_right_in[18]
  PIN chanx_right_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.78 71.93 113.16 72.23 ;
    END
  END chanx_right_in[19]
  PIN right_top_grid_pin_1_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.87 102 110.01 103.36 ;
    END
  END right_top_grid_pin_1_[0]
  PIN chany_bottom_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.71 0 65.85 1.36 ;
    END
  END chany_bottom_in[0]
  PIN chany_bottom_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.65 0 14.79 1.36 ;
    END
  END chany_bottom_in[1]
  PIN chany_bottom_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.23 0 71.37 1.36 ;
    END
  END chany_bottom_in[2]
  PIN chany_bottom_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.73 0 13.87 1.36 ;
    END
  END chany_bottom_in[3]
  PIN chany_bottom_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.07 0 73.21 1.36 ;
    END
  END chany_bottom_in[4]
  PIN chany_bottom_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.15 0 49.29 1.36 ;
    END
  END chany_bottom_in[5]
  PIN chany_bottom_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.83 0 52.97 1.36 ;
    END
  END chany_bottom_in[6]
  PIN chany_bottom_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.01 0 22.15 1.36 ;
    END
  END chany_bottom_in[7]
  PIN chany_bottom_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.85 0 23.99 1.36 ;
    END
  END chany_bottom_in[8]
  PIN chany_bottom_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.93 0 23.07 1.36 ;
    END
  END chany_bottom_in[9]
  PIN chany_bottom_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.91 0 52.05 1.36 ;
    END
  END chany_bottom_in[10]
  PIN chany_bottom_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.75 0 30.89 1.36 ;
    END
  END chany_bottom_in[11]
  PIN chany_bottom_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.87 0 64.01 1.36 ;
    END
  END chany_bottom_in[12]
  PIN chany_bottom_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.15 0 72.29 1.36 ;
    END
  END chany_bottom_in[13]
  PIN chany_bottom_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.63 0 43.77 1.36 ;
    END
  END chany_bottom_in[14]
  PIN chany_bottom_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.39 0 46.53 1.36 ;
    END
  END chany_bottom_in[15]
  PIN chany_bottom_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.79 0 41.93 1.36 ;
    END
  END chany_bottom_in[16]
  PIN chany_bottom_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.83 0 29.97 1.36 ;
    END
  END chany_bottom_in[17]
  PIN chany_bottom_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.61 0 26.75 1.36 ;
    END
  END chany_bottom_in[18]
  PIN chany_bottom_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.77 0 24.91 1.36 ;
    END
  END chany_bottom_in[19]
  PIN bottom_left_grid_pin_1_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.23 0 2.37 1.36 ;
    END
  END bottom_left_grid_pin_1_[0]
  PIN ccff_head[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.79 102 110.93 103.36 ;
    END
  END ccff_head[0]
  PIN chanx_right_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.78 73.29 113.16 73.59 ;
    END
  END chanx_right_out[0]
  PIN chanx_right_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.78 47.45 113.16 47.75 ;
    END
  END chanx_right_out[1]
  PIN chanx_right_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.78 52.89 113.16 53.19 ;
    END
  END chanx_right_out[2]
  PIN chanx_right_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.78 82.81 113.16 83.11 ;
    END
  END chanx_right_out[3]
  PIN chanx_right_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.78 78.73 113.16 79.03 ;
    END
  END chanx_right_out[4]
  PIN chanx_right_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.78 95.05 113.16 95.35 ;
    END
  END chanx_right_out[5]
  PIN chanx_right_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.78 84.17 113.16 84.47 ;
    END
  END chanx_right_out[6]
  PIN chanx_right_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.78 93.69 113.16 93.99 ;
    END
  END chanx_right_out[7]
  PIN chanx_right_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.78 85.53 113.16 85.83 ;
    END
  END chanx_right_out[8]
  PIN chanx_right_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.78 44.73 113.16 45.03 ;
    END
  END chanx_right_out[9]
  PIN chanx_right_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.78 51.53 113.16 51.83 ;
    END
  END chanx_right_out[10]
  PIN chanx_right_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.78 69.21 113.16 69.51 ;
    END
  END chanx_right_out[11]
  PIN chanx_right_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.78 42.01 113.16 42.31 ;
    END
  END chanx_right_out[12]
  PIN chanx_right_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.78 66.49 113.16 66.79 ;
    END
  END chanx_right_out[13]
  PIN chanx_right_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.78 90.97 113.16 91.27 ;
    END
  END chanx_right_out[14]
  PIN chanx_right_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.78 67.85 113.16 68.15 ;
    END
  END chanx_right_out[15]
  PIN chanx_right_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.78 63.77 113.16 64.07 ;
    END
  END chanx_right_out[16]
  PIN chanx_right_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.78 88.25 113.16 88.55 ;
    END
  END chanx_right_out[17]
  PIN chanx_right_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.78 89.61 113.16 89.91 ;
    END
  END chanx_right_out[18]
  PIN chanx_right_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.78 46.09 113.16 46.39 ;
    END
  END chanx_right_out[19]
  PIN chany_bottom_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.07 0 50.21 1.36 ;
    END
  END chany_bottom_out[0]
  PIN chany_bottom_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.43 0 34.57 1.36 ;
    END
  END chany_bottom_out[1]
  PIN chany_bottom_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.63 0 66.77 1.36 ;
    END
  END chany_bottom_out[2]
  PIN chany_bottom_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.55 0 44.69 1.36 ;
    END
  END chany_bottom_out[3]
  PIN chany_bottom_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.99 0 51.13 1.36 ;
    END
  END chany_bottom_out[4]
  PIN chany_bottom_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.47 0 45.61 1.36 ;
    END
  END chany_bottom_out[5]
  PIN chany_bottom_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.31 0 70.45 1.36 ;
    END
  END chany_bottom_out[6]
  PIN chany_bottom_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.47 0 68.61 1.36 ;
    END
  END chany_bottom_out[7]
  PIN chany_bottom_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.39 0 69.53 1.36 ;
    END
  END chany_bottom_out[8]
  PIN chany_bottom_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.69 0 25.83 1.36 ;
    END
  END chany_bottom_out[9]
  PIN chany_bottom_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.71 0 42.85 1.36 ;
    END
  END chany_bottom_out[10]
  PIN chany_bottom_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.23 0 48.37 1.36 ;
    END
  END chany_bottom_out[11]
  PIN chany_bottom_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.55 0 67.69 1.36 ;
    END
  END chany_bottom_out[12]
  PIN chany_bottom_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 49.53 0 49.83 1.36 ;
    END
  END chany_bottom_out[13]
  PIN chany_bottom_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 45.85 0 46.15 1.36 ;
    END
  END chany_bottom_out[14]
  PIN chany_bottom_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 47.69 0 47.99 1.36 ;
    END
  END chany_bottom_out[15]
  PIN chany_bottom_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.45 0 28.59 1.36 ;
    END
  END chany_bottom_out[16]
  PIN chany_bottom_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.31 0 47.45 1.36 ;
    END
  END chany_bottom_out[17]
  PIN chany_bottom_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 23.77 0 24.07 1.36 ;
    END
  END chany_bottom_out[18]
  PIN chany_bottom_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 25.61 0 25.91 1.36 ;
    END
  END chany_bottom_out[19]
  PIN ccff_tail[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.21 0 54.35 1.36 ;
    END
  END ccff_tail[0]
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 0.48 2.96 ;
        RECT 84.16 2.48 84.64 2.96 ;
        RECT 0 7.92 0.48 8.4 ;
        RECT 84.16 7.92 84.64 8.4 ;
        RECT 0 13.36 0.48 13.84 ;
        RECT 84.16 13.36 84.64 13.84 ;
        RECT 0 18.8 0.48 19.28 ;
        RECT 84.16 18.8 84.64 19.28 ;
        RECT 0 24.24 0.48 24.72 ;
        RECT 84.16 24.24 84.64 24.72 ;
        RECT 0 29.68 0.48 30.16 ;
        RECT 112.68 29.68 113.16 30.16 ;
        RECT 0 35.12 0.48 35.6 ;
        RECT 112.68 35.12 113.16 35.6 ;
        RECT 0 40.56 0.48 41.04 ;
        RECT 112.68 40.56 113.16 41.04 ;
        RECT 0 46 0.48 46.48 ;
        RECT 112.68 46 113.16 46.48 ;
        RECT 0 51.44 0.48 51.92 ;
        RECT 112.68 51.44 113.16 51.92 ;
        RECT 0 56.88 0.48 57.36 ;
        RECT 112.68 56.88 113.16 57.36 ;
        RECT 0 62.32 0.48 62.8 ;
        RECT 112.68 62.32 113.16 62.8 ;
        RECT 0 67.76 0.48 68.24 ;
        RECT 112.68 67.76 113.16 68.24 ;
        RECT 0 73.2 0.48 73.68 ;
        RECT 112.68 73.2 113.16 73.68 ;
        RECT 0 78.64 0.48 79.12 ;
        RECT 112.68 78.64 113.16 79.12 ;
        RECT 0 84.08 0.48 84.56 ;
        RECT 112.68 84.08 113.16 84.56 ;
        RECT 0 89.52 0.48 90 ;
        RECT 112.68 89.52 113.16 90 ;
        RECT 0 94.96 0.48 95.44 ;
        RECT 112.68 94.96 113.16 95.44 ;
        RECT 0 100.4 0.48 100.88 ;
        RECT 112.68 100.4 113.16 100.88 ;
      LAYER met4 ;
        RECT 12.58 0 13.18 0.6 ;
        RECT 42.02 0 42.62 0.6 ;
        RECT 71.46 0 72.06 0.6 ;
        RECT 106.42 27.2 107.02 27.8 ;
        RECT 12.58 102.76 13.18 103.36 ;
        RECT 42.02 102.76 42.62 103.36 ;
        RECT 71.46 102.76 72.06 103.36 ;
        RECT 106.42 102.76 107.02 103.36 ;
      LAYER met5 ;
        RECT 0 43.28 3.2 46.48 ;
        RECT 109.96 43.28 113.16 46.48 ;
        RECT 0 84.08 3.2 87.28 ;
        RECT 109.96 84.08 113.16 87.28 ;
    END
  END VDD
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 0 84.64 0.24 ;
        RECT 0 5.2 0.48 5.68 ;
        RECT 84.16 5.2 84.64 5.68 ;
        RECT 0 10.64 0.48 11.12 ;
        RECT 84.16 10.64 84.64 11.12 ;
        RECT 0 16.08 0.48 16.56 ;
        RECT 84.16 16.08 84.64 16.56 ;
        RECT 0 21.52 0.48 22 ;
        RECT 84.16 21.52 84.64 22 ;
        RECT 0 26.96 113.16 27.44 ;
        RECT 0 32.4 0.48 32.88 ;
        RECT 112.68 32.4 113.16 32.88 ;
        RECT 0 37.84 0.48 38.32 ;
        RECT 112.68 37.84 113.16 38.32 ;
        RECT 0 43.28 0.48 43.76 ;
        RECT 112.68 43.28 113.16 43.76 ;
        RECT 0 48.72 0.48 49.2 ;
        RECT 112.68 48.72 113.16 49.2 ;
        RECT 0 54.16 0.48 54.64 ;
        RECT 112.68 54.16 113.16 54.64 ;
        RECT 0 59.6 0.48 60.08 ;
        RECT 112.68 59.6 113.16 60.08 ;
        RECT 0 65.04 0.48 65.52 ;
        RECT 112.68 65.04 113.16 65.52 ;
        RECT 0 70.48 0.48 70.96 ;
        RECT 112.68 70.48 113.16 70.96 ;
        RECT 0 75.92 0.48 76.4 ;
        RECT 112.68 75.92 113.16 76.4 ;
        RECT 0 81.36 0.48 81.84 ;
        RECT 112.68 81.36 113.16 81.84 ;
        RECT 0 86.8 0.48 87.28 ;
        RECT 112.68 86.8 113.16 87.28 ;
        RECT 0 92.24 0.48 92.72 ;
        RECT 112.68 92.24 113.16 92.72 ;
        RECT 0 97.68 0.48 98.16 ;
        RECT 112.68 97.68 113.16 98.16 ;
        RECT 0 103.12 113.16 103.36 ;
      LAYER met5 ;
        RECT 0 4.52 3.2 7.72 ;
        RECT 81.44 4.52 84.64 7.72 ;
        RECT 0 63.68 3.2 66.88 ;
        RECT 109.96 63.68 113.16 66.88 ;
      LAYER met4 ;
        RECT 27.3 0 27.9 0.6 ;
        RECT 56.74 0 57.34 0.6 ;
        RECT 27.3 102.76 27.9 103.36 ;
        RECT 56.74 102.76 57.34 103.36 ;
    END
  END VSS
  OBS
    LAYER li1 ;
      RECT 0 103.275 113.16 103.445 ;
      RECT 112.24 100.555 113.16 100.725 ;
      RECT 0 100.555 3.68 100.725 ;
      RECT 112.24 97.835 113.16 98.005 ;
      RECT 0 97.835 3.68 98.005 ;
      RECT 112.24 95.115 113.16 95.285 ;
      RECT 0 95.115 3.68 95.285 ;
      RECT 112.24 92.395 113.16 92.565 ;
      RECT 0 92.395 3.68 92.565 ;
      RECT 112.24 89.675 113.16 89.845 ;
      RECT 0 89.675 3.68 89.845 ;
      RECT 112.24 86.955 113.16 87.125 ;
      RECT 0 86.955 3.68 87.125 ;
      RECT 112.24 84.235 113.16 84.405 ;
      RECT 0 84.235 3.68 84.405 ;
      RECT 112.24 81.515 113.16 81.685 ;
      RECT 0 81.515 3.68 81.685 ;
      RECT 112.24 78.795 113.16 78.965 ;
      RECT 0 78.795 3.68 78.965 ;
      RECT 112.24 76.075 113.16 76.245 ;
      RECT 0 76.075 3.68 76.245 ;
      RECT 112.24 73.355 113.16 73.525 ;
      RECT 0 73.355 3.68 73.525 ;
      RECT 112.24 70.635 113.16 70.805 ;
      RECT 0 70.635 3.68 70.805 ;
      RECT 112.24 67.915 113.16 68.085 ;
      RECT 0 67.915 3.68 68.085 ;
      RECT 112.24 65.195 113.16 65.365 ;
      RECT 0 65.195 3.68 65.365 ;
      RECT 112.24 62.475 113.16 62.645 ;
      RECT 0 62.475 3.68 62.645 ;
      RECT 112.24 59.755 113.16 59.925 ;
      RECT 0 59.755 3.68 59.925 ;
      RECT 112.24 57.035 113.16 57.205 ;
      RECT 0 57.035 3.68 57.205 ;
      RECT 112.24 54.315 113.16 54.485 ;
      RECT 0 54.315 3.68 54.485 ;
      RECT 112.24 51.595 113.16 51.765 ;
      RECT 0 51.595 3.68 51.765 ;
      RECT 112.24 48.875 113.16 49.045 ;
      RECT 0 48.875 3.68 49.045 ;
      RECT 112.24 46.155 113.16 46.325 ;
      RECT 0 46.155 3.68 46.325 ;
      RECT 112.24 43.435 113.16 43.605 ;
      RECT 0 43.435 3.68 43.605 ;
      RECT 112.24 40.715 113.16 40.885 ;
      RECT 0 40.715 3.68 40.885 ;
      RECT 112.7 37.995 113.16 38.165 ;
      RECT 0 37.995 3.68 38.165 ;
      RECT 112.7 35.275 113.16 35.445 ;
      RECT 0 35.275 3.68 35.445 ;
      RECT 112.24 32.555 113.16 32.725 ;
      RECT 0 32.555 3.68 32.725 ;
      RECT 112.24 29.835 113.16 30.005 ;
      RECT 0 29.835 3.68 30.005 ;
      RECT 80.96 27.115 113.16 27.285 ;
      RECT 0 27.115 3.68 27.285 ;
      RECT 83.72 24.395 84.64 24.565 ;
      RECT 0 24.395 3.68 24.565 ;
      RECT 83.72 21.675 84.64 21.845 ;
      RECT 0 21.675 3.68 21.845 ;
      RECT 83.72 18.955 84.64 19.125 ;
      RECT 0 18.955 3.68 19.125 ;
      RECT 84.18 16.235 84.64 16.405 ;
      RECT 0 16.235 3.68 16.405 ;
      RECT 80.96 13.515 84.64 13.685 ;
      RECT 0 13.515 3.68 13.685 ;
      RECT 80.96 10.795 84.64 10.965 ;
      RECT 0 10.795 3.68 10.965 ;
      RECT 83.72 8.075 84.64 8.245 ;
      RECT 0 8.075 3.68 8.245 ;
      RECT 83.72 5.355 84.64 5.525 ;
      RECT 0 5.355 3.68 5.525 ;
      RECT 80.96 2.635 84.64 2.805 ;
      RECT 0 2.635 3.68 2.805 ;
      RECT 0 -0.085 84.64 0.085 ;
    LAYER met2 ;
      RECT 56.9 103.175 57.18 103.545 ;
      RECT 27.46 103.175 27.74 103.545 ;
      RECT 56.9 -0.185 57.18 0.185 ;
      RECT 27.46 -0.185 27.74 0.185 ;
      POLYGON 112.88 103.08 112.88 27.48 84.36 27.48 84.36 0.28 73.49 0.28 73.49 1.64 72.79 1.64 72.79 0.28 72.57 0.28 72.57 1.64 71.87 1.64 71.87 0.28 71.65 0.28 71.65 1.64 70.95 1.64 70.95 0.28 70.73 0.28 70.73 1.64 70.03 1.64 70.03 0.28 69.81 0.28 69.81 1.64 69.11 1.64 69.11 0.28 68.89 0.28 68.89 1.64 68.19 1.64 68.19 0.28 67.97 0.28 67.97 1.64 67.27 1.64 67.27 0.28 67.05 0.28 67.05 1.64 66.35 1.64 66.35 0.28 66.13 0.28 66.13 1.64 65.43 1.64 65.43 0.28 64.29 0.28 64.29 1.64 63.59 1.64 63.59 0.28 54.63 0.28 54.63 1.64 53.93 1.64 53.93 0.28 53.25 0.28 53.25 1.64 52.55 1.64 52.55 0.28 52.33 0.28 52.33 1.64 51.63 1.64 51.63 0.28 51.41 0.28 51.41 1.64 50.71 1.64 50.71 0.28 50.49 0.28 50.49 1.64 49.79 1.64 49.79 0.28 49.57 0.28 49.57 1.64 48.87 1.64 48.87 0.28 48.65 0.28 48.65 1.64 47.95 1.64 47.95 0.28 47.73 0.28 47.73 1.64 47.03 1.64 47.03 0.28 46.81 0.28 46.81 1.64 46.11 1.64 46.11 0.28 45.89 0.28 45.89 1.64 45.19 1.64 45.19 0.28 44.97 0.28 44.97 1.64 44.27 1.64 44.27 0.28 44.05 0.28 44.05 1.64 43.35 1.64 43.35 0.28 43.13 0.28 43.13 1.64 42.43 1.64 42.43 0.28 42.21 0.28 42.21 1.64 41.51 1.64 41.51 0.28 36.69 0.28 36.69 1.64 35.99 1.64 35.99 0.28 34.85 0.28 34.85 1.64 34.15 1.64 34.15 0.28 31.17 0.28 31.17 1.64 30.47 1.64 30.47 0.28 30.25 0.28 30.25 1.64 29.55 1.64 29.55 0.28 28.87 0.28 28.87 1.64 28.17 1.64 28.17 0.28 27.03 0.28 27.03 1.64 26.33 1.64 26.33 0.28 26.11 0.28 26.11 1.64 25.41 1.64 25.41 0.28 25.19 0.28 25.19 1.64 24.49 1.64 24.49 0.28 24.27 0.28 24.27 1.64 23.57 1.64 23.57 0.28 23.35 0.28 23.35 1.64 22.65 1.64 22.65 0.28 22.43 0.28 22.43 1.64 21.73 1.64 21.73 0.28 15.07 0.28 15.07 1.64 14.37 1.64 14.37 0.28 14.15 0.28 14.15 1.64 13.45 1.64 13.45 0.28 2.65 0.28 2.65 1.64 1.95 1.64 1.95 0.28 0.28 0.28 0.28 103.08 109.59 103.08 109.59 101.72 110.29 101.72 110.29 103.08 110.51 103.08 110.51 101.72 111.21 101.72 111.21 103.08 ;
    LAYER met3 ;
      POLYGON 57.205 103.525 57.205 103.52 57.42 103.52 57.42 103.2 57.205 103.2 57.205 103.195 56.875 103.195 56.875 103.2 56.66 103.2 56.66 103.52 56.875 103.52 56.875 103.525 ;
      POLYGON 27.765 103.525 27.765 103.52 27.98 103.52 27.98 103.2 27.765 103.2 27.765 103.195 27.435 103.195 27.435 103.2 27.22 103.2 27.22 103.52 27.435 103.52 27.435 103.525 ;
      POLYGON 57.205 0.165 57.205 0.16 57.42 0.16 57.42 -0.16 57.205 -0.16 57.205 -0.165 56.875 -0.165 56.875 -0.16 56.66 -0.16 56.66 0.16 56.875 0.16 56.875 0.165 ;
      POLYGON 27.765 0.165 27.765 0.16 27.98 0.16 27.98 -0.16 27.765 -0.16 27.765 -0.165 27.435 -0.165 27.435 -0.16 27.22 -0.16 27.22 0.16 27.435 0.16 27.435 0.165 ;
      POLYGON 112.76 102.96 112.76 99.83 111.38 99.83 111.38 98.73 112.76 98.73 112.76 97.11 111.38 97.11 111.38 96.01 112.76 96.01 112.76 95.75 111.38 95.75 111.38 94.65 112.76 94.65 112.76 94.39 111.38 94.39 111.38 93.29 112.76 93.29 112.76 91.67 111.38 91.67 111.38 90.57 112.76 90.57 112.76 90.31 111.38 90.31 111.38 89.21 112.76 89.21 112.76 88.95 111.38 88.95 111.38 87.85 112.76 87.85 112.76 87.59 111.38 87.59 111.38 86.49 112.76 86.49 112.76 86.23 111.38 86.23 111.38 85.13 112.76 85.13 112.76 84.87 111.38 84.87 111.38 83.77 112.76 83.77 112.76 83.51 111.38 83.51 111.38 82.41 112.76 82.41 112.76 80.79 111.38 80.79 111.38 79.69 112.76 79.69 112.76 79.43 111.38 79.43 111.38 78.33 112.76 78.33 112.76 78.07 111.38 78.07 111.38 76.97 112.76 76.97 112.76 75.35 111.38 75.35 111.38 74.25 112.76 74.25 112.76 73.99 111.38 73.99 111.38 72.89 112.76 72.89 112.76 72.63 111.38 72.63 111.38 71.53 112.76 71.53 112.76 69.91 111.38 69.91 111.38 68.81 112.76 68.81 112.76 68.55 111.38 68.55 111.38 67.45 112.76 67.45 112.76 67.19 111.38 67.19 111.38 66.09 112.76 66.09 112.76 64.47 111.38 64.47 111.38 63.37 112.76 63.37 112.76 63.11 111.38 63.11 111.38 62.01 112.76 62.01 112.76 61.75 111.38 61.75 111.38 60.65 112.76 60.65 112.76 59.03 111.38 59.03 111.38 57.93 112.76 57.93 112.76 57.67 111.38 57.67 111.38 56.57 112.76 56.57 112.76 56.31 111.38 56.31 111.38 55.21 112.76 55.21 112.76 53.59 111.38 53.59 111.38 52.49 112.76 52.49 112.76 52.23 111.38 52.23 111.38 51.13 112.76 51.13 112.76 50.87 111.38 50.87 111.38 49.77 112.76 49.77 112.76 48.15 111.38 48.15 111.38 47.05 112.76 47.05 112.76 46.79 111.38 46.79 111.38 45.69 112.76 45.69 112.76 45.43 111.38 45.43 111.38 44.33 112.76 44.33 112.76 44.07 111.38 44.07 111.38 42.97 112.76 42.97 112.76 42.71 111.38 42.71 111.38 41.61 112.76 41.61 112.76 41.35 111.38 41.35 111.38 40.25 112.76 40.25 112.76 39.99 111.38 39.99 111.38 38.89 112.76 38.89 112.76 37.27 111.38 37.27 111.38 36.17 112.76 36.17 112.76 35.91 111.38 35.91 111.38 34.81 112.76 34.81 112.76 34.55 111.38 34.55 111.38 33.45 112.76 33.45 112.76 31.83 111.38 31.83 111.38 30.73 112.76 30.73 112.76 27.6 84.24 27.6 84.24 0.4 0.4 0.4 0.4 102.96 ;
    LAYER met4 ;
      POLYGON 112.76 102.96 112.76 27.6 107.42 27.6 107.42 28.2 106.02 28.2 106.02 27.6 84.24 27.6 84.24 0.4 72.46 0.4 72.46 1 71.06 1 71.06 0.4 57.74 0.4 57.74 1 56.34 1 56.34 0.4 50.23 0.4 50.23 1.76 49.13 1.76 49.13 0.4 48.39 0.4 48.39 1.76 47.29 1.76 47.29 0.4 46.55 0.4 46.55 1.76 45.45 1.76 45.45 0.4 43.02 0.4 43.02 1 41.62 1 41.62 0.4 28.3 0.4 28.3 1 26.9 1 26.9 0.4 26.31 0.4 26.31 1.76 25.21 1.76 25.21 0.4 24.47 0.4 24.47 1.76 23.37 1.76 23.37 0.4 13.58 0.4 13.58 1 12.18 1 12.18 0.4 0.4 0.4 0.4 102.96 12.18 102.96 12.18 102.36 13.58 102.36 13.58 102.96 26.9 102.96 26.9 102.36 28.3 102.36 28.3 102.96 41.62 102.96 41.62 102.36 43.02 102.36 43.02 102.96 56.34 102.96 56.34 102.36 57.74 102.36 57.74 102.96 71.06 102.96 71.06 102.36 72.46 102.36 72.46 102.96 106.02 102.96 106.02 102.36 107.42 102.36 107.42 102.96 ;
    LAYER met5 ;
      POLYGON 109.96 100.16 109.96 90.48 106.76 90.48 106.76 80.88 109.96 80.88 109.96 70.08 106.76 70.08 106.76 60.48 109.96 60.48 109.96 49.68 106.76 49.68 106.76 40.08 109.96 40.08 109.96 30.4 81.44 30.4 81.44 10.92 78.24 10.92 78.24 3.2 6.4 3.2 6.4 10.92 3.2 10.92 3.2 40.08 6.4 40.08 6.4 49.68 3.2 49.68 3.2 60.48 6.4 60.48 6.4 70.08 3.2 70.08 3.2 80.88 6.4 80.88 6.4 90.48 3.2 90.48 3.2 100.16 ;
    LAYER met1 ;
      POLYGON 112.88 102.84 112.88 101.16 112.4 101.16 112.4 100.12 112.88 100.12 112.88 98.44 112.4 98.44 112.4 97.4 112.88 97.4 112.88 95.72 112.4 95.72 112.4 94.68 112.88 94.68 112.88 93 112.4 93 112.4 91.96 112.88 91.96 112.88 90.28 112.4 90.28 112.4 89.24 112.88 89.24 112.88 87.56 112.4 87.56 112.4 86.52 112.88 86.52 112.88 84.84 112.4 84.84 112.4 83.8 112.88 83.8 112.88 82.12 112.4 82.12 112.4 81.08 112.88 81.08 112.88 79.4 112.4 79.4 112.4 78.36 112.88 78.36 112.88 76.68 112.4 76.68 112.4 75.64 112.88 75.64 112.88 73.96 112.4 73.96 112.4 72.92 112.88 72.92 112.88 71.24 112.4 71.24 112.4 70.2 112.88 70.2 112.88 68.52 112.4 68.52 112.4 67.48 112.88 67.48 112.88 65.8 112.4 65.8 112.4 64.76 112.88 64.76 112.88 63.08 112.4 63.08 112.4 62.04 112.88 62.04 112.88 60.36 112.4 60.36 112.4 59.32 112.88 59.32 112.88 57.64 112.4 57.64 112.4 56.6 112.88 56.6 112.88 54.92 112.4 54.92 112.4 53.88 112.88 53.88 112.88 52.2 112.4 52.2 112.4 51.16 112.88 51.16 112.88 49.48 112.4 49.48 112.4 48.44 112.88 48.44 112.88 46.76 112.4 46.76 112.4 45.72 112.88 45.72 112.88 44.04 112.4 44.04 112.4 43 112.88 43 112.88 41.32 112.4 41.32 112.4 40.28 112.88 40.28 112.88 38.6 112.4 38.6 112.4 37.56 112.88 37.56 112.88 35.88 112.4 35.88 112.4 34.84 112.88 34.84 112.88 33.16 112.4 33.16 112.4 32.12 112.88 32.12 112.88 30.44 112.4 30.44 112.4 29.4 112.88 29.4 112.88 27.72 0.28 27.72 0.28 29.4 0.76 29.4 0.76 30.44 0.28 30.44 0.28 32.12 0.76 32.12 0.76 33.16 0.28 33.16 0.28 34.84 0.76 34.84 0.76 35.88 0.28 35.88 0.28 37.56 0.76 37.56 0.76 38.6 0.28 38.6 0.28 40.28 0.76 40.28 0.76 41.32 0.28 41.32 0.28 43 0.76 43 0.76 44.04 0.28 44.04 0.28 45.72 0.76 45.72 0.76 46.76 0.28 46.76 0.28 48.44 0.76 48.44 0.76 49.48 0.28 49.48 0.28 51.16 0.76 51.16 0.76 52.2 0.28 52.2 0.28 53.88 0.76 53.88 0.76 54.92 0.28 54.92 0.28 56.6 0.76 56.6 0.76 57.64 0.28 57.64 0.28 59.32 0.76 59.32 0.76 60.36 0.28 60.36 0.28 62.04 0.76 62.04 0.76 63.08 0.28 63.08 0.28 64.76 0.76 64.76 0.76 65.8 0.28 65.8 0.28 67.48 0.76 67.48 0.76 68.52 0.28 68.52 0.28 70.2 0.76 70.2 0.76 71.24 0.28 71.24 0.28 72.92 0.76 72.92 0.76 73.96 0.28 73.96 0.28 75.64 0.76 75.64 0.76 76.68 0.28 76.68 0.28 78.36 0.76 78.36 0.76 79.4 0.28 79.4 0.28 81.08 0.76 81.08 0.76 82.12 0.28 82.12 0.28 83.8 0.76 83.8 0.76 84.84 0.28 84.84 0.28 86.52 0.76 86.52 0.76 87.56 0.28 87.56 0.28 89.24 0.76 89.24 0.76 90.28 0.28 90.28 0.28 91.96 0.76 91.96 0.76 93 0.28 93 0.28 94.68 0.76 94.68 0.76 95.72 0.28 95.72 0.28 97.4 0.76 97.4 0.76 98.44 0.28 98.44 0.28 100.12 0.76 100.12 0.76 101.16 0.28 101.16 0.28 102.84 ;
      POLYGON 84.36 26.68 84.36 25 83.88 25 83.88 23.96 84.36 23.96 84.36 22.28 83.88 22.28 83.88 21.24 84.36 21.24 84.36 19.56 83.88 19.56 83.88 18.52 84.36 18.52 84.36 16.84 83.88 16.84 83.88 15.8 84.36 15.8 84.36 14.12 83.88 14.12 83.88 13.08 84.36 13.08 84.36 11.4 83.88 11.4 83.88 10.36 84.36 10.36 84.36 8.68 83.88 8.68 83.88 7.64 84.36 7.64 84.36 5.96 83.88 5.96 83.88 4.92 84.36 4.92 84.36 3.24 83.88 3.24 83.88 2.2 84.36 2.2 84.36 0.52 0.28 0.52 0.28 2.2 0.76 2.2 0.76 3.24 0.28 3.24 0.28 4.92 0.76 4.92 0.76 5.96 0.28 5.96 0.28 7.64 0.76 7.64 0.76 8.68 0.28 8.68 0.28 10.36 0.76 10.36 0.76 11.4 0.28 11.4 0.28 13.08 0.76 13.08 0.76 14.12 0.28 14.12 0.28 15.8 0.76 15.8 0.76 16.84 0.28 16.84 0.28 18.52 0.76 18.52 0.76 19.56 0.28 19.56 0.28 21.24 0.76 21.24 0.76 22.28 0.28 22.28 0.28 23.96 0.76 23.96 0.76 25 0.28 25 0.28 26.68 ;
    LAYER li1 ;
      POLYGON 112.82 103.02 112.82 27.54 84.3 27.54 84.3 0.34 0.34 0.34 0.34 103.02 ;
    LAYER mcon ;
      RECT 112.845 103.275 113.015 103.445 ;
      RECT 112.385 103.275 112.555 103.445 ;
      RECT 111.925 103.275 112.095 103.445 ;
      RECT 111.465 103.275 111.635 103.445 ;
      RECT 111.005 103.275 111.175 103.445 ;
      RECT 110.545 103.275 110.715 103.445 ;
      RECT 110.085 103.275 110.255 103.445 ;
      RECT 109.625 103.275 109.795 103.445 ;
      RECT 109.165 103.275 109.335 103.445 ;
      RECT 108.705 103.275 108.875 103.445 ;
      RECT 108.245 103.275 108.415 103.445 ;
      RECT 107.785 103.275 107.955 103.445 ;
      RECT 107.325 103.275 107.495 103.445 ;
      RECT 106.865 103.275 107.035 103.445 ;
      RECT 106.405 103.275 106.575 103.445 ;
      RECT 105.945 103.275 106.115 103.445 ;
      RECT 105.485 103.275 105.655 103.445 ;
      RECT 105.025 103.275 105.195 103.445 ;
      RECT 104.565 103.275 104.735 103.445 ;
      RECT 104.105 103.275 104.275 103.445 ;
      RECT 103.645 103.275 103.815 103.445 ;
      RECT 103.185 103.275 103.355 103.445 ;
      RECT 102.725 103.275 102.895 103.445 ;
      RECT 102.265 103.275 102.435 103.445 ;
      RECT 101.805 103.275 101.975 103.445 ;
      RECT 101.345 103.275 101.515 103.445 ;
      RECT 100.885 103.275 101.055 103.445 ;
      RECT 100.425 103.275 100.595 103.445 ;
      RECT 99.965 103.275 100.135 103.445 ;
      RECT 99.505 103.275 99.675 103.445 ;
      RECT 99.045 103.275 99.215 103.445 ;
      RECT 98.585 103.275 98.755 103.445 ;
      RECT 98.125 103.275 98.295 103.445 ;
      RECT 97.665 103.275 97.835 103.445 ;
      RECT 97.205 103.275 97.375 103.445 ;
      RECT 96.745 103.275 96.915 103.445 ;
      RECT 96.285 103.275 96.455 103.445 ;
      RECT 95.825 103.275 95.995 103.445 ;
      RECT 95.365 103.275 95.535 103.445 ;
      RECT 94.905 103.275 95.075 103.445 ;
      RECT 94.445 103.275 94.615 103.445 ;
      RECT 93.985 103.275 94.155 103.445 ;
      RECT 93.525 103.275 93.695 103.445 ;
      RECT 93.065 103.275 93.235 103.445 ;
      RECT 92.605 103.275 92.775 103.445 ;
      RECT 92.145 103.275 92.315 103.445 ;
      RECT 91.685 103.275 91.855 103.445 ;
      RECT 91.225 103.275 91.395 103.445 ;
      RECT 90.765 103.275 90.935 103.445 ;
      RECT 90.305 103.275 90.475 103.445 ;
      RECT 89.845 103.275 90.015 103.445 ;
      RECT 89.385 103.275 89.555 103.445 ;
      RECT 88.925 103.275 89.095 103.445 ;
      RECT 88.465 103.275 88.635 103.445 ;
      RECT 88.005 103.275 88.175 103.445 ;
      RECT 87.545 103.275 87.715 103.445 ;
      RECT 87.085 103.275 87.255 103.445 ;
      RECT 86.625 103.275 86.795 103.445 ;
      RECT 86.165 103.275 86.335 103.445 ;
      RECT 85.705 103.275 85.875 103.445 ;
      RECT 85.245 103.275 85.415 103.445 ;
      RECT 84.785 103.275 84.955 103.445 ;
      RECT 84.325 103.275 84.495 103.445 ;
      RECT 83.865 103.275 84.035 103.445 ;
      RECT 83.405 103.275 83.575 103.445 ;
      RECT 82.945 103.275 83.115 103.445 ;
      RECT 82.485 103.275 82.655 103.445 ;
      RECT 82.025 103.275 82.195 103.445 ;
      RECT 81.565 103.275 81.735 103.445 ;
      RECT 81.105 103.275 81.275 103.445 ;
      RECT 80.645 103.275 80.815 103.445 ;
      RECT 80.185 103.275 80.355 103.445 ;
      RECT 79.725 103.275 79.895 103.445 ;
      RECT 79.265 103.275 79.435 103.445 ;
      RECT 78.805 103.275 78.975 103.445 ;
      RECT 78.345 103.275 78.515 103.445 ;
      RECT 77.885 103.275 78.055 103.445 ;
      RECT 77.425 103.275 77.595 103.445 ;
      RECT 76.965 103.275 77.135 103.445 ;
      RECT 76.505 103.275 76.675 103.445 ;
      RECT 76.045 103.275 76.215 103.445 ;
      RECT 75.585 103.275 75.755 103.445 ;
      RECT 75.125 103.275 75.295 103.445 ;
      RECT 74.665 103.275 74.835 103.445 ;
      RECT 74.205 103.275 74.375 103.445 ;
      RECT 73.745 103.275 73.915 103.445 ;
      RECT 73.285 103.275 73.455 103.445 ;
      RECT 72.825 103.275 72.995 103.445 ;
      RECT 72.365 103.275 72.535 103.445 ;
      RECT 71.905 103.275 72.075 103.445 ;
      RECT 71.445 103.275 71.615 103.445 ;
      RECT 70.985 103.275 71.155 103.445 ;
      RECT 70.525 103.275 70.695 103.445 ;
      RECT 70.065 103.275 70.235 103.445 ;
      RECT 69.605 103.275 69.775 103.445 ;
      RECT 69.145 103.275 69.315 103.445 ;
      RECT 68.685 103.275 68.855 103.445 ;
      RECT 68.225 103.275 68.395 103.445 ;
      RECT 67.765 103.275 67.935 103.445 ;
      RECT 67.305 103.275 67.475 103.445 ;
      RECT 66.845 103.275 67.015 103.445 ;
      RECT 66.385 103.275 66.555 103.445 ;
      RECT 65.925 103.275 66.095 103.445 ;
      RECT 65.465 103.275 65.635 103.445 ;
      RECT 65.005 103.275 65.175 103.445 ;
      RECT 64.545 103.275 64.715 103.445 ;
      RECT 64.085 103.275 64.255 103.445 ;
      RECT 63.625 103.275 63.795 103.445 ;
      RECT 63.165 103.275 63.335 103.445 ;
      RECT 62.705 103.275 62.875 103.445 ;
      RECT 62.245 103.275 62.415 103.445 ;
      RECT 61.785 103.275 61.955 103.445 ;
      RECT 61.325 103.275 61.495 103.445 ;
      RECT 60.865 103.275 61.035 103.445 ;
      RECT 60.405 103.275 60.575 103.445 ;
      RECT 59.945 103.275 60.115 103.445 ;
      RECT 59.485 103.275 59.655 103.445 ;
      RECT 59.025 103.275 59.195 103.445 ;
      RECT 58.565 103.275 58.735 103.445 ;
      RECT 58.105 103.275 58.275 103.445 ;
      RECT 57.645 103.275 57.815 103.445 ;
      RECT 57.185 103.275 57.355 103.445 ;
      RECT 56.725 103.275 56.895 103.445 ;
      RECT 56.265 103.275 56.435 103.445 ;
      RECT 55.805 103.275 55.975 103.445 ;
      RECT 55.345 103.275 55.515 103.445 ;
      RECT 54.885 103.275 55.055 103.445 ;
      RECT 54.425 103.275 54.595 103.445 ;
      RECT 53.965 103.275 54.135 103.445 ;
      RECT 53.505 103.275 53.675 103.445 ;
      RECT 53.045 103.275 53.215 103.445 ;
      RECT 52.585 103.275 52.755 103.445 ;
      RECT 52.125 103.275 52.295 103.445 ;
      RECT 51.665 103.275 51.835 103.445 ;
      RECT 51.205 103.275 51.375 103.445 ;
      RECT 50.745 103.275 50.915 103.445 ;
      RECT 50.285 103.275 50.455 103.445 ;
      RECT 49.825 103.275 49.995 103.445 ;
      RECT 49.365 103.275 49.535 103.445 ;
      RECT 48.905 103.275 49.075 103.445 ;
      RECT 48.445 103.275 48.615 103.445 ;
      RECT 47.985 103.275 48.155 103.445 ;
      RECT 47.525 103.275 47.695 103.445 ;
      RECT 47.065 103.275 47.235 103.445 ;
      RECT 46.605 103.275 46.775 103.445 ;
      RECT 46.145 103.275 46.315 103.445 ;
      RECT 45.685 103.275 45.855 103.445 ;
      RECT 45.225 103.275 45.395 103.445 ;
      RECT 44.765 103.275 44.935 103.445 ;
      RECT 44.305 103.275 44.475 103.445 ;
      RECT 43.845 103.275 44.015 103.445 ;
      RECT 43.385 103.275 43.555 103.445 ;
      RECT 42.925 103.275 43.095 103.445 ;
      RECT 42.465 103.275 42.635 103.445 ;
      RECT 42.005 103.275 42.175 103.445 ;
      RECT 41.545 103.275 41.715 103.445 ;
      RECT 41.085 103.275 41.255 103.445 ;
      RECT 40.625 103.275 40.795 103.445 ;
      RECT 40.165 103.275 40.335 103.445 ;
      RECT 39.705 103.275 39.875 103.445 ;
      RECT 39.245 103.275 39.415 103.445 ;
      RECT 38.785 103.275 38.955 103.445 ;
      RECT 38.325 103.275 38.495 103.445 ;
      RECT 37.865 103.275 38.035 103.445 ;
      RECT 37.405 103.275 37.575 103.445 ;
      RECT 36.945 103.275 37.115 103.445 ;
      RECT 36.485 103.275 36.655 103.445 ;
      RECT 36.025 103.275 36.195 103.445 ;
      RECT 35.565 103.275 35.735 103.445 ;
      RECT 35.105 103.275 35.275 103.445 ;
      RECT 34.645 103.275 34.815 103.445 ;
      RECT 34.185 103.275 34.355 103.445 ;
      RECT 33.725 103.275 33.895 103.445 ;
      RECT 33.265 103.275 33.435 103.445 ;
      RECT 32.805 103.275 32.975 103.445 ;
      RECT 32.345 103.275 32.515 103.445 ;
      RECT 31.885 103.275 32.055 103.445 ;
      RECT 31.425 103.275 31.595 103.445 ;
      RECT 30.965 103.275 31.135 103.445 ;
      RECT 30.505 103.275 30.675 103.445 ;
      RECT 30.045 103.275 30.215 103.445 ;
      RECT 29.585 103.275 29.755 103.445 ;
      RECT 29.125 103.275 29.295 103.445 ;
      RECT 28.665 103.275 28.835 103.445 ;
      RECT 28.205 103.275 28.375 103.445 ;
      RECT 27.745 103.275 27.915 103.445 ;
      RECT 27.285 103.275 27.455 103.445 ;
      RECT 26.825 103.275 26.995 103.445 ;
      RECT 26.365 103.275 26.535 103.445 ;
      RECT 25.905 103.275 26.075 103.445 ;
      RECT 25.445 103.275 25.615 103.445 ;
      RECT 24.985 103.275 25.155 103.445 ;
      RECT 24.525 103.275 24.695 103.445 ;
      RECT 24.065 103.275 24.235 103.445 ;
      RECT 23.605 103.275 23.775 103.445 ;
      RECT 23.145 103.275 23.315 103.445 ;
      RECT 22.685 103.275 22.855 103.445 ;
      RECT 22.225 103.275 22.395 103.445 ;
      RECT 21.765 103.275 21.935 103.445 ;
      RECT 21.305 103.275 21.475 103.445 ;
      RECT 20.845 103.275 21.015 103.445 ;
      RECT 20.385 103.275 20.555 103.445 ;
      RECT 19.925 103.275 20.095 103.445 ;
      RECT 19.465 103.275 19.635 103.445 ;
      RECT 19.005 103.275 19.175 103.445 ;
      RECT 18.545 103.275 18.715 103.445 ;
      RECT 18.085 103.275 18.255 103.445 ;
      RECT 17.625 103.275 17.795 103.445 ;
      RECT 17.165 103.275 17.335 103.445 ;
      RECT 16.705 103.275 16.875 103.445 ;
      RECT 16.245 103.275 16.415 103.445 ;
      RECT 15.785 103.275 15.955 103.445 ;
      RECT 15.325 103.275 15.495 103.445 ;
      RECT 14.865 103.275 15.035 103.445 ;
      RECT 14.405 103.275 14.575 103.445 ;
      RECT 13.945 103.275 14.115 103.445 ;
      RECT 13.485 103.275 13.655 103.445 ;
      RECT 13.025 103.275 13.195 103.445 ;
      RECT 12.565 103.275 12.735 103.445 ;
      RECT 12.105 103.275 12.275 103.445 ;
      RECT 11.645 103.275 11.815 103.445 ;
      RECT 11.185 103.275 11.355 103.445 ;
      RECT 10.725 103.275 10.895 103.445 ;
      RECT 10.265 103.275 10.435 103.445 ;
      RECT 9.805 103.275 9.975 103.445 ;
      RECT 9.345 103.275 9.515 103.445 ;
      RECT 8.885 103.275 9.055 103.445 ;
      RECT 8.425 103.275 8.595 103.445 ;
      RECT 7.965 103.275 8.135 103.445 ;
      RECT 7.505 103.275 7.675 103.445 ;
      RECT 7.045 103.275 7.215 103.445 ;
      RECT 6.585 103.275 6.755 103.445 ;
      RECT 6.125 103.275 6.295 103.445 ;
      RECT 5.665 103.275 5.835 103.445 ;
      RECT 5.205 103.275 5.375 103.445 ;
      RECT 4.745 103.275 4.915 103.445 ;
      RECT 4.285 103.275 4.455 103.445 ;
      RECT 3.825 103.275 3.995 103.445 ;
      RECT 3.365 103.275 3.535 103.445 ;
      RECT 2.905 103.275 3.075 103.445 ;
      RECT 2.445 103.275 2.615 103.445 ;
      RECT 1.985 103.275 2.155 103.445 ;
      RECT 1.525 103.275 1.695 103.445 ;
      RECT 1.065 103.275 1.235 103.445 ;
      RECT 0.605 103.275 0.775 103.445 ;
      RECT 0.145 103.275 0.315 103.445 ;
      RECT 112.845 100.555 113.015 100.725 ;
      RECT 112.385 100.555 112.555 100.725 ;
      RECT 0.605 100.555 0.775 100.725 ;
      RECT 0.145 100.555 0.315 100.725 ;
      RECT 112.845 97.835 113.015 98.005 ;
      RECT 112.385 97.835 112.555 98.005 ;
      RECT 0.605 97.835 0.775 98.005 ;
      RECT 0.145 97.835 0.315 98.005 ;
      RECT 112.845 95.115 113.015 95.285 ;
      RECT 112.385 95.115 112.555 95.285 ;
      RECT 0.605 95.115 0.775 95.285 ;
      RECT 0.145 95.115 0.315 95.285 ;
      RECT 112.845 92.395 113.015 92.565 ;
      RECT 112.385 92.395 112.555 92.565 ;
      RECT 0.605 92.395 0.775 92.565 ;
      RECT 0.145 92.395 0.315 92.565 ;
      RECT 112.845 89.675 113.015 89.845 ;
      RECT 112.385 89.675 112.555 89.845 ;
      RECT 0.605 89.675 0.775 89.845 ;
      RECT 0.145 89.675 0.315 89.845 ;
      RECT 112.845 86.955 113.015 87.125 ;
      RECT 112.385 86.955 112.555 87.125 ;
      RECT 0.605 86.955 0.775 87.125 ;
      RECT 0.145 86.955 0.315 87.125 ;
      RECT 112.845 84.235 113.015 84.405 ;
      RECT 112.385 84.235 112.555 84.405 ;
      RECT 0.605 84.235 0.775 84.405 ;
      RECT 0.145 84.235 0.315 84.405 ;
      RECT 112.845 81.515 113.015 81.685 ;
      RECT 112.385 81.515 112.555 81.685 ;
      RECT 0.605 81.515 0.775 81.685 ;
      RECT 0.145 81.515 0.315 81.685 ;
      RECT 112.845 78.795 113.015 78.965 ;
      RECT 112.385 78.795 112.555 78.965 ;
      RECT 0.605 78.795 0.775 78.965 ;
      RECT 0.145 78.795 0.315 78.965 ;
      RECT 112.845 76.075 113.015 76.245 ;
      RECT 112.385 76.075 112.555 76.245 ;
      RECT 0.605 76.075 0.775 76.245 ;
      RECT 0.145 76.075 0.315 76.245 ;
      RECT 112.845 73.355 113.015 73.525 ;
      RECT 112.385 73.355 112.555 73.525 ;
      RECT 0.605 73.355 0.775 73.525 ;
      RECT 0.145 73.355 0.315 73.525 ;
      RECT 112.845 70.635 113.015 70.805 ;
      RECT 112.385 70.635 112.555 70.805 ;
      RECT 0.605 70.635 0.775 70.805 ;
      RECT 0.145 70.635 0.315 70.805 ;
      RECT 112.845 67.915 113.015 68.085 ;
      RECT 112.385 67.915 112.555 68.085 ;
      RECT 0.605 67.915 0.775 68.085 ;
      RECT 0.145 67.915 0.315 68.085 ;
      RECT 112.845 65.195 113.015 65.365 ;
      RECT 112.385 65.195 112.555 65.365 ;
      RECT 0.605 65.195 0.775 65.365 ;
      RECT 0.145 65.195 0.315 65.365 ;
      RECT 112.845 62.475 113.015 62.645 ;
      RECT 112.385 62.475 112.555 62.645 ;
      RECT 0.605 62.475 0.775 62.645 ;
      RECT 0.145 62.475 0.315 62.645 ;
      RECT 112.845 59.755 113.015 59.925 ;
      RECT 112.385 59.755 112.555 59.925 ;
      RECT 0.605 59.755 0.775 59.925 ;
      RECT 0.145 59.755 0.315 59.925 ;
      RECT 112.845 57.035 113.015 57.205 ;
      RECT 112.385 57.035 112.555 57.205 ;
      RECT 0.605 57.035 0.775 57.205 ;
      RECT 0.145 57.035 0.315 57.205 ;
      RECT 112.845 54.315 113.015 54.485 ;
      RECT 112.385 54.315 112.555 54.485 ;
      RECT 0.605 54.315 0.775 54.485 ;
      RECT 0.145 54.315 0.315 54.485 ;
      RECT 112.845 51.595 113.015 51.765 ;
      RECT 112.385 51.595 112.555 51.765 ;
      RECT 0.605 51.595 0.775 51.765 ;
      RECT 0.145 51.595 0.315 51.765 ;
      RECT 112.845 48.875 113.015 49.045 ;
      RECT 112.385 48.875 112.555 49.045 ;
      RECT 0.605 48.875 0.775 49.045 ;
      RECT 0.145 48.875 0.315 49.045 ;
      RECT 112.845 46.155 113.015 46.325 ;
      RECT 112.385 46.155 112.555 46.325 ;
      RECT 0.605 46.155 0.775 46.325 ;
      RECT 0.145 46.155 0.315 46.325 ;
      RECT 112.845 43.435 113.015 43.605 ;
      RECT 112.385 43.435 112.555 43.605 ;
      RECT 0.605 43.435 0.775 43.605 ;
      RECT 0.145 43.435 0.315 43.605 ;
      RECT 112.845 40.715 113.015 40.885 ;
      RECT 112.385 40.715 112.555 40.885 ;
      RECT 0.605 40.715 0.775 40.885 ;
      RECT 0.145 40.715 0.315 40.885 ;
      RECT 112.845 37.995 113.015 38.165 ;
      RECT 112.385 37.995 112.555 38.165 ;
      RECT 0.605 37.995 0.775 38.165 ;
      RECT 0.145 37.995 0.315 38.165 ;
      RECT 112.845 35.275 113.015 35.445 ;
      RECT 112.385 35.275 112.555 35.445 ;
      RECT 0.605 35.275 0.775 35.445 ;
      RECT 0.145 35.275 0.315 35.445 ;
      RECT 112.845 32.555 113.015 32.725 ;
      RECT 112.385 32.555 112.555 32.725 ;
      RECT 0.605 32.555 0.775 32.725 ;
      RECT 0.145 32.555 0.315 32.725 ;
      RECT 112.845 29.835 113.015 30.005 ;
      RECT 112.385 29.835 112.555 30.005 ;
      RECT 0.605 29.835 0.775 30.005 ;
      RECT 0.145 29.835 0.315 30.005 ;
      RECT 112.845 27.115 113.015 27.285 ;
      RECT 112.385 27.115 112.555 27.285 ;
      RECT 111.925 27.115 112.095 27.285 ;
      RECT 111.465 27.115 111.635 27.285 ;
      RECT 111.005 27.115 111.175 27.285 ;
      RECT 110.545 27.115 110.715 27.285 ;
      RECT 110.085 27.115 110.255 27.285 ;
      RECT 109.625 27.115 109.795 27.285 ;
      RECT 109.165 27.115 109.335 27.285 ;
      RECT 108.705 27.115 108.875 27.285 ;
      RECT 108.245 27.115 108.415 27.285 ;
      RECT 107.785 27.115 107.955 27.285 ;
      RECT 107.325 27.115 107.495 27.285 ;
      RECT 106.865 27.115 107.035 27.285 ;
      RECT 106.405 27.115 106.575 27.285 ;
      RECT 105.945 27.115 106.115 27.285 ;
      RECT 105.485 27.115 105.655 27.285 ;
      RECT 105.025 27.115 105.195 27.285 ;
      RECT 104.565 27.115 104.735 27.285 ;
      RECT 104.105 27.115 104.275 27.285 ;
      RECT 103.645 27.115 103.815 27.285 ;
      RECT 103.185 27.115 103.355 27.285 ;
      RECT 102.725 27.115 102.895 27.285 ;
      RECT 102.265 27.115 102.435 27.285 ;
      RECT 101.805 27.115 101.975 27.285 ;
      RECT 101.345 27.115 101.515 27.285 ;
      RECT 100.885 27.115 101.055 27.285 ;
      RECT 100.425 27.115 100.595 27.285 ;
      RECT 99.965 27.115 100.135 27.285 ;
      RECT 99.505 27.115 99.675 27.285 ;
      RECT 99.045 27.115 99.215 27.285 ;
      RECT 98.585 27.115 98.755 27.285 ;
      RECT 98.125 27.115 98.295 27.285 ;
      RECT 97.665 27.115 97.835 27.285 ;
      RECT 97.205 27.115 97.375 27.285 ;
      RECT 96.745 27.115 96.915 27.285 ;
      RECT 96.285 27.115 96.455 27.285 ;
      RECT 95.825 27.115 95.995 27.285 ;
      RECT 95.365 27.115 95.535 27.285 ;
      RECT 94.905 27.115 95.075 27.285 ;
      RECT 94.445 27.115 94.615 27.285 ;
      RECT 93.985 27.115 94.155 27.285 ;
      RECT 93.525 27.115 93.695 27.285 ;
      RECT 93.065 27.115 93.235 27.285 ;
      RECT 92.605 27.115 92.775 27.285 ;
      RECT 92.145 27.115 92.315 27.285 ;
      RECT 91.685 27.115 91.855 27.285 ;
      RECT 91.225 27.115 91.395 27.285 ;
      RECT 90.765 27.115 90.935 27.285 ;
      RECT 90.305 27.115 90.475 27.285 ;
      RECT 89.845 27.115 90.015 27.285 ;
      RECT 89.385 27.115 89.555 27.285 ;
      RECT 88.925 27.115 89.095 27.285 ;
      RECT 88.465 27.115 88.635 27.285 ;
      RECT 88.005 27.115 88.175 27.285 ;
      RECT 87.545 27.115 87.715 27.285 ;
      RECT 87.085 27.115 87.255 27.285 ;
      RECT 86.625 27.115 86.795 27.285 ;
      RECT 86.165 27.115 86.335 27.285 ;
      RECT 85.705 27.115 85.875 27.285 ;
      RECT 85.245 27.115 85.415 27.285 ;
      RECT 84.785 27.115 84.955 27.285 ;
      RECT 84.325 27.115 84.495 27.285 ;
      RECT 83.865 27.115 84.035 27.285 ;
      RECT 83.405 27.115 83.575 27.285 ;
      RECT 82.945 27.115 83.115 27.285 ;
      RECT 82.485 27.115 82.655 27.285 ;
      RECT 82.025 27.115 82.195 27.285 ;
      RECT 81.565 27.115 81.735 27.285 ;
      RECT 81.105 27.115 81.275 27.285 ;
      RECT 80.645 27.115 80.815 27.285 ;
      RECT 80.185 27.115 80.355 27.285 ;
      RECT 79.725 27.115 79.895 27.285 ;
      RECT 79.265 27.115 79.435 27.285 ;
      RECT 78.805 27.115 78.975 27.285 ;
      RECT 78.345 27.115 78.515 27.285 ;
      RECT 77.885 27.115 78.055 27.285 ;
      RECT 77.425 27.115 77.595 27.285 ;
      RECT 76.965 27.115 77.135 27.285 ;
      RECT 76.505 27.115 76.675 27.285 ;
      RECT 76.045 27.115 76.215 27.285 ;
      RECT 75.585 27.115 75.755 27.285 ;
      RECT 75.125 27.115 75.295 27.285 ;
      RECT 74.665 27.115 74.835 27.285 ;
      RECT 74.205 27.115 74.375 27.285 ;
      RECT 73.745 27.115 73.915 27.285 ;
      RECT 73.285 27.115 73.455 27.285 ;
      RECT 72.825 27.115 72.995 27.285 ;
      RECT 72.365 27.115 72.535 27.285 ;
      RECT 71.905 27.115 72.075 27.285 ;
      RECT 71.445 27.115 71.615 27.285 ;
      RECT 70.985 27.115 71.155 27.285 ;
      RECT 70.525 27.115 70.695 27.285 ;
      RECT 70.065 27.115 70.235 27.285 ;
      RECT 69.605 27.115 69.775 27.285 ;
      RECT 69.145 27.115 69.315 27.285 ;
      RECT 68.685 27.115 68.855 27.285 ;
      RECT 68.225 27.115 68.395 27.285 ;
      RECT 67.765 27.115 67.935 27.285 ;
      RECT 67.305 27.115 67.475 27.285 ;
      RECT 66.845 27.115 67.015 27.285 ;
      RECT 66.385 27.115 66.555 27.285 ;
      RECT 65.925 27.115 66.095 27.285 ;
      RECT 65.465 27.115 65.635 27.285 ;
      RECT 65.005 27.115 65.175 27.285 ;
      RECT 64.545 27.115 64.715 27.285 ;
      RECT 64.085 27.115 64.255 27.285 ;
      RECT 63.625 27.115 63.795 27.285 ;
      RECT 63.165 27.115 63.335 27.285 ;
      RECT 62.705 27.115 62.875 27.285 ;
      RECT 62.245 27.115 62.415 27.285 ;
      RECT 61.785 27.115 61.955 27.285 ;
      RECT 61.325 27.115 61.495 27.285 ;
      RECT 60.865 27.115 61.035 27.285 ;
      RECT 60.405 27.115 60.575 27.285 ;
      RECT 59.945 27.115 60.115 27.285 ;
      RECT 59.485 27.115 59.655 27.285 ;
      RECT 59.025 27.115 59.195 27.285 ;
      RECT 58.565 27.115 58.735 27.285 ;
      RECT 58.105 27.115 58.275 27.285 ;
      RECT 57.645 27.115 57.815 27.285 ;
      RECT 57.185 27.115 57.355 27.285 ;
      RECT 56.725 27.115 56.895 27.285 ;
      RECT 56.265 27.115 56.435 27.285 ;
      RECT 55.805 27.115 55.975 27.285 ;
      RECT 55.345 27.115 55.515 27.285 ;
      RECT 54.885 27.115 55.055 27.285 ;
      RECT 54.425 27.115 54.595 27.285 ;
      RECT 53.965 27.115 54.135 27.285 ;
      RECT 53.505 27.115 53.675 27.285 ;
      RECT 53.045 27.115 53.215 27.285 ;
      RECT 52.585 27.115 52.755 27.285 ;
      RECT 52.125 27.115 52.295 27.285 ;
      RECT 51.665 27.115 51.835 27.285 ;
      RECT 51.205 27.115 51.375 27.285 ;
      RECT 50.745 27.115 50.915 27.285 ;
      RECT 50.285 27.115 50.455 27.285 ;
      RECT 49.825 27.115 49.995 27.285 ;
      RECT 49.365 27.115 49.535 27.285 ;
      RECT 48.905 27.115 49.075 27.285 ;
      RECT 48.445 27.115 48.615 27.285 ;
      RECT 47.985 27.115 48.155 27.285 ;
      RECT 47.525 27.115 47.695 27.285 ;
      RECT 47.065 27.115 47.235 27.285 ;
      RECT 46.605 27.115 46.775 27.285 ;
      RECT 46.145 27.115 46.315 27.285 ;
      RECT 45.685 27.115 45.855 27.285 ;
      RECT 45.225 27.115 45.395 27.285 ;
      RECT 44.765 27.115 44.935 27.285 ;
      RECT 44.305 27.115 44.475 27.285 ;
      RECT 43.845 27.115 44.015 27.285 ;
      RECT 43.385 27.115 43.555 27.285 ;
      RECT 42.925 27.115 43.095 27.285 ;
      RECT 42.465 27.115 42.635 27.285 ;
      RECT 42.005 27.115 42.175 27.285 ;
      RECT 41.545 27.115 41.715 27.285 ;
      RECT 41.085 27.115 41.255 27.285 ;
      RECT 40.625 27.115 40.795 27.285 ;
      RECT 40.165 27.115 40.335 27.285 ;
      RECT 39.705 27.115 39.875 27.285 ;
      RECT 39.245 27.115 39.415 27.285 ;
      RECT 38.785 27.115 38.955 27.285 ;
      RECT 38.325 27.115 38.495 27.285 ;
      RECT 37.865 27.115 38.035 27.285 ;
      RECT 37.405 27.115 37.575 27.285 ;
      RECT 36.945 27.115 37.115 27.285 ;
      RECT 36.485 27.115 36.655 27.285 ;
      RECT 36.025 27.115 36.195 27.285 ;
      RECT 35.565 27.115 35.735 27.285 ;
      RECT 35.105 27.115 35.275 27.285 ;
      RECT 34.645 27.115 34.815 27.285 ;
      RECT 34.185 27.115 34.355 27.285 ;
      RECT 33.725 27.115 33.895 27.285 ;
      RECT 33.265 27.115 33.435 27.285 ;
      RECT 32.805 27.115 32.975 27.285 ;
      RECT 32.345 27.115 32.515 27.285 ;
      RECT 31.885 27.115 32.055 27.285 ;
      RECT 31.425 27.115 31.595 27.285 ;
      RECT 30.965 27.115 31.135 27.285 ;
      RECT 30.505 27.115 30.675 27.285 ;
      RECT 30.045 27.115 30.215 27.285 ;
      RECT 29.585 27.115 29.755 27.285 ;
      RECT 29.125 27.115 29.295 27.285 ;
      RECT 28.665 27.115 28.835 27.285 ;
      RECT 28.205 27.115 28.375 27.285 ;
      RECT 27.745 27.115 27.915 27.285 ;
      RECT 27.285 27.115 27.455 27.285 ;
      RECT 26.825 27.115 26.995 27.285 ;
      RECT 26.365 27.115 26.535 27.285 ;
      RECT 25.905 27.115 26.075 27.285 ;
      RECT 25.445 27.115 25.615 27.285 ;
      RECT 24.985 27.115 25.155 27.285 ;
      RECT 24.525 27.115 24.695 27.285 ;
      RECT 24.065 27.115 24.235 27.285 ;
      RECT 23.605 27.115 23.775 27.285 ;
      RECT 23.145 27.115 23.315 27.285 ;
      RECT 22.685 27.115 22.855 27.285 ;
      RECT 22.225 27.115 22.395 27.285 ;
      RECT 21.765 27.115 21.935 27.285 ;
      RECT 21.305 27.115 21.475 27.285 ;
      RECT 20.845 27.115 21.015 27.285 ;
      RECT 20.385 27.115 20.555 27.285 ;
      RECT 19.925 27.115 20.095 27.285 ;
      RECT 19.465 27.115 19.635 27.285 ;
      RECT 19.005 27.115 19.175 27.285 ;
      RECT 18.545 27.115 18.715 27.285 ;
      RECT 18.085 27.115 18.255 27.285 ;
      RECT 17.625 27.115 17.795 27.285 ;
      RECT 17.165 27.115 17.335 27.285 ;
      RECT 16.705 27.115 16.875 27.285 ;
      RECT 16.245 27.115 16.415 27.285 ;
      RECT 15.785 27.115 15.955 27.285 ;
      RECT 15.325 27.115 15.495 27.285 ;
      RECT 14.865 27.115 15.035 27.285 ;
      RECT 14.405 27.115 14.575 27.285 ;
      RECT 13.945 27.115 14.115 27.285 ;
      RECT 13.485 27.115 13.655 27.285 ;
      RECT 13.025 27.115 13.195 27.285 ;
      RECT 12.565 27.115 12.735 27.285 ;
      RECT 12.105 27.115 12.275 27.285 ;
      RECT 11.645 27.115 11.815 27.285 ;
      RECT 11.185 27.115 11.355 27.285 ;
      RECT 10.725 27.115 10.895 27.285 ;
      RECT 10.265 27.115 10.435 27.285 ;
      RECT 9.805 27.115 9.975 27.285 ;
      RECT 9.345 27.115 9.515 27.285 ;
      RECT 8.885 27.115 9.055 27.285 ;
      RECT 8.425 27.115 8.595 27.285 ;
      RECT 7.965 27.115 8.135 27.285 ;
      RECT 7.505 27.115 7.675 27.285 ;
      RECT 7.045 27.115 7.215 27.285 ;
      RECT 6.585 27.115 6.755 27.285 ;
      RECT 6.125 27.115 6.295 27.285 ;
      RECT 5.665 27.115 5.835 27.285 ;
      RECT 5.205 27.115 5.375 27.285 ;
      RECT 4.745 27.115 4.915 27.285 ;
      RECT 4.285 27.115 4.455 27.285 ;
      RECT 3.825 27.115 3.995 27.285 ;
      RECT 3.365 27.115 3.535 27.285 ;
      RECT 2.905 27.115 3.075 27.285 ;
      RECT 2.445 27.115 2.615 27.285 ;
      RECT 1.985 27.115 2.155 27.285 ;
      RECT 1.525 27.115 1.695 27.285 ;
      RECT 1.065 27.115 1.235 27.285 ;
      RECT 0.605 27.115 0.775 27.285 ;
      RECT 0.145 27.115 0.315 27.285 ;
      RECT 84.325 24.395 84.495 24.565 ;
      RECT 83.865 24.395 84.035 24.565 ;
      RECT 0.605 24.395 0.775 24.565 ;
      RECT 0.145 24.395 0.315 24.565 ;
      RECT 84.325 21.675 84.495 21.845 ;
      RECT 83.865 21.675 84.035 21.845 ;
      RECT 0.605 21.675 0.775 21.845 ;
      RECT 0.145 21.675 0.315 21.845 ;
      RECT 84.325 18.955 84.495 19.125 ;
      RECT 83.865 18.955 84.035 19.125 ;
      RECT 0.605 18.955 0.775 19.125 ;
      RECT 0.145 18.955 0.315 19.125 ;
      RECT 84.325 16.235 84.495 16.405 ;
      RECT 83.865 16.235 84.035 16.405 ;
      RECT 0.605 16.235 0.775 16.405 ;
      RECT 0.145 16.235 0.315 16.405 ;
      RECT 84.325 13.515 84.495 13.685 ;
      RECT 83.865 13.515 84.035 13.685 ;
      RECT 0.605 13.515 0.775 13.685 ;
      RECT 0.145 13.515 0.315 13.685 ;
      RECT 84.325 10.795 84.495 10.965 ;
      RECT 83.865 10.795 84.035 10.965 ;
      RECT 0.605 10.795 0.775 10.965 ;
      RECT 0.145 10.795 0.315 10.965 ;
      RECT 84.325 8.075 84.495 8.245 ;
      RECT 83.865 8.075 84.035 8.245 ;
      RECT 0.605 8.075 0.775 8.245 ;
      RECT 0.145 8.075 0.315 8.245 ;
      RECT 84.325 5.355 84.495 5.525 ;
      RECT 83.865 5.355 84.035 5.525 ;
      RECT 0.605 5.355 0.775 5.525 ;
      RECT 0.145 5.355 0.315 5.525 ;
      RECT 84.325 2.635 84.495 2.805 ;
      RECT 83.865 2.635 84.035 2.805 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 84.325 -0.085 84.495 0.085 ;
      RECT 83.865 -0.085 84.035 0.085 ;
      RECT 83.405 -0.085 83.575 0.085 ;
      RECT 82.945 -0.085 83.115 0.085 ;
      RECT 82.485 -0.085 82.655 0.085 ;
      RECT 82.025 -0.085 82.195 0.085 ;
      RECT 81.565 -0.085 81.735 0.085 ;
      RECT 81.105 -0.085 81.275 0.085 ;
      RECT 80.645 -0.085 80.815 0.085 ;
      RECT 80.185 -0.085 80.355 0.085 ;
      RECT 79.725 -0.085 79.895 0.085 ;
      RECT 79.265 -0.085 79.435 0.085 ;
      RECT 78.805 -0.085 78.975 0.085 ;
      RECT 78.345 -0.085 78.515 0.085 ;
      RECT 77.885 -0.085 78.055 0.085 ;
      RECT 77.425 -0.085 77.595 0.085 ;
      RECT 76.965 -0.085 77.135 0.085 ;
      RECT 76.505 -0.085 76.675 0.085 ;
      RECT 76.045 -0.085 76.215 0.085 ;
      RECT 75.585 -0.085 75.755 0.085 ;
      RECT 75.125 -0.085 75.295 0.085 ;
      RECT 74.665 -0.085 74.835 0.085 ;
      RECT 74.205 -0.085 74.375 0.085 ;
      RECT 73.745 -0.085 73.915 0.085 ;
      RECT 73.285 -0.085 73.455 0.085 ;
      RECT 72.825 -0.085 72.995 0.085 ;
      RECT 72.365 -0.085 72.535 0.085 ;
      RECT 71.905 -0.085 72.075 0.085 ;
      RECT 71.445 -0.085 71.615 0.085 ;
      RECT 70.985 -0.085 71.155 0.085 ;
      RECT 70.525 -0.085 70.695 0.085 ;
      RECT 70.065 -0.085 70.235 0.085 ;
      RECT 69.605 -0.085 69.775 0.085 ;
      RECT 69.145 -0.085 69.315 0.085 ;
      RECT 68.685 -0.085 68.855 0.085 ;
      RECT 68.225 -0.085 68.395 0.085 ;
      RECT 67.765 -0.085 67.935 0.085 ;
      RECT 67.305 -0.085 67.475 0.085 ;
      RECT 66.845 -0.085 67.015 0.085 ;
      RECT 66.385 -0.085 66.555 0.085 ;
      RECT 65.925 -0.085 66.095 0.085 ;
      RECT 65.465 -0.085 65.635 0.085 ;
      RECT 65.005 -0.085 65.175 0.085 ;
      RECT 64.545 -0.085 64.715 0.085 ;
      RECT 64.085 -0.085 64.255 0.085 ;
      RECT 63.625 -0.085 63.795 0.085 ;
      RECT 63.165 -0.085 63.335 0.085 ;
      RECT 62.705 -0.085 62.875 0.085 ;
      RECT 62.245 -0.085 62.415 0.085 ;
      RECT 61.785 -0.085 61.955 0.085 ;
      RECT 61.325 -0.085 61.495 0.085 ;
      RECT 60.865 -0.085 61.035 0.085 ;
      RECT 60.405 -0.085 60.575 0.085 ;
      RECT 59.945 -0.085 60.115 0.085 ;
      RECT 59.485 -0.085 59.655 0.085 ;
      RECT 59.025 -0.085 59.195 0.085 ;
      RECT 58.565 -0.085 58.735 0.085 ;
      RECT 58.105 -0.085 58.275 0.085 ;
      RECT 57.645 -0.085 57.815 0.085 ;
      RECT 57.185 -0.085 57.355 0.085 ;
      RECT 56.725 -0.085 56.895 0.085 ;
      RECT 56.265 -0.085 56.435 0.085 ;
      RECT 55.805 -0.085 55.975 0.085 ;
      RECT 55.345 -0.085 55.515 0.085 ;
      RECT 54.885 -0.085 55.055 0.085 ;
      RECT 54.425 -0.085 54.595 0.085 ;
      RECT 53.965 -0.085 54.135 0.085 ;
      RECT 53.505 -0.085 53.675 0.085 ;
      RECT 53.045 -0.085 53.215 0.085 ;
      RECT 52.585 -0.085 52.755 0.085 ;
      RECT 52.125 -0.085 52.295 0.085 ;
      RECT 51.665 -0.085 51.835 0.085 ;
      RECT 51.205 -0.085 51.375 0.085 ;
      RECT 50.745 -0.085 50.915 0.085 ;
      RECT 50.285 -0.085 50.455 0.085 ;
      RECT 49.825 -0.085 49.995 0.085 ;
      RECT 49.365 -0.085 49.535 0.085 ;
      RECT 48.905 -0.085 49.075 0.085 ;
      RECT 48.445 -0.085 48.615 0.085 ;
      RECT 47.985 -0.085 48.155 0.085 ;
      RECT 47.525 -0.085 47.695 0.085 ;
      RECT 47.065 -0.085 47.235 0.085 ;
      RECT 46.605 -0.085 46.775 0.085 ;
      RECT 46.145 -0.085 46.315 0.085 ;
      RECT 45.685 -0.085 45.855 0.085 ;
      RECT 45.225 -0.085 45.395 0.085 ;
      RECT 44.765 -0.085 44.935 0.085 ;
      RECT 44.305 -0.085 44.475 0.085 ;
      RECT 43.845 -0.085 44.015 0.085 ;
      RECT 43.385 -0.085 43.555 0.085 ;
      RECT 42.925 -0.085 43.095 0.085 ;
      RECT 42.465 -0.085 42.635 0.085 ;
      RECT 42.005 -0.085 42.175 0.085 ;
      RECT 41.545 -0.085 41.715 0.085 ;
      RECT 41.085 -0.085 41.255 0.085 ;
      RECT 40.625 -0.085 40.795 0.085 ;
      RECT 40.165 -0.085 40.335 0.085 ;
      RECT 39.705 -0.085 39.875 0.085 ;
      RECT 39.245 -0.085 39.415 0.085 ;
      RECT 38.785 -0.085 38.955 0.085 ;
      RECT 38.325 -0.085 38.495 0.085 ;
      RECT 37.865 -0.085 38.035 0.085 ;
      RECT 37.405 -0.085 37.575 0.085 ;
      RECT 36.945 -0.085 37.115 0.085 ;
      RECT 36.485 -0.085 36.655 0.085 ;
      RECT 36.025 -0.085 36.195 0.085 ;
      RECT 35.565 -0.085 35.735 0.085 ;
      RECT 35.105 -0.085 35.275 0.085 ;
      RECT 34.645 -0.085 34.815 0.085 ;
      RECT 34.185 -0.085 34.355 0.085 ;
      RECT 33.725 -0.085 33.895 0.085 ;
      RECT 33.265 -0.085 33.435 0.085 ;
      RECT 32.805 -0.085 32.975 0.085 ;
      RECT 32.345 -0.085 32.515 0.085 ;
      RECT 31.885 -0.085 32.055 0.085 ;
      RECT 31.425 -0.085 31.595 0.085 ;
      RECT 30.965 -0.085 31.135 0.085 ;
      RECT 30.505 -0.085 30.675 0.085 ;
      RECT 30.045 -0.085 30.215 0.085 ;
      RECT 29.585 -0.085 29.755 0.085 ;
      RECT 29.125 -0.085 29.295 0.085 ;
      RECT 28.665 -0.085 28.835 0.085 ;
      RECT 28.205 -0.085 28.375 0.085 ;
      RECT 27.745 -0.085 27.915 0.085 ;
      RECT 27.285 -0.085 27.455 0.085 ;
      RECT 26.825 -0.085 26.995 0.085 ;
      RECT 26.365 -0.085 26.535 0.085 ;
      RECT 25.905 -0.085 26.075 0.085 ;
      RECT 25.445 -0.085 25.615 0.085 ;
      RECT 24.985 -0.085 25.155 0.085 ;
      RECT 24.525 -0.085 24.695 0.085 ;
      RECT 24.065 -0.085 24.235 0.085 ;
      RECT 23.605 -0.085 23.775 0.085 ;
      RECT 23.145 -0.085 23.315 0.085 ;
      RECT 22.685 -0.085 22.855 0.085 ;
      RECT 22.225 -0.085 22.395 0.085 ;
      RECT 21.765 -0.085 21.935 0.085 ;
      RECT 21.305 -0.085 21.475 0.085 ;
      RECT 20.845 -0.085 21.015 0.085 ;
      RECT 20.385 -0.085 20.555 0.085 ;
      RECT 19.925 -0.085 20.095 0.085 ;
      RECT 19.465 -0.085 19.635 0.085 ;
      RECT 19.005 -0.085 19.175 0.085 ;
      RECT 18.545 -0.085 18.715 0.085 ;
      RECT 18.085 -0.085 18.255 0.085 ;
      RECT 17.625 -0.085 17.795 0.085 ;
      RECT 17.165 -0.085 17.335 0.085 ;
      RECT 16.705 -0.085 16.875 0.085 ;
      RECT 16.245 -0.085 16.415 0.085 ;
      RECT 15.785 -0.085 15.955 0.085 ;
      RECT 15.325 -0.085 15.495 0.085 ;
      RECT 14.865 -0.085 15.035 0.085 ;
      RECT 14.405 -0.085 14.575 0.085 ;
      RECT 13.945 -0.085 14.115 0.085 ;
      RECT 13.485 -0.085 13.655 0.085 ;
      RECT 13.025 -0.085 13.195 0.085 ;
      RECT 12.565 -0.085 12.735 0.085 ;
      RECT 12.105 -0.085 12.275 0.085 ;
      RECT 11.645 -0.085 11.815 0.085 ;
      RECT 11.185 -0.085 11.355 0.085 ;
      RECT 10.725 -0.085 10.895 0.085 ;
      RECT 10.265 -0.085 10.435 0.085 ;
      RECT 9.805 -0.085 9.975 0.085 ;
      RECT 9.345 -0.085 9.515 0.085 ;
      RECT 8.885 -0.085 9.055 0.085 ;
      RECT 8.425 -0.085 8.595 0.085 ;
      RECT 7.965 -0.085 8.135 0.085 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.145 -0.085 0.315 0.085 ;
    LAYER via ;
      RECT 56.965 103.285 57.115 103.435 ;
      RECT 27.525 103.285 27.675 103.435 ;
      RECT 109.865 101.585 110.015 101.735 ;
      RECT 56.965 27.125 57.115 27.275 ;
      RECT 27.525 27.125 27.675 27.275 ;
      RECT 54.205 1.625 54.355 1.775 ;
      RECT 22.925 1.625 23.075 1.775 ;
      RECT 56.965 -0.075 57.115 0.075 ;
      RECT 27.525 -0.075 27.675 0.075 ;
    LAYER via2 ;
      RECT 56.94 103.26 57.14 103.46 ;
      RECT 27.5 103.26 27.7 103.46 ;
      RECT 111.68 93.74 111.88 93.94 ;
      RECT 111.68 88.3 111.88 88.5 ;
      RECT 111.68 82.86 111.88 83.06 ;
      RECT 111.68 50.22 111.88 50.42 ;
      RECT 111.22 47.5 111.42 47.7 ;
      RECT 111.68 46.14 111.88 46.34 ;
      RECT 111.68 42.06 111.88 42.26 ;
      RECT 56.94 -0.1 57.14 0.1 ;
      RECT 27.5 -0.1 27.7 0.1 ;
    LAYER via3 ;
      RECT 56.94 103.26 57.14 103.46 ;
      RECT 27.5 103.26 27.7 103.46 ;
      RECT 56.94 -0.1 57.14 0.1 ;
      RECT 27.5 -0.1 27.7 0.1 ;
    LAYER via4 ;
      RECT 106.32 86.08 107.12 86.88 ;
      RECT 106.32 84.48 107.12 85.28 ;
      RECT 106.32 45.28 107.12 46.08 ;
      RECT 106.32 43.68 107.12 44.48 ;
    LAYER fieldpoly ;
      POLYGON 113.02 103.22 113.02 27.34 84.5 27.34 84.5 0.14 0.14 0.14 0.14 103.22 ;
    LAYER diff ;
      POLYGON 113.16 103.36 113.16 27.2 84.64 27.2 84.64 0 0 0 0 103.36 ;
    LAYER nwell ;
      RECT 112.05 99.225 113.35 102.055 ;
      RECT -0.19 99.225 3.87 102.055 ;
      RECT 112.05 93.785 113.35 96.615 ;
      RECT -0.19 93.785 3.87 96.615 ;
      RECT 112.05 88.345 113.35 91.175 ;
      RECT -0.19 88.345 3.87 91.175 ;
      RECT 112.05 82.905 113.35 85.735 ;
      RECT -0.19 82.905 3.87 85.735 ;
      POLYGON 113.35 80.295 113.35 77.465 112.51 77.465 112.51 78.69 112.05 78.69 112.05 80.295 ;
      RECT -0.19 77.465 3.87 80.295 ;
      RECT 112.05 72.025 113.35 74.855 ;
      RECT -0.19 72.025 3.87 74.855 ;
      RECT 112.05 66.585 113.35 69.415 ;
      RECT -0.19 66.585 3.87 69.415 ;
      RECT 112.05 61.145 113.35 63.975 ;
      RECT -0.19 61.145 3.87 63.975 ;
      POLYGON 113.35 58.535 113.35 55.705 112.05 55.705 112.05 57.31 112.51 57.31 112.51 58.535 ;
      RECT -0.19 55.705 3.87 58.535 ;
      RECT 112.05 50.265 113.35 53.095 ;
      RECT -0.19 50.265 3.87 53.095 ;
      RECT 112.05 44.825 113.35 47.655 ;
      RECT -0.19 44.825 3.87 47.655 ;
      POLYGON 113.35 42.215 113.35 39.385 112.51 39.385 112.51 40.61 112.05 40.61 112.05 42.215 ;
      RECT -0.19 39.385 3.87 42.215 ;
      RECT 112.51 33.945 113.35 36.775 ;
      RECT -0.19 33.945 3.87 36.775 ;
      RECT 112.05 28.505 113.35 31.335 ;
      RECT -0.19 28.505 3.87 31.335 ;
      POLYGON 84.83 25.895 84.83 23.065 83.99 23.065 83.99 24.29 83.53 24.29 83.53 25.895 ;
      RECT -0.19 23.065 3.87 25.895 ;
      POLYGON 84.83 20.455 84.83 17.625 83.99 17.625 83.99 18.85 83.53 18.85 83.53 20.455 ;
      RECT -0.19 17.625 3.87 20.455 ;
      POLYGON 84.83 15.015 84.83 12.185 80.77 12.185 80.77 13.79 83.99 13.79 83.99 15.015 ;
      RECT -0.19 12.185 3.87 15.015 ;
      POLYGON 84.83 9.575 84.83 6.745 83.53 6.745 83.53 8.35 83.99 8.35 83.99 9.575 ;
      RECT -0.19 6.745 3.87 9.575 ;
      POLYGON 84.83 4.135 84.83 1.305 80.77 1.305 80.77 2.91 83.99 2.91 83.99 4.135 ;
      RECT -0.19 1.305 3.87 4.135 ;
      POLYGON 113.16 103.36 113.16 27.2 84.64 27.2 84.64 0 0 0 0 103.36 ;
    LAYER pwell ;
      RECT 106.85 103.31 107.07 103.48 ;
      RECT 103.17 103.31 103.39 103.48 ;
      RECT 99.49 103.31 99.71 103.48 ;
      RECT 95.81 103.31 96.03 103.48 ;
      RECT 92.13 103.31 92.35 103.48 ;
      RECT 88.45 103.31 88.67 103.48 ;
      RECT 84.77 103.31 84.99 103.48 ;
      RECT 81.09 103.31 81.31 103.48 ;
      RECT 77.41 103.31 77.63 103.48 ;
      RECT 73.73 103.31 73.95 103.48 ;
      RECT 70.05 103.31 70.27 103.48 ;
      RECT 66.37 103.31 66.59 103.48 ;
      RECT 62.69 103.31 62.91 103.48 ;
      RECT 59.01 103.31 59.23 103.48 ;
      RECT 55.33 103.31 55.55 103.48 ;
      RECT 51.65 103.31 51.87 103.48 ;
      RECT 47.97 103.31 48.19 103.48 ;
      RECT 44.29 103.31 44.51 103.48 ;
      RECT 40.61 103.31 40.83 103.48 ;
      RECT 36.93 103.31 37.15 103.48 ;
      RECT 33.25 103.31 33.47 103.48 ;
      RECT 29.57 103.31 29.79 103.48 ;
      RECT 25.89 103.31 26.11 103.48 ;
      RECT 22.21 103.31 22.43 103.48 ;
      RECT 18.53 103.31 18.75 103.48 ;
      RECT 14.85 103.31 15.07 103.48 ;
      RECT 11.17 103.31 11.39 103.48 ;
      RECT 7.49 103.31 7.71 103.48 ;
      RECT 3.81 103.31 4.03 103.48 ;
      RECT 0.13 103.31 0.35 103.48 ;
      RECT 110.575 103.3 110.685 103.42 ;
      RECT 112.395 103.3 112.555 103.41 ;
      RECT 112.395 27.15 112.555 27.26 ;
      RECT 110.575 27.14 110.685 27.26 ;
      RECT 106.85 27.08 107.07 27.25 ;
      RECT 103.17 27.08 103.39 27.25 ;
      RECT 99.49 27.08 99.71 27.25 ;
      RECT 95.81 27.08 96.03 27.25 ;
      RECT 92.13 27.08 92.35 27.25 ;
      RECT 88.45 27.08 88.67 27.25 ;
      RECT 84.77 27.08 84.99 27.25 ;
      RECT 81.09 -0.12 81.31 0.05 ;
      RECT 77.41 -0.12 77.63 0.05 ;
      RECT 73.73 -0.12 73.95 0.05 ;
      RECT 70.05 -0.12 70.27 0.05 ;
      RECT 66.37 -0.12 66.59 0.05 ;
      RECT 62.69 -0.12 62.91 0.05 ;
      RECT 59.01 -0.12 59.23 0.05 ;
      RECT 55.33 -0.12 55.55 0.05 ;
      RECT 51.65 -0.12 51.87 0.05 ;
      RECT 47.97 -0.12 48.19 0.05 ;
      RECT 44.29 -0.12 44.51 0.05 ;
      RECT 40.61 -0.12 40.83 0.05 ;
      RECT 36.93 -0.12 37.15 0.05 ;
      RECT 33.25 -0.12 33.47 0.05 ;
      RECT 29.57 -0.12 29.79 0.05 ;
      RECT 25.89 -0.12 26.11 0.05 ;
      RECT 22.21 -0.12 22.43 0.05 ;
      RECT 18.53 -0.12 18.75 0.05 ;
      RECT 14.85 -0.12 15.07 0.05 ;
      RECT 11.17 -0.12 11.39 0.05 ;
      RECT 7.49 -0.12 7.71 0.05 ;
      RECT 3.81 -0.12 4.03 0.05 ;
      RECT 0.13 -0.12 0.35 0.05 ;
      POLYGON 113.16 103.36 113.16 27.2 84.64 27.2 84.64 0 0 0 0 103.36 ;
    LAYER OVERLAP ;
      POLYGON 0 0 0 103.36 113.16 103.36 113.16 27.2 84.64 27.2 84.64 0 ;
  END
END sb_0__2_

END LIBRARY
