VERSION 5.7 ;
BUSBITCHARS "[]" ;

UNITS
  DATABASE MICRONS 1000 ;
END UNITS

MANUFACTURINGGRID 0.005 ;

LAYER li1
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.46 ;
  WIDTH 0.17 ;
END li1

LAYER mcon
  TYPE CUT ;
END mcon

LAYER met1
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.34 ;
  WIDTH 0.14 ;
END met1

LAYER via
  TYPE CUT ;
END via

LAYER met2
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.46 ;
  WIDTH 0.14 ;
END met2

LAYER via2
  TYPE CUT ;
END via2

LAYER met3
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.68 ;
  WIDTH 0.3 ;
END met3

LAYER via3
  TYPE CUT ;
END via3

LAYER met4
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.92 ;
  WIDTH 0.3 ;
END met4

LAYER via4
  TYPE CUT ;
END via4

LAYER met5
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 3.4 ;
  WIDTH 1.6 ;
END met5

LAYER nwell
  TYPE MASTERSLICE ;
END nwell

LAYER pwell
  TYPE MASTERSLICE ;
END pwell

LAYER OVERLAP
  TYPE OVERLAP ;
END OVERLAP

VIA L1M1_PR
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.145 -0.115 0.145 0.115 ;
END L1M1_PR

VIA L1M1_PR_R
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.115 -0.145 0.115 0.145 ;
END L1M1_PR_R

VIA L1M1_PR_M
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.115 -0.145 0.115 0.145 ;
END L1M1_PR_M

VIA L1M1_PR_MR
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.145 -0.115 0.145 0.115 ;
END L1M1_PR_MR

VIA L1M1_PR_C
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.145 -0.145 0.145 0.145 ;
END L1M1_PR_C

VIA M1M2_PR
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR

VIA M1M2_PR_Enc
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_Enc

VIA M1M2_PR_R
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_R

VIA M1M2_PR_R_Enc
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR_R_Enc

VIA M1M2_PR_M
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_M

VIA M1M2_PR_M_Enc
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR_M_Enc

VIA M1M2_PR_MR
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR_MR

VIA M1M2_PR_MR_Enc
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_MR_Enc

VIA M1M2_PR_C
  LAYER met1 ;
    RECT -0.16 -0.16 0.16 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.16 0.16 0.16 ;
END M1M2_PR_C

VIA M2M3_PR
  LAYER met2 ;
    RECT -0.14 -0.185 0.14 0.185 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR

VIA M2M3_PR_R
  LAYER met2 ;
    RECT -0.185 -0.14 0.185 0.14 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_R

VIA M2M3_PR_M
  LAYER met2 ;
    RECT -0.14 -0.185 0.14 0.185 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_M

VIA M2M3_PR_MR
  LAYER met2 ;
    RECT -0.185 -0.14 0.185 0.14 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_MR

VIA M2M3_PR_C
  LAYER met2 ;
    RECT -0.185 -0.185 0.185 0.185 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_C

VIA M3M4_PR
  LAYER met3 ;
    RECT -0.19 -0.16 0.19 0.16 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR

VIA M3M4_PR_R
  LAYER met3 ;
    RECT -0.16 -0.19 0.16 0.19 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_R

VIA M3M4_PR_M
  LAYER met3 ;
    RECT -0.19 -0.16 0.19 0.16 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_M

VIA M3M4_PR_MR
  LAYER met3 ;
    RECT -0.16 -0.19 0.16 0.19 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_MR

VIA M3M4_PR_C
  LAYER met3 ;
    RECT -0.19 -0.19 0.19 0.19 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_C

VIA M4M5_PR
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR

VIA M4M5_PR_R
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_R

VIA M4M5_PR_M
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_M

VIA M4M5_PR_MR
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_MR

VIA M4M5_PR_C
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_C

SITE unit
  CLASS CORE ;
  SYMMETRY Y ;
  SIZE 0.46 BY 2.72 ;
END unit

SITE unithddbl
  CLASS CORE ;
  SIZE 0.46 BY 5.44 ;
END unithddbl

MACRO cby_0__1_
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  SIZE 66.24 BY 76.16 ;
  SYMMETRY X Y ;
  PIN chany_bottom_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.72 0 62.86 0.485 ;
    END
  END chany_bottom_in[0]
  PIN chany_bottom_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.18 0 40.32 0.485 ;
    END
  END chany_bottom_in[1]
  PIN chany_bottom_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.68 0 51.82 0.485 ;
    END
  END chany_bottom_in[2]
  PIN chany_bottom_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.28 0 56.42 0.485 ;
    END
  END chany_bottom_in[3]
  PIN chany_bottom_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.52 0 53.66 0.485 ;
    END
  END chany_bottom_in[4]
  PIN chany_bottom_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.66 0 34.8 0.485 ;
    END
  END chany_bottom_in[5]
  PIN chany_bottom_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.96 0 14.1 0.485 ;
    END
  END chany_bottom_in[6]
  PIN chany_bottom_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.72 0 16.86 0.485 ;
    END
  END chany_bottom_in[7]
  PIN chany_bottom_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.26 0 39.4 0.485 ;
    END
  END chany_bottom_in[8]
  PIN chany_bottom_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.58 0 35.72 0.485 ;
    END
  END chany_bottom_in[9]
  PIN chany_bottom_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.8 0 61.94 0.485 ;
    END
  END chany_bottom_in[10]
  PIN chany_bottom_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.12 0 58.26 0.485 ;
    END
  END chany_bottom_in[11]
  PIN chany_bottom_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.74 0 33.88 0.485 ;
    END
  END chany_bottom_in[12]
  PIN chany_bottom_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.34 0 38.48 0.485 ;
    END
  END chany_bottom_in[13]
  PIN chany_bottom_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.88 0 15.02 0.485 ;
    END
  END chany_bottom_in[14]
  PIN chany_bottom_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.5 0 36.64 0.485 ;
    END
  END chany_bottom_in[15]
  PIN chany_bottom_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.96 0 60.1 0.485 ;
    END
  END chany_bottom_in[16]
  PIN chany_bottom_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.8 0 15.94 0.485 ;
    END
  END chany_bottom_in[17]
  PIN chany_bottom_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.42 0 37.56 0.485 ;
    END
  END chany_bottom_in[18]
  PIN chany_bottom_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.2 0 57.34 0.485 ;
    END
  END chany_bottom_in[19]
  PIN chany_top_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.76 75.675 50.9 76.16 ;
    END
  END chany_top_in[0]
  PIN chany_top_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.2 75.675 57.34 76.16 ;
    END
  END chany_top_in[1]
  PIN chany_top_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.1 75.675 41.24 76.16 ;
    END
  END chany_top_in[2]
  PIN chany_top_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.2 75.675 11.34 76.16 ;
    END
  END chany_top_in[3]
  PIN chany_top_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.74 75.675 33.88 76.16 ;
    END
  END chany_top_in[4]
  PIN chany_top_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.48 75.675 19.62 76.16 ;
    END
  END chany_top_in[5]
  PIN chany_top_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.12 75.675 12.26 76.16 ;
    END
  END chany_top_in[6]
  PIN chany_top_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.5 75.675 36.64 76.16 ;
    END
  END chany_top_in[7]
  PIN chany_top_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.56 75.675 18.7 76.16 ;
    END
  END chany_top_in[8]
  PIN chany_top_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.04 75.675 13.18 76.16 ;
    END
  END chany_top_in[9]
  PIN chany_top_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.04 75.675 59.18 76.16 ;
    END
  END chany_top_in[10]
  PIN chany_top_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.64 75.675 17.78 76.16 ;
    END
  END chany_top_in[11]
  PIN chany_top_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.28 75.675 10.42 76.16 ;
    END
  END chany_top_in[12]
  PIN chany_top_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.96 75.675 14.1 76.16 ;
    END
  END chany_top_in[13]
  PIN chany_top_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.42 75.675 37.56 76.16 ;
    END
  END chany_top_in[14]
  PIN chany_top_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.72 75.675 16.86 76.16 ;
    END
  END chany_top_in[15]
  PIN chany_top_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.44 75.675 54.58 76.16 ;
    END
  END chany_top_in[16]
  PIN chany_top_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.88 75.675 15.02 76.16 ;
    END
  END chany_top_in[17]
  PIN chany_top_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.46 75.675 2.6 76.16 ;
    END
  END chany_top_in[18]
  PIN chany_top_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.8 75.675 15.94 76.16 ;
    END
  END chany_top_in[19]
  PIN ccff_head[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.66 75.675 34.8 76.16 ;
    END
  END ccff_head[0]
  PIN chany_bottom_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48 0 48.14 0.485 ;
    END
  END chany_bottom_out[0]
  PIN chany_bottom_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.44 0 54.58 0.485 ;
    END
  END chany_bottom_out[1]
  PIN chany_bottom_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.08 0 47.22 0.485 ;
    END
  END chany_bottom_out[2]
  PIN chany_bottom_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.88 0 61.02 0.485 ;
    END
  END chany_bottom_out[3]
  PIN chany_bottom_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.76 0 50.9 0.485 ;
    END
  END chany_bottom_out[4]
  PIN chany_bottom_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.02 0 42.16 0.485 ;
    END
  END chany_bottom_out[5]
  PIN chany_bottom_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.9 0 32.04 0.485 ;
    END
  END chany_bottom_out[6]
  PIN chany_bottom_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.94 0 43.08 0.485 ;
    END
  END chany_bottom_out[7]
  PIN chany_bottom_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.04 0 13.18 0.485 ;
    END
  END chany_bottom_out[8]
  PIN chany_bottom_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.56 0 18.7 0.485 ;
    END
  END chany_bottom_out[9]
  PIN chany_bottom_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.84 0 49.98 0.485 ;
    END
  END chany_bottom_out[10]
  PIN chany_bottom_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.6 0 52.74 0.485 ;
    END
  END chany_bottom_out[11]
  PIN chany_bottom_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.04 0 59.18 0.485 ;
    END
  END chany_bottom_out[12]
  PIN chany_bottom_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.1 0 41.24 0.485 ;
    END
  END chany_bottom_out[13]
  PIN chany_bottom_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.82 0 32.96 0.485 ;
    END
  END chany_bottom_out[14]
  PIN chany_bottom_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.64 0 17.78 0.485 ;
    END
  END chany_bottom_out[15]
  PIN chany_bottom_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25 0 25.14 0.485 ;
    END
  END chany_bottom_out[16]
  PIN chany_bottom_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.98 0 31.12 0.485 ;
    END
  END chany_bottom_out[17]
  PIN chany_bottom_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.64 0 63.78 0.485 ;
    END
  END chany_bottom_out[18]
  PIN chany_bottom_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.92 0 49.06 0.485 ;
    END
  END chany_bottom_out[19]
  PIN chany_top_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.84 75.675 49.98 76.16 ;
    END
  END chany_top_out[0]
  PIN chany_top_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.96 75.675 60.1 76.16 ;
    END
  END chany_top_out[1]
  PIN chany_top_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.88 75.675 61.02 76.16 ;
    END
  END chany_top_out[2]
  PIN chany_top_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.64 75.675 63.78 76.16 ;
    END
  END chany_top_out[3]
  PIN chany_top_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.6 75.675 52.74 76.16 ;
    END
  END chany_top_out[4]
  PIN chany_top_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.26 75.675 39.4 76.16 ;
    END
  END chany_top_out[5]
  PIN chany_top_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.58 75.675 35.72 76.16 ;
    END
  END chany_top_out[6]
  PIN chany_top_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.72 75.675 62.86 76.16 ;
    END
  END chany_top_out[7]
  PIN chany_top_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.36 75.675 9.5 76.16 ;
    END
  END chany_top_out[8]
  PIN chany_top_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.44 75.675 8.58 76.16 ;
    END
  END chany_top_out[9]
  PIN chany_top_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.38 75.675 26.52 76.16 ;
    END
  END chany_top_out[10]
  PIN chany_top_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.68 75.675 51.82 76.16 ;
    END
  END chany_top_out[11]
  PIN chany_top_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.52 75.675 53.66 76.16 ;
    END
  END chany_top_out[12]
  PIN chany_top_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.28 75.675 56.42 76.16 ;
    END
  END chany_top_out[13]
  PIN chany_top_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.12 75.675 58.26 76.16 ;
    END
  END chany_top_out[14]
  PIN chany_top_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.34 75.675 38.48 76.16 ;
    END
  END chany_top_out[15]
  PIN chany_top_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.8 75.675 61.94 76.16 ;
    END
  END chany_top_out[16]
  PIN chany_top_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.82 75.675 32.96 76.16 ;
    END
  END chany_top_out[17]
  PIN chany_top_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.32 75.675 21.46 76.16 ;
    END
  END chany_top_out[18]
  PIN chany_top_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.18 75.675 40.32 76.16 ;
    END
  END chany_top_out[19]
  PIN left_grid_pin_0_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 20.59 0.8 20.89 ;
    END
  END left_grid_pin_0_[0]
  PIN ccff_tail[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 65.44 23.99 66.24 24.29 ;
    END
  END ccff_tail[0]
  PIN IO_ISOL_N[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 65.44 3.59 66.24 3.89 ;
    END
  END IO_ISOL_N[0]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 13.79 0.8 14.09 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN[0]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 8.35 0.8 8.65 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[0]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 9.71 0.8 10.01 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[0]
  PIN right_width_0_height_0__pin_0_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 21.95 0.8 22.25 ;
    END
  END right_width_0_height_0__pin_0_[0]
  PIN right_width_0_height_0__pin_1_upper[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.4 75.675 20.54 76.16 ;
    END
  END right_width_0_height_0__pin_1_upper[0]
  PIN right_width_0_height_0__pin_1_lower[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.38 0 26.52 0.485 ;
    END
  END right_width_0_height_0__pin_1_lower[0]
  PIN prog_clk_0_E_in
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER met3 ;
        RECT 65.44 10.39 66.24 10.69 ;
    END
  END prog_clk_0_E_in
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 0.48 2.96 ;
        RECT 65.76 2.48 66.24 2.96 ;
        RECT 0 7.92 0.48 8.4 ;
        RECT 65.76 7.92 66.24 8.4 ;
        RECT 0 13.36 0.48 13.84 ;
        RECT 65.76 13.36 66.24 13.84 ;
        RECT 0 18.8 0.48 19.28 ;
        RECT 65.76 18.8 66.24 19.28 ;
        RECT 0 24.24 0.48 24.72 ;
        RECT 65.76 24.24 66.24 24.72 ;
        RECT 0 29.68 0.48 30.16 ;
        RECT 65.76 29.68 66.24 30.16 ;
        RECT 0 35.12 0.48 35.6 ;
        RECT 65.76 35.12 66.24 35.6 ;
        RECT 0 40.56 0.48 41.04 ;
        RECT 65.76 40.56 66.24 41.04 ;
        RECT 0 46 0.48 46.48 ;
        RECT 65.76 46 66.24 46.48 ;
        RECT 0 51.44 0.48 51.92 ;
        RECT 65.76 51.44 66.24 51.92 ;
        RECT 0 56.88 0.48 57.36 ;
        RECT 65.76 56.88 66.24 57.36 ;
        RECT 0 62.32 0.48 62.8 ;
        RECT 65.76 62.32 66.24 62.8 ;
        RECT 0 67.76 0.48 68.24 ;
        RECT 65.76 67.76 66.24 68.24 ;
        RECT 0 73.2 0.48 73.68 ;
        RECT 65.76 73.2 66.24 73.68 ;
      LAYER met4 ;
        RECT 10.74 0 11.34 0.6 ;
        RECT 40.18 0 40.78 0.6 ;
        RECT 10.74 75.56 11.34 76.16 ;
        RECT 40.18 75.56 40.78 76.16 ;
      LAYER met5 ;
        RECT 0 5.88 3.2 9.08 ;
        RECT 63.04 5.88 66.24 9.08 ;
        RECT 0 46.68 3.2 49.88 ;
        RECT 63.04 46.68 66.24 49.88 ;
    END
  END VDD
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 0 45.4 0.24 ;
        RECT 46.6 0 66.24 0.24 ;
        RECT 0 5.2 0.48 5.68 ;
        RECT 65.76 5.2 66.24 5.68 ;
        RECT 0 10.64 0.48 11.12 ;
        RECT 65.76 10.64 66.24 11.12 ;
        RECT 0 16.08 0.48 16.56 ;
        RECT 65.76 16.08 66.24 16.56 ;
        RECT 0 21.52 0.48 22 ;
        RECT 65.76 21.52 66.24 22 ;
        RECT 0 26.96 0.48 27.44 ;
        RECT 65.76 26.96 66.24 27.44 ;
        RECT 0 32.4 0.48 32.88 ;
        RECT 65.76 32.4 66.24 32.88 ;
        RECT 0 37.84 0.48 38.32 ;
        RECT 65.76 37.84 66.24 38.32 ;
        RECT 0 43.28 0.48 43.76 ;
        RECT 65.76 43.28 66.24 43.76 ;
        RECT 0 48.72 0.48 49.2 ;
        RECT 65.76 48.72 66.24 49.2 ;
        RECT 0 54.16 0.48 54.64 ;
        RECT 65.76 54.16 66.24 54.64 ;
        RECT 0 59.6 0.48 60.08 ;
        RECT 65.76 59.6 66.24 60.08 ;
        RECT 0 65.04 0.48 65.52 ;
        RECT 65.76 65.04 66.24 65.52 ;
        RECT 0 70.48 0.48 70.96 ;
        RECT 65.76 70.48 66.24 70.96 ;
        RECT 0 75.92 45.4 76.16 ;
        RECT 46.6 75.92 66.24 76.16 ;
      LAYER met4 ;
        RECT 25.46 0 26.06 0.6 ;
        RECT 54.9 0 55.5 0.6 ;
        RECT 25.46 75.56 26.06 76.16 ;
        RECT 54.9 75.56 55.5 76.16 ;
      LAYER met5 ;
        RECT 0 26.28 3.2 29.48 ;
        RECT 63.04 26.28 66.24 29.48 ;
        RECT 0 67.08 3.2 70.28 ;
        RECT 63.04 67.08 66.24 70.28 ;
    END
  END VSS
  OBS
    LAYER met2 ;
      RECT 55.06 75.975 55.34 76.345 ;
      RECT 25.62 75.975 25.9 76.345 ;
      POLYGON 39.9 76.06 39.9 75.92 39.86 75.92 39.86 71.84 39.72 71.84 39.72 76.06 ;
      POLYGON 11.8 76.06 11.8 47.7 11.66 47.7 11.66 75.92 11.62 75.92 11.62 76.06 ;
      RECT 36.9 75.15 37.16 75.47 ;
      POLYGON 39.86 6.7 39.86 0.24 39.9 0.24 39.9 0.1 39.72 0.1 39.72 6.7 ;
      RECT 55.06 -0.185 55.34 0.185 ;
      RECT 25.62 -0.185 25.9 0.185 ;
      POLYGON 65.96 75.88 65.96 0.28 64.06 0.28 64.06 0.765 63.36 0.765 63.36 0.28 63.14 0.28 63.14 0.765 62.44 0.765 62.44 0.28 62.22 0.28 62.22 0.765 61.52 0.765 61.52 0.28 61.3 0.28 61.3 0.765 60.6 0.765 60.6 0.28 60.38 0.28 60.38 0.765 59.68 0.765 59.68 0.28 59.46 0.28 59.46 0.765 58.76 0.765 58.76 0.28 58.54 0.28 58.54 0.765 57.84 0.765 57.84 0.28 57.62 0.28 57.62 0.765 56.92 0.765 56.92 0.28 56.7 0.28 56.7 0.765 56 0.765 56 0.28 54.86 0.28 54.86 0.765 54.16 0.765 54.16 0.28 53.94 0.28 53.94 0.765 53.24 0.765 53.24 0.28 53.02 0.28 53.02 0.765 52.32 0.765 52.32 0.28 52.1 0.28 52.1 0.765 51.4 0.765 51.4 0.28 51.18 0.28 51.18 0.765 50.48 0.765 50.48 0.28 50.26 0.28 50.26 0.765 49.56 0.765 49.56 0.28 49.34 0.28 49.34 0.765 48.64 0.765 48.64 0.28 48.42 0.28 48.42 0.765 47.72 0.765 47.72 0.28 47.5 0.28 47.5 0.765 46.8 0.765 46.8 0.28 43.36 0.28 43.36 0.765 42.66 0.765 42.66 0.28 42.44 0.28 42.44 0.765 41.74 0.765 41.74 0.28 41.52 0.28 41.52 0.765 40.82 0.765 40.82 0.28 40.6 0.28 40.6 0.765 39.9 0.765 39.9 0.28 39.68 0.28 39.68 0.765 38.98 0.765 38.98 0.28 38.76 0.28 38.76 0.765 38.06 0.765 38.06 0.28 37.84 0.28 37.84 0.765 37.14 0.765 37.14 0.28 36.92 0.28 36.92 0.765 36.22 0.765 36.22 0.28 36 0.28 36 0.765 35.3 0.765 35.3 0.28 35.08 0.28 35.08 0.765 34.38 0.765 34.38 0.28 34.16 0.28 34.16 0.765 33.46 0.765 33.46 0.28 33.24 0.28 33.24 0.765 32.54 0.765 32.54 0.28 32.32 0.28 32.32 0.765 31.62 0.765 31.62 0.28 31.4 0.28 31.4 0.765 30.7 0.765 30.7 0.28 26.8 0.28 26.8 0.765 26.1 0.765 26.1 0.28 25.42 0.28 25.42 0.765 24.72 0.765 24.72 0.28 18.98 0.28 18.98 0.765 18.28 0.765 18.28 0.28 18.06 0.28 18.06 0.765 17.36 0.765 17.36 0.28 17.14 0.28 17.14 0.765 16.44 0.765 16.44 0.28 16.22 0.28 16.22 0.765 15.52 0.765 15.52 0.28 15.3 0.28 15.3 0.765 14.6 0.765 14.6 0.28 14.38 0.28 14.38 0.765 13.68 0.765 13.68 0.28 13.46 0.28 13.46 0.765 12.76 0.765 12.76 0.28 0.28 0.28 0.28 75.88 2.18 75.88 2.18 75.395 2.88 75.395 2.88 75.88 8.16 75.88 8.16 75.395 8.86 75.395 8.86 75.88 9.08 75.88 9.08 75.395 9.78 75.395 9.78 75.88 10 75.88 10 75.395 10.7 75.395 10.7 75.88 10.92 75.88 10.92 75.395 11.62 75.395 11.62 75.88 11.84 75.88 11.84 75.395 12.54 75.395 12.54 75.88 12.76 75.88 12.76 75.395 13.46 75.395 13.46 75.88 13.68 75.88 13.68 75.395 14.38 75.395 14.38 75.88 14.6 75.88 14.6 75.395 15.3 75.395 15.3 75.88 15.52 75.88 15.52 75.395 16.22 75.395 16.22 75.88 16.44 75.88 16.44 75.395 17.14 75.395 17.14 75.88 17.36 75.88 17.36 75.395 18.06 75.395 18.06 75.88 18.28 75.88 18.28 75.395 18.98 75.395 18.98 75.88 19.2 75.88 19.2 75.395 19.9 75.395 19.9 75.88 20.12 75.88 20.12 75.395 20.82 75.395 20.82 75.88 21.04 75.88 21.04 75.395 21.74 75.395 21.74 75.88 26.1 75.88 26.1 75.395 26.8 75.395 26.8 75.88 32.54 75.88 32.54 75.395 33.24 75.395 33.24 75.88 33.46 75.88 33.46 75.395 34.16 75.395 34.16 75.88 34.38 75.88 34.38 75.395 35.08 75.395 35.08 75.88 35.3 75.88 35.3 75.395 36 75.395 36 75.88 36.22 75.88 36.22 75.395 36.92 75.395 36.92 75.88 37.14 75.88 37.14 75.395 37.84 75.395 37.84 75.88 38.06 75.88 38.06 75.395 38.76 75.395 38.76 75.88 38.98 75.88 38.98 75.395 39.68 75.395 39.68 75.88 39.9 75.88 39.9 75.395 40.6 75.395 40.6 75.88 40.82 75.88 40.82 75.395 41.52 75.395 41.52 75.88 49.56 75.88 49.56 75.395 50.26 75.395 50.26 75.88 50.48 75.88 50.48 75.395 51.18 75.395 51.18 75.88 51.4 75.88 51.4 75.395 52.1 75.395 52.1 75.88 52.32 75.88 52.32 75.395 53.02 75.395 53.02 75.88 53.24 75.88 53.24 75.395 53.94 75.395 53.94 75.88 54.16 75.88 54.16 75.395 54.86 75.395 54.86 75.88 56 75.88 56 75.395 56.7 75.395 56.7 75.88 56.92 75.88 56.92 75.395 57.62 75.395 57.62 75.88 57.84 75.88 57.84 75.395 58.54 75.395 58.54 75.88 58.76 75.88 58.76 75.395 59.46 75.395 59.46 75.88 59.68 75.88 59.68 75.395 60.38 75.395 60.38 75.88 60.6 75.88 60.6 75.395 61.3 75.395 61.3 75.88 61.52 75.88 61.52 75.395 62.22 75.395 62.22 75.88 62.44 75.88 62.44 75.395 63.14 75.395 63.14 75.88 63.36 75.88 63.36 75.395 64.06 75.395 64.06 75.88 ;
    LAYER met3 ;
      POLYGON 55.365 76.325 55.365 76.32 55.58 76.32 55.58 76 55.365 76 55.365 75.995 55.035 75.995 55.035 76 54.82 76 54.82 76.32 55.035 76.32 55.035 76.325 ;
      POLYGON 25.925 76.325 25.925 76.32 26.14 76.32 26.14 76 25.925 76 25.925 75.995 25.595 75.995 25.595 76 25.38 76 25.38 76.32 25.595 76.32 25.595 76.325 ;
      POLYGON 55.365 0.165 55.365 0.16 55.58 0.16 55.58 -0.16 55.365 -0.16 55.365 -0.165 55.035 -0.165 55.035 -0.16 54.82 -0.16 54.82 0.16 55.035 0.16 55.035 0.165 ;
      POLYGON 25.925 0.165 25.925 0.16 26.14 0.16 26.14 -0.16 25.925 -0.16 25.925 -0.165 25.595 -0.165 25.595 -0.16 25.38 -0.16 25.38 0.16 25.595 0.16 25.595 0.165 ;
      POLYGON 65.84 75.76 65.84 24.69 65.04 24.69 65.04 23.59 65.84 23.59 65.84 11.09 65.04 11.09 65.04 9.99 65.84 9.99 65.84 4.29 65.04 4.29 65.04 3.19 65.84 3.19 65.84 0.4 0.4 0.4 0.4 7.95 1.2 7.95 1.2 9.05 0.4 9.05 0.4 9.31 1.2 9.31 1.2 10.41 0.4 10.41 0.4 13.39 1.2 13.39 1.2 14.49 0.4 14.49 0.4 20.19 1.2 20.19 1.2 21.29 0.4 21.29 0.4 21.55 1.2 21.55 1.2 22.65 0.4 22.65 0.4 75.76 ;
    LAYER met5 ;
      POLYGON 64.64 74.56 64.64 71.88 61.44 71.88 61.44 65.48 64.64 65.48 64.64 51.48 61.44 51.48 61.44 45.08 64.64 45.08 64.64 31.08 61.44 31.08 61.44 24.68 64.64 24.68 64.64 10.68 61.44 10.68 61.44 4.28 64.64 4.28 64.64 1.6 1.6 1.6 1.6 4.28 4.8 4.28 4.8 10.68 1.6 10.68 1.6 24.68 4.8 24.68 4.8 31.08 1.6 31.08 1.6 45.08 4.8 45.08 4.8 51.48 1.6 51.48 1.6 65.48 4.8 65.48 4.8 71.88 1.6 71.88 1.6 74.56 ;
    LAYER met4 ;
      POLYGON 65.84 75.76 65.84 0.4 55.9 0.4 55.9 1 54.5 1 54.5 0.4 41.18 0.4 41.18 1 39.78 1 39.78 0.4 26.46 0.4 26.46 1 25.06 1 25.06 0.4 11.74 0.4 11.74 1 10.34 1 10.34 0.4 0.4 0.4 0.4 75.76 10.34 75.76 10.34 75.16 11.74 75.16 11.74 75.76 25.06 75.76 25.06 75.16 26.46 75.16 26.46 75.76 39.78 75.76 39.78 75.16 41.18 75.16 41.18 75.76 54.5 75.76 54.5 75.16 55.9 75.16 55.9 75.76 ;
    LAYER met1 ;
      RECT 45.68 75.92 46.32 76.4 ;
      RECT 45.68 -0.24 46.32 0.24 ;
      POLYGON 46.32 75.88 46.32 75.64 65.96 75.64 65.96 73.96 65.48 73.96 65.48 72.92 65.96 72.92 65.96 71.24 65.48 71.24 65.48 70.2 65.96 70.2 65.96 68.52 65.48 68.52 65.48 67.48 65.96 67.48 65.96 65.8 65.48 65.8 65.48 64.76 65.96 64.76 65.96 63.08 65.48 63.08 65.48 62.04 65.96 62.04 65.96 60.36 65.48 60.36 65.48 59.32 65.96 59.32 65.96 57.64 65.48 57.64 65.48 56.6 65.96 56.6 65.96 54.92 65.48 54.92 65.48 53.88 65.96 53.88 65.96 52.2 65.48 52.2 65.48 51.16 65.96 51.16 65.96 49.48 65.48 49.48 65.48 48.44 65.96 48.44 65.96 46.76 65.48 46.76 65.48 45.72 65.96 45.72 65.96 44.04 65.48 44.04 65.48 43 65.96 43 65.96 41.32 65.48 41.32 65.48 40.28 65.96 40.28 65.96 38.6 65.48 38.6 65.48 37.56 65.96 37.56 65.96 35.88 65.48 35.88 65.48 34.84 65.96 34.84 65.96 33.16 65.48 33.16 65.48 32.12 65.96 32.12 65.96 30.44 65.48 30.44 65.48 29.4 65.96 29.4 65.96 27.72 65.48 27.72 65.48 26.68 65.96 26.68 65.96 25 65.48 25 65.48 23.96 65.96 23.96 65.96 22.28 65.48 22.28 65.48 21.24 65.96 21.24 65.96 19.56 65.48 19.56 65.48 18.52 65.96 18.52 65.96 16.84 65.48 16.84 65.48 15.8 65.96 15.8 65.96 14.12 65.48 14.12 65.48 13.08 65.96 13.08 65.96 11.4 65.48 11.4 65.48 10.36 65.96 10.36 65.96 8.68 65.48 8.68 65.48 7.64 65.96 7.64 65.96 5.96 65.48 5.96 65.48 4.92 65.96 4.92 65.96 3.24 65.48 3.24 65.48 2.2 65.96 2.2 65.96 0.52 46.32 0.52 46.32 0.28 45.68 0.28 45.68 0.52 0.28 0.52 0.28 2.2 0.76 2.2 0.76 3.24 0.28 3.24 0.28 4.92 0.76 4.92 0.76 5.96 0.28 5.96 0.28 7.64 0.76 7.64 0.76 8.68 0.28 8.68 0.28 10.36 0.76 10.36 0.76 11.4 0.28 11.4 0.28 13.08 0.76 13.08 0.76 14.12 0.28 14.12 0.28 15.8 0.76 15.8 0.76 16.84 0.28 16.84 0.28 18.52 0.76 18.52 0.76 19.56 0.28 19.56 0.28 21.24 0.76 21.24 0.76 22.28 0.28 22.28 0.28 23.96 0.76 23.96 0.76 25 0.28 25 0.28 26.68 0.76 26.68 0.76 27.72 0.28 27.72 0.28 29.4 0.76 29.4 0.76 30.44 0.28 30.44 0.28 32.12 0.76 32.12 0.76 33.16 0.28 33.16 0.28 34.84 0.76 34.84 0.76 35.88 0.28 35.88 0.28 37.56 0.76 37.56 0.76 38.6 0.28 38.6 0.28 40.28 0.76 40.28 0.76 41.32 0.28 41.32 0.28 43 0.76 43 0.76 44.04 0.28 44.04 0.28 45.72 0.76 45.72 0.76 46.76 0.28 46.76 0.28 48.44 0.76 48.44 0.76 49.48 0.28 49.48 0.28 51.16 0.76 51.16 0.76 52.2 0.28 52.2 0.28 53.88 0.76 53.88 0.76 54.92 0.28 54.92 0.28 56.6 0.76 56.6 0.76 57.64 0.28 57.64 0.28 59.32 0.76 59.32 0.76 60.36 0.28 60.36 0.28 62.04 0.76 62.04 0.76 63.08 0.28 63.08 0.28 64.76 0.76 64.76 0.76 65.8 0.28 65.8 0.28 67.48 0.76 67.48 0.76 68.52 0.28 68.52 0.28 70.2 0.76 70.2 0.76 71.24 0.28 71.24 0.28 72.92 0.76 72.92 0.76 73.96 0.28 73.96 0.28 75.64 45.68 75.64 45.68 75.88 ;
    LAYER li1 ;
      POLYGON 66.24 76.245 66.24 76.075 59.715 76.075 59.715 75.35 59.425 75.35 59.425 76.075 52.355 76.075 52.355 75.35 52.065 75.35 52.065 76.075 37.635 76.075 37.635 75.35 37.345 75.35 37.345 76.075 22.455 76.075 22.455 75.35 22.165 75.35 22.165 76.075 16.005 76.075 16.005 75.275 15.675 75.275 15.675 76.075 15.165 76.075 15.165 75.595 14.835 75.595 14.835 76.075 14.325 76.075 14.325 75.595 13.995 75.595 13.995 76.075 13.405 76.075 13.405 75.595 13.235 75.595 13.235 76.075 12.565 76.075 12.565 75.595 12.395 75.595 12.395 76.075 7.735 76.075 7.735 75.35 7.445 75.35 7.445 76.075 0 76.075 0 76.245 ;
      RECT 65.32 73.355 66.24 73.525 ;
      RECT 0 73.355 3.68 73.525 ;
      RECT 65.32 70.635 66.24 70.805 ;
      RECT 0 70.635 3.68 70.805 ;
      RECT 65.32 67.915 66.24 68.085 ;
      RECT 0 67.915 3.68 68.085 ;
      RECT 65.32 65.195 66.24 65.365 ;
      RECT 0 65.195 3.68 65.365 ;
      RECT 65.32 62.475 66.24 62.645 ;
      RECT 0 62.475 3.68 62.645 ;
      RECT 65.32 59.755 66.24 59.925 ;
      RECT 0 59.755 3.68 59.925 ;
      RECT 65.32 57.035 66.24 57.205 ;
      RECT 0 57.035 3.68 57.205 ;
      RECT 65.32 54.315 66.24 54.485 ;
      RECT 0 54.315 3.68 54.485 ;
      RECT 65.32 51.595 66.24 51.765 ;
      RECT 0 51.595 3.68 51.765 ;
      RECT 65.32 48.875 66.24 49.045 ;
      RECT 0 48.875 3.68 49.045 ;
      RECT 65.32 46.155 66.24 46.325 ;
      RECT 0 46.155 3.68 46.325 ;
      RECT 65.32 43.435 66.24 43.605 ;
      RECT 0 43.435 3.68 43.605 ;
      RECT 65.32 40.715 66.24 40.885 ;
      RECT 0 40.715 3.68 40.885 ;
      RECT 65.32 37.995 66.24 38.165 ;
      RECT 0 37.995 3.68 38.165 ;
      RECT 65.32 35.275 66.24 35.445 ;
      RECT 0 35.275 3.68 35.445 ;
      RECT 65.32 32.555 66.24 32.725 ;
      RECT 0 32.555 3.68 32.725 ;
      RECT 65.32 29.835 66.24 30.005 ;
      RECT 0 29.835 3.68 30.005 ;
      RECT 65.32 27.115 66.24 27.285 ;
      RECT 0 27.115 3.68 27.285 ;
      RECT 65.32 24.395 66.24 24.565 ;
      RECT 0 24.395 3.68 24.565 ;
      RECT 65.32 21.675 66.24 21.845 ;
      RECT 0 21.675 3.68 21.845 ;
      RECT 65.32 18.955 66.24 19.125 ;
      RECT 0 18.955 3.68 19.125 ;
      RECT 65.32 16.235 66.24 16.405 ;
      RECT 0 16.235 3.68 16.405 ;
      RECT 65.32 13.515 66.24 13.685 ;
      RECT 0 13.515 3.68 13.685 ;
      RECT 65.32 10.795 66.24 10.965 ;
      RECT 0 10.795 3.68 10.965 ;
      RECT 65.32 8.075 66.24 8.245 ;
      RECT 0 8.075 3.68 8.245 ;
      RECT 65.32 5.355 66.24 5.525 ;
      RECT 0 5.355 3.68 5.525 ;
      RECT 65.32 2.635 66.24 2.805 ;
      RECT 0 2.635 3.68 2.805 ;
      POLYGON 57.865 0.885 57.865 0.085 59.425 0.085 59.425 0.81 59.715 0.81 59.715 0.085 66.24 0.085 66.24 -0.085 0 -0.085 0 0.085 7.445 0.085 7.445 0.81 7.735 0.81 7.735 0.085 22.165 0.085 22.165 0.81 22.455 0.81 22.455 0.085 22.975 0.085 22.975 0.565 23.145 0.565 23.145 0.085 23.815 0.085 23.815 0.565 23.985 0.565 23.985 0.085 24.575 0.085 24.575 0.565 24.905 0.565 24.905 0.085 25.415 0.085 25.415 0.565 25.745 0.565 25.745 0.085 26.255 0.085 26.255 0.885 26.585 0.885 26.585 0.085 31.715 0.085 31.715 0.565 31.885 0.565 31.885 0.085 32.555 0.085 32.555 0.565 32.725 0.565 32.725 0.085 33.315 0.085 33.315 0.565 33.645 0.565 33.645 0.085 34.155 0.085 34.155 0.565 34.485 0.565 34.485 0.085 34.995 0.085 34.995 0.885 35.325 0.885 35.325 0.085 37.345 0.085 37.345 0.81 37.635 0.81 37.635 0.085 38.155 0.085 38.155 0.565 38.325 0.565 38.325 0.085 38.995 0.085 38.995 0.565 39.165 0.565 39.165 0.085 39.755 0.085 39.755 0.565 40.085 0.565 40.085 0.085 40.595 0.085 40.595 0.565 40.925 0.565 40.925 0.085 41.435 0.085 41.435 0.885 41.765 0.885 41.765 0.085 46.935 0.085 46.935 0.885 47.265 0.885 47.265 0.085 47.775 0.085 47.775 0.565 48.105 0.565 48.105 0.085 48.615 0.085 48.615 0.565 48.945 0.565 48.945 0.085 49.455 0.085 49.455 0.565 49.785 0.565 49.785 0.085 50.295 0.085 50.295 0.565 50.625 0.565 50.625 0.085 51.135 0.085 51.135 0.565 51.465 0.565 51.465 0.085 52.065 0.085 52.065 0.81 52.355 0.81 52.355 0.085 54.255 0.085 54.255 0.565 54.425 0.565 54.425 0.085 55.095 0.085 55.095 0.565 55.265 0.565 55.265 0.085 55.855 0.085 55.855 0.565 56.185 0.565 56.185 0.085 56.695 0.085 56.695 0.565 57.025 0.565 57.025 0.085 57.535 0.085 57.535 0.885 ;
      RECT 0.17 0.17 66.07 75.99 ;
    LAYER via ;
      RECT 55.125 76.085 55.275 76.235 ;
      RECT 25.685 76.085 25.835 76.235 ;
      RECT 55.125 -0.075 55.275 0.075 ;
      RECT 25.685 -0.075 25.835 0.075 ;
    LAYER via2 ;
      RECT 55.1 76.06 55.3 76.26 ;
      RECT 25.66 76.06 25.86 76.26 ;
      RECT 55.1 -0.1 55.3 0.1 ;
      RECT 25.66 -0.1 25.86 0.1 ;
    LAYER via3 ;
      RECT 55.1 76.06 55.3 76.26 ;
      RECT 25.66 76.06 25.86 76.26 ;
      RECT 55.1 -0.1 55.3 0.1 ;
      RECT 25.66 -0.1 25.86 0.1 ;
    LAYER OVERLAP ;
      POLYGON 0 0 0 76.16 66.24 76.16 66.24 0 ;
  END
END cby_0__1_

END LIBRARY
