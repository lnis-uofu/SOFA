VERSION 5.7 ;
BUSBITCHARS "[]" ;

UNITS
  DATABASE MICRONS 1000 ;
END UNITS

MANUFACTURINGGRID 0.005 ;

LAYER nwell
  TYPE MASTERSLICE ;
END nwell

LAYER pwell
  TYPE MASTERSLICE ;
END pwell

LAYER fieldpoly
  TYPE MASTERSLICE ;
END fieldpoly

LAYER li1
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.46 ;
  WIDTH 0.17 ;
END li1

LAYER mcon
  TYPE CUT ;
END mcon

LAYER met1
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.34 ;
  WIDTH 0.14 ;
END met1

LAYER via
  TYPE CUT ;
END via

LAYER met2
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.46 ;
  WIDTH 0.14 ;
END met2

LAYER via2
  TYPE CUT ;
END via2

LAYER met3
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.68 ;
  WIDTH 0.3 ;
END met3

LAYER via3
  TYPE CUT ;
END via3

LAYER met4
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.92 ;
  WIDTH 0.3 ;
END met4

LAYER via4
  TYPE CUT ;
END via4

LAYER met5
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 3.4 ;
  WIDTH 1.6 ;
END met5

LAYER diff
  TYPE MASTERSLICE ;
END diff

LAYER licon1
  TYPE MASTERSLICE ;
END licon1

LAYER OVERLAP
  TYPE OVERLAP ;
END OVERLAP

VIA L1M1_PR
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.145 -0.115 0.145 0.115 ;
END L1M1_PR

VIA L1M1_PR_R
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.115 -0.145 0.115 0.145 ;
END L1M1_PR_R

VIA L1M1_PR_M
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.115 -0.145 0.115 0.145 ;
END L1M1_PR_M

VIA L1M1_PR_MR
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.145 -0.115 0.145 0.115 ;
END L1M1_PR_MR

VIA L1M1_PR_C
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.145 -0.145 0.145 0.145 ;
END L1M1_PR_C

VIA M1M2_PR
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR

VIA M1M2_PR_Enc
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_Enc

VIA M1M2_PR_R
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_R

VIA M1M2_PR_R_Enc
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR_R_Enc

VIA M1M2_PR_M
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_M

VIA M1M2_PR_M_Enc
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR_M_Enc

VIA M1M2_PR_MR
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR_MR

VIA M1M2_PR_MR_Enc
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_MR_Enc

VIA M1M2_PR_C
  LAYER met1 ;
    RECT -0.16 -0.16 0.16 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.16 0.16 0.16 ;
END M1M2_PR_C

VIA M2M3_PR
  LAYER met2 ;
    RECT -0.14 -0.185 0.14 0.185 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR

VIA M2M3_PR_R
  LAYER met2 ;
    RECT -0.185 -0.14 0.185 0.14 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_R

VIA M2M3_PR_M
  LAYER met2 ;
    RECT -0.14 -0.185 0.14 0.185 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_M

VIA M2M3_PR_MR
  LAYER met2 ;
    RECT -0.185 -0.14 0.185 0.14 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_MR

VIA M2M3_PR_C
  LAYER met2 ;
    RECT -0.185 -0.185 0.185 0.185 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_C

VIA M3M4_PR
  LAYER met3 ;
    RECT -0.19 -0.16 0.19 0.16 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR

VIA M3M4_PR_R
  LAYER met3 ;
    RECT -0.16 -0.19 0.16 0.19 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_R

VIA M3M4_PR_M
  LAYER met3 ;
    RECT -0.19 -0.16 0.19 0.16 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_M

VIA M3M4_PR_MR
  LAYER met3 ;
    RECT -0.16 -0.19 0.16 0.19 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_MR

VIA M3M4_PR_C
  LAYER met3 ;
    RECT -0.19 -0.19 0.19 0.19 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_C

VIA M4M5_PR
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR

VIA M4M5_PR_R
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_R

VIA M4M5_PR_M
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_M

VIA M4M5_PR_MR
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_MR

VIA M4M5_PR_C
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_C

SITE unit
  CLASS CORE ;
  SYMMETRY Y ;
  SIZE 0.46 BY 2.72 ;
END unit

SITE unithddbl
  CLASS CORE ;
  SIZE 0.46 BY 5.44 ;
END unithddbl

MACRO cby_0__1_
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  SIZE 84.64 BY 108.8 ;
  SYMMETRY X Y ;
  PIN prog_clk[0]
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER met3 ;
        RECT 0 3.25 1.38 3.55 ;
    END
  END prog_clk[0]
  PIN chany_bottom_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.71 0 42.85 1.36 ;
    END
  END chany_bottom_in[0]
  PIN chany_bottom_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.69 0 25.83 1.36 ;
    END
  END chany_bottom_in[1]
  PIN chany_bottom_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.23 0 71.37 1.36 ;
    END
  END chany_bottom_in[2]
  PIN chany_bottom_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.15 0 49.29 1.36 ;
    END
  END chany_bottom_in[3]
  PIN chany_bottom_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.27 0 36.41 1.36 ;
    END
  END chany_bottom_in[4]
  PIN chany_bottom_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.55 0 44.69 1.36 ;
    END
  END chany_bottom_in[5]
  PIN chany_bottom_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 5.37 0 5.67 1.36 ;
    END
  END chany_bottom_in[6]
  PIN chany_bottom_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 68.85 0 69.15 1.36 ;
    END
  END chany_bottom_in[7]
  PIN chany_bottom_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 21.93 0 22.23 1.36 ;
    END
  END chany_bottom_in[8]
  PIN chany_bottom_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 9.05 0 9.35 1.36 ;
    END
  END chany_bottom_in[9]
  PIN chany_bottom_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.39 0 46.53 1.36 ;
    END
  END chany_bottom_in[10]
  PIN chany_bottom_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.99 0 51.13 1.36 ;
    END
  END chany_bottom_in[11]
  PIN chany_bottom_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.29 0 7.43 1.36 ;
    END
  END chany_bottom_in[12]
  PIN chany_bottom_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 23.77 0 24.07 1.36 ;
    END
  END chany_bottom_in[13]
  PIN chany_bottom_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 7.21 0 7.51 1.36 ;
    END
  END chany_bottom_in[14]
  PIN chany_bottom_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 45.85 0 46.15 1.36 ;
    END
  END chany_bottom_in[15]
  PIN chany_bottom_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.23 0 48.37 1.36 ;
    END
  END chany_bottom_in[16]
  PIN chany_bottom_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.83 0 52.97 1.36 ;
    END
  END chany_bottom_in[17]
  PIN chany_bottom_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 47.69 0 47.99 1.36 ;
    END
  END chany_bottom_in[18]
  PIN chany_bottom_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 25.61 0 25.91 1.36 ;
    END
  END chany_bottom_in[19]
  PIN chany_top_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.07 107.44 50.21 108.8 ;
    END
  END chany_top_in[0]
  PIN chany_top_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.43 107.44 34.57 108.8 ;
    END
  END chany_top_in[1]
  PIN chany_top_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.63 107.44 66.77 108.8 ;
    END
  END chany_top_in[2]
  PIN chany_top_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.55 107.44 44.69 108.8 ;
    END
  END chany_top_in[3]
  PIN chany_top_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.99 107.44 51.13 108.8 ;
    END
  END chany_top_in[4]
  PIN chany_top_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.47 107.44 45.61 108.8 ;
    END
  END chany_top_in[5]
  PIN chany_top_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.31 107.44 70.45 108.8 ;
    END
  END chany_top_in[6]
  PIN chany_top_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.47 107.44 68.61 108.8 ;
    END
  END chany_top_in[7]
  PIN chany_top_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.39 107.44 69.53 108.8 ;
    END
  END chany_top_in[8]
  PIN chany_top_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.69 107.44 25.83 108.8 ;
    END
  END chany_top_in[9]
  PIN chany_top_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.71 107.44 42.85 108.8 ;
    END
  END chany_top_in[10]
  PIN chany_top_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.23 107.44 48.37 108.8 ;
    END
  END chany_top_in[11]
  PIN chany_top_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.55 107.44 67.69 108.8 ;
    END
  END chany_top_in[12]
  PIN chany_top_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 49.53 107.44 49.83 108.8 ;
    END
  END chany_top_in[13]
  PIN chany_top_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 45.85 107.44 46.15 108.8 ;
    END
  END chany_top_in[14]
  PIN chany_top_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 47.69 107.44 47.99 108.8 ;
    END
  END chany_top_in[15]
  PIN chany_top_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.45 107.44 28.59 108.8 ;
    END
  END chany_top_in[16]
  PIN chany_top_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.31 107.44 47.45 108.8 ;
    END
  END chany_top_in[17]
  PIN chany_top_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 23.77 107.44 24.07 108.8 ;
    END
  END chany_top_in[18]
  PIN chany_top_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 25.61 107.44 25.91 108.8 ;
    END
  END chany_top_in[19]
  PIN ccff_head[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.21 107.44 54.35 108.8 ;
    END
  END ccff_head[0]
  PIN chany_bottom_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.55 0 67.69 1.36 ;
    END
  END chany_bottom_out[0]
  PIN chany_bottom_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.03 0 62.17 1.36 ;
    END
  END chany_bottom_out[1]
  PIN chany_bottom_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.31 0 70.45 1.36 ;
    END
  END chany_bottom_out[2]
  PIN chany_bottom_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.47 0 45.61 1.36 ;
    END
  END chany_bottom_out[3]
  PIN chany_bottom_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.63 0 43.77 1.36 ;
    END
  END chany_bottom_out[4]
  PIN chany_bottom_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.91 0 29.05 1.36 ;
    END
  END chany_bottom_out[5]
  PIN chany_bottom_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.39 0 69.53 1.36 ;
    END
  END chany_bottom_out[6]
  PIN chany_bottom_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.47 0 68.61 1.36 ;
    END
  END chany_bottom_out[7]
  PIN chany_bottom_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.95 0 63.09 1.36 ;
    END
  END chany_bottom_out[8]
  PIN chany_bottom_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.91 0 52.05 1.36 ;
    END
  END chany_bottom_out[9]
  PIN chany_bottom_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.07 0 50.21 1.36 ;
    END
  END chany_bottom_out[10]
  PIN chany_bottom_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.79 0 41.93 1.36 ;
    END
  END chany_bottom_out[11]
  PIN chany_bottom_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.15 0 72.29 1.36 ;
    END
  END chany_bottom_out[12]
  PIN chany_bottom_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 20.09 0 20.39 1.36 ;
    END
  END chany_bottom_out[13]
  PIN chany_bottom_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 29.29 0 29.59 1.36 ;
    END
  END chany_bottom_out[14]
  PIN chany_bottom_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 49.53 0 49.83 1.36 ;
    END
  END chany_bottom_out[15]
  PIN chany_bottom_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 58.73 0 59.03 1.36 ;
    END
  END chany_bottom_out[16]
  PIN chany_bottom_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 14.57 0 14.87 1.36 ;
    END
  END chany_bottom_out[17]
  PIN chany_bottom_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 44.01 0 44.31 1.36 ;
    END
  END chany_bottom_out[18]
  PIN chany_bottom_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.31 0 47.45 1.36 ;
    END
  END chany_bottom_out[19]
  PIN chany_top_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.71 107.44 65.85 108.8 ;
    END
  END chany_top_out[0]
  PIN chany_top_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.65 107.44 14.79 108.8 ;
    END
  END chany_top_out[1]
  PIN chany_top_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.23 107.44 71.37 108.8 ;
    END
  END chany_top_out[2]
  PIN chany_top_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.73 107.44 13.87 108.8 ;
    END
  END chany_top_out[3]
  PIN chany_top_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.07 107.44 73.21 108.8 ;
    END
  END chany_top_out[4]
  PIN chany_top_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.15 107.44 49.29 108.8 ;
    END
  END chany_top_out[5]
  PIN chany_top_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.83 107.44 52.97 108.8 ;
    END
  END chany_top_out[6]
  PIN chany_top_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.01 107.44 22.15 108.8 ;
    END
  END chany_top_out[7]
  PIN chany_top_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.85 107.44 23.99 108.8 ;
    END
  END chany_top_out[8]
  PIN chany_top_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.93 107.44 23.07 108.8 ;
    END
  END chany_top_out[9]
  PIN chany_top_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.91 107.44 52.05 108.8 ;
    END
  END chany_top_out[10]
  PIN chany_top_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.75 107.44 30.89 108.8 ;
    END
  END chany_top_out[11]
  PIN chany_top_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.87 107.44 64.01 108.8 ;
    END
  END chany_top_out[12]
  PIN chany_top_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.15 107.44 72.29 108.8 ;
    END
  END chany_top_out[13]
  PIN chany_top_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.63 107.44 43.77 108.8 ;
    END
  END chany_top_out[14]
  PIN chany_top_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.39 107.44 46.53 108.8 ;
    END
  END chany_top_out[15]
  PIN chany_top_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.79 107.44 41.93 108.8 ;
    END
  END chany_top_out[16]
  PIN chany_top_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.83 107.44 29.97 108.8 ;
    END
  END chany_top_out[17]
  PIN chany_top_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.61 107.44 26.75 108.8 ;
    END
  END chany_top_out[18]
  PIN chany_top_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.77 107.44 24.91 108.8 ;
    END
  END chany_top_out[19]
  PIN right_grid_pin_52_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 83.26 78.73 84.64 79.03 ;
    END
  END right_grid_pin_52_[0]
  PIN left_grid_pin_0_[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 99.13 1.38 99.43 ;
    END
  END left_grid_pin_0_[0]
  PIN ccff_tail[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 78.73 1.38 79.03 ;
    END
  END ccff_tail[0]
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0 22.2 3.2 25.4 ;
        RECT 81.44 22.2 84.64 25.4 ;
        RECT 0 63 3.2 66.2 ;
        RECT 81.44 63 84.64 66.2 ;
        RECT 0 103.8 3.2 107 ;
        RECT 81.44 103.8 84.64 107 ;
      LAYER met4 ;
        RECT 12.58 0 13.18 0.6 ;
        RECT 42.02 0 42.62 0.6 ;
        RECT 71.46 0 72.06 0.6 ;
        RECT 12.58 108.2 13.18 108.8 ;
        RECT 42.02 108.2 42.62 108.8 ;
        RECT 71.46 108.2 72.06 108.8 ;
      LAYER met1 ;
        RECT 0 2.48 0.48 2.96 ;
        RECT 84.16 2.48 84.64 2.96 ;
        RECT 0 7.92 0.48 8.4 ;
        RECT 84.16 7.92 84.64 8.4 ;
        RECT 0 13.36 0.48 13.84 ;
        RECT 84.16 13.36 84.64 13.84 ;
        RECT 0 18.8 0.48 19.28 ;
        RECT 84.16 18.8 84.64 19.28 ;
        RECT 0 24.24 0.48 24.72 ;
        RECT 84.16 24.24 84.64 24.72 ;
        RECT 0 29.68 0.48 30.16 ;
        RECT 84.16 29.68 84.64 30.16 ;
        RECT 0 35.12 0.48 35.6 ;
        RECT 84.16 35.12 84.64 35.6 ;
        RECT 0 40.56 0.48 41.04 ;
        RECT 84.16 40.56 84.64 41.04 ;
        RECT 0 46 0.48 46.48 ;
        RECT 84.16 46 84.64 46.48 ;
        RECT 0 51.44 0.48 51.92 ;
        RECT 84.16 51.44 84.64 51.92 ;
        RECT 0 56.88 0.48 57.36 ;
        RECT 84.16 56.88 84.64 57.36 ;
        RECT 0 62.32 0.48 62.8 ;
        RECT 84.16 62.32 84.64 62.8 ;
        RECT 0 67.76 0.48 68.24 ;
        RECT 84.16 67.76 84.64 68.24 ;
        RECT 0 73.2 0.48 73.68 ;
        RECT 84.16 73.2 84.64 73.68 ;
        RECT 0 78.64 0.48 79.12 ;
        RECT 84.16 78.64 84.64 79.12 ;
        RECT 0 84.08 0.48 84.56 ;
        RECT 84.16 84.08 84.64 84.56 ;
        RECT 0 89.52 0.48 90 ;
        RECT 84.16 89.52 84.64 90 ;
        RECT 0 94.96 0.48 95.44 ;
        RECT 84.16 94.96 84.64 95.44 ;
        RECT 0 100.4 0.48 100.88 ;
        RECT 84.16 100.4 84.64 100.88 ;
        RECT 0 105.84 0.48 106.32 ;
        RECT 84.16 105.84 84.64 106.32 ;
    END
  END VDD
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0 1.8 3.2 5 ;
        RECT 81.44 1.8 84.64 5 ;
        RECT 0 42.6 3.2 45.8 ;
        RECT 81.44 42.6 84.64 45.8 ;
        RECT 0 83.4 3.2 86.6 ;
        RECT 81.44 83.4 84.64 86.6 ;
      LAYER met4 ;
        RECT 27.3 0 27.9 0.6 ;
        RECT 56.74 0 57.34 0.6 ;
        RECT 27.3 108.2 27.9 108.8 ;
        RECT 56.74 108.2 57.34 108.8 ;
      LAYER met1 ;
        RECT 0 0 84.64 0.24 ;
        RECT 0 5.2 0.48 5.68 ;
        RECT 84.16 5.2 84.64 5.68 ;
        RECT 0 10.64 0.48 11.12 ;
        RECT 84.16 10.64 84.64 11.12 ;
        RECT 0 16.08 0.48 16.56 ;
        RECT 84.16 16.08 84.64 16.56 ;
        RECT 0 21.52 0.48 22 ;
        RECT 84.16 21.52 84.64 22 ;
        RECT 0 26.96 0.48 27.44 ;
        RECT 84.16 26.96 84.64 27.44 ;
        RECT 0 32.4 0.48 32.88 ;
        RECT 84.16 32.4 84.64 32.88 ;
        RECT 0 37.84 0.48 38.32 ;
        RECT 84.16 37.84 84.64 38.32 ;
        RECT 0 43.28 0.48 43.76 ;
        RECT 84.16 43.28 84.64 43.76 ;
        RECT 0 48.72 0.48 49.2 ;
        RECT 84.16 48.72 84.64 49.2 ;
        RECT 0 54.16 0.48 54.64 ;
        RECT 84.16 54.16 84.64 54.64 ;
        RECT 0 59.6 0.48 60.08 ;
        RECT 84.16 59.6 84.64 60.08 ;
        RECT 0 65.04 0.48 65.52 ;
        RECT 84.16 65.04 84.64 65.52 ;
        RECT 0 70.48 0.48 70.96 ;
        RECT 84.16 70.48 84.64 70.96 ;
        RECT 0 75.92 0.48 76.4 ;
        RECT 84.16 75.92 84.64 76.4 ;
        RECT 0 81.36 0.48 81.84 ;
        RECT 84.16 81.36 84.64 81.84 ;
        RECT 0 86.8 0.48 87.28 ;
        RECT 84.16 86.8 84.64 87.28 ;
        RECT 0 92.24 0.48 92.72 ;
        RECT 84.16 92.24 84.64 92.72 ;
        RECT 0 97.68 0.48 98.16 ;
        RECT 84.16 97.68 84.64 98.16 ;
        RECT 0 103.12 0.48 103.6 ;
        RECT 84.16 103.12 84.64 103.6 ;
        RECT 0 108.56 84.64 108.8 ;
    END
  END VSS
  OBS
    LAYER li1 ;
      RECT 0 108.715 84.64 108.885 ;
      RECT 80.96 105.995 84.64 106.165 ;
      RECT 0 105.995 3.68 106.165 ;
      RECT 83.72 103.275 84.64 103.445 ;
      RECT 0 103.275 3.68 103.445 ;
      RECT 83.72 100.555 84.64 100.725 ;
      RECT 0 100.555 3.68 100.725 ;
      RECT 84.18 97.835 84.64 98.005 ;
      RECT 0 97.835 3.68 98.005 ;
      RECT 84.18 95.115 84.64 95.285 ;
      RECT 0 95.115 3.68 95.285 ;
      RECT 84.18 92.395 84.64 92.565 ;
      RECT 0 92.395 3.68 92.565 ;
      RECT 84.18 89.675 84.64 89.845 ;
      RECT 0 89.675 3.68 89.845 ;
      RECT 84.18 86.955 84.64 87.125 ;
      RECT 0 86.955 3.68 87.125 ;
      RECT 83.72 84.235 84.64 84.405 ;
      RECT 0 84.235 1.84 84.405 ;
      RECT 83.72 81.515 84.64 81.685 ;
      RECT 0 81.515 1.84 81.685 ;
      RECT 83.72 78.795 84.64 78.965 ;
      RECT 0 78.795 3.68 78.965 ;
      RECT 80.96 76.075 84.64 76.245 ;
      RECT 0 76.075 3.68 76.245 ;
      RECT 80.96 73.355 84.64 73.525 ;
      RECT 0 73.355 3.68 73.525 ;
      RECT 82.8 70.635 84.64 70.805 ;
      RECT 0 70.635 3.68 70.805 ;
      RECT 82.8 67.915 84.64 68.085 ;
      RECT 0 67.915 3.68 68.085 ;
      RECT 83.72 65.195 84.64 65.365 ;
      RECT 0 65.195 3.68 65.365 ;
      RECT 83.72 62.475 84.64 62.645 ;
      RECT 0 62.475 3.68 62.645 ;
      RECT 83.72 59.755 84.64 59.925 ;
      RECT 0 59.755 3.68 59.925 ;
      RECT 80.96 57.035 84.64 57.205 ;
      RECT 0 57.035 3.68 57.205 ;
      RECT 80.96 54.315 84.64 54.485 ;
      RECT 0 54.315 3.68 54.485 ;
      RECT 80.96 51.595 84.64 51.765 ;
      RECT 0 51.595 3.68 51.765 ;
      RECT 80.96 48.875 84.64 49.045 ;
      RECT 0 48.875 3.68 49.045 ;
      RECT 80.96 46.155 84.64 46.325 ;
      RECT 0 46.155 3.68 46.325 ;
      RECT 80.96 43.435 84.64 43.605 ;
      RECT 0 43.435 3.68 43.605 ;
      RECT 80.96 40.715 84.64 40.885 ;
      RECT 0 40.715 3.68 40.885 ;
      RECT 80.96 37.995 84.64 38.165 ;
      RECT 0 37.995 3.68 38.165 ;
      RECT 80.96 35.275 84.64 35.445 ;
      RECT 0 35.275 3.68 35.445 ;
      RECT 80.96 32.555 84.64 32.725 ;
      RECT 0 32.555 3.68 32.725 ;
      RECT 80.96 29.835 84.64 30.005 ;
      RECT 0 29.835 3.68 30.005 ;
      RECT 80.96 27.115 84.64 27.285 ;
      RECT 0 27.115 3.68 27.285 ;
      RECT 82.8 24.395 84.64 24.565 ;
      RECT 0 24.395 3.68 24.565 ;
      RECT 82.8 21.675 84.64 21.845 ;
      RECT 0 21.675 3.68 21.845 ;
      RECT 82.8 18.955 84.64 19.125 ;
      RECT 0 18.955 3.68 19.125 ;
      RECT 82.8 16.235 84.64 16.405 ;
      RECT 0 16.235 3.68 16.405 ;
      RECT 84.18 13.515 84.64 13.685 ;
      RECT 0 13.515 3.68 13.685 ;
      RECT 84.18 10.795 84.64 10.965 ;
      RECT 0 10.795 3.68 10.965 ;
      RECT 83.72 8.075 84.64 8.245 ;
      RECT 0 8.075 3.68 8.245 ;
      RECT 80.96 5.355 84.64 5.525 ;
      RECT 0 5.355 3.68 5.525 ;
      RECT 80.96 2.635 84.64 2.805 ;
      RECT 0 2.635 3.68 2.805 ;
      RECT 0 -0.085 84.64 0.085 ;
    LAYER met3 ;
      POLYGON 57.205 108.965 57.205 108.96 57.42 108.96 57.42 108.64 57.205 108.64 57.205 108.635 56.875 108.635 56.875 108.64 56.66 108.64 56.66 108.96 56.875 108.96 56.875 108.965 ;
      POLYGON 27.765 108.965 27.765 108.96 27.98 108.96 27.98 108.64 27.765 108.64 27.765 108.635 27.435 108.635 27.435 108.64 27.22 108.64 27.22 108.96 27.435 108.96 27.435 108.965 ;
      POLYGON 57.205 0.165 57.205 0.16 57.42 0.16 57.42 -0.16 57.205 -0.16 57.205 -0.165 56.875 -0.165 56.875 -0.16 56.66 -0.16 56.66 0.16 56.875 0.16 56.875 0.165 ;
      POLYGON 27.765 0.165 27.765 0.16 27.98 0.16 27.98 -0.16 27.765 -0.16 27.765 -0.165 27.435 -0.165 27.435 -0.16 27.22 -0.16 27.22 0.16 27.435 0.16 27.435 0.165 ;
      POLYGON 84.24 108.4 84.24 79.43 82.86 79.43 82.86 78.33 84.24 78.33 84.24 0.4 0.4 0.4 0.4 2.85 1.78 2.85 1.78 3.95 0.4 3.95 0.4 78.33 1.78 78.33 1.78 79.43 0.4 79.43 0.4 98.73 1.78 98.73 1.78 99.83 0.4 99.83 0.4 108.4 ;
    LAYER met2 ;
      RECT 56.9 108.615 57.18 108.985 ;
      RECT 27.46 108.615 27.74 108.985 ;
      RECT 51.39 106.94 51.65 107.26 ;
      RECT 41.27 106.94 41.53 107.26 ;
      RECT 56.9 -0.185 57.18 0.185 ;
      RECT 27.46 -0.185 27.74 0.185 ;
      POLYGON 84.36 108.52 84.36 0.28 72.57 0.28 72.57 1.64 71.87 1.64 71.87 0.28 71.65 0.28 71.65 1.64 70.95 1.64 70.95 0.28 70.73 0.28 70.73 1.64 70.03 1.64 70.03 0.28 69.81 0.28 69.81 1.64 69.11 1.64 69.11 0.28 68.89 0.28 68.89 1.64 68.19 1.64 68.19 0.28 67.97 0.28 67.97 1.64 67.27 1.64 67.27 0.28 63.37 0.28 63.37 1.64 62.67 1.64 62.67 0.28 62.45 0.28 62.45 1.64 61.75 1.64 61.75 0.28 53.25 0.28 53.25 1.64 52.55 1.64 52.55 0.28 52.33 0.28 52.33 1.64 51.63 1.64 51.63 0.28 51.41 0.28 51.41 1.64 50.71 1.64 50.71 0.28 50.49 0.28 50.49 1.64 49.79 1.64 49.79 0.28 49.57 0.28 49.57 1.64 48.87 1.64 48.87 0.28 48.65 0.28 48.65 1.64 47.95 1.64 47.95 0.28 47.73 0.28 47.73 1.64 47.03 1.64 47.03 0.28 46.81 0.28 46.81 1.64 46.11 1.64 46.11 0.28 45.89 0.28 45.89 1.64 45.19 1.64 45.19 0.28 44.97 0.28 44.97 1.64 44.27 1.64 44.27 0.28 44.05 0.28 44.05 1.64 43.35 1.64 43.35 0.28 43.13 0.28 43.13 1.64 42.43 1.64 42.43 0.28 42.21 0.28 42.21 1.64 41.51 1.64 41.51 0.28 36.69 0.28 36.69 1.64 35.99 1.64 35.99 0.28 29.33 0.28 29.33 1.64 28.63 1.64 28.63 0.28 26.11 0.28 26.11 1.64 25.41 1.64 25.41 0.28 7.71 0.28 7.71 1.64 7.01 1.64 7.01 0.28 0.28 0.28 0.28 108.52 13.45 108.52 13.45 107.16 14.15 107.16 14.15 108.52 14.37 108.52 14.37 107.16 15.07 107.16 15.07 108.52 21.73 108.52 21.73 107.16 22.43 107.16 22.43 108.52 22.65 108.52 22.65 107.16 23.35 107.16 23.35 108.52 23.57 108.52 23.57 107.16 24.27 107.16 24.27 108.52 24.49 108.52 24.49 107.16 25.19 107.16 25.19 108.52 25.41 108.52 25.41 107.16 26.11 107.16 26.11 108.52 26.33 108.52 26.33 107.16 27.03 107.16 27.03 108.52 28.17 108.52 28.17 107.16 28.87 107.16 28.87 108.52 29.55 108.52 29.55 107.16 30.25 107.16 30.25 108.52 30.47 108.52 30.47 107.16 31.17 107.16 31.17 108.52 34.15 108.52 34.15 107.16 34.85 107.16 34.85 108.52 41.51 108.52 41.51 107.16 42.21 107.16 42.21 108.52 42.43 108.52 42.43 107.16 43.13 107.16 43.13 108.52 43.35 108.52 43.35 107.16 44.05 107.16 44.05 108.52 44.27 108.52 44.27 107.16 44.97 107.16 44.97 108.52 45.19 108.52 45.19 107.16 45.89 107.16 45.89 108.52 46.11 108.52 46.11 107.16 46.81 107.16 46.81 108.52 47.03 108.52 47.03 107.16 47.73 107.16 47.73 108.52 47.95 108.52 47.95 107.16 48.65 107.16 48.65 108.52 48.87 108.52 48.87 107.16 49.57 107.16 49.57 108.52 49.79 108.52 49.79 107.16 50.49 107.16 50.49 108.52 50.71 108.52 50.71 107.16 51.41 107.16 51.41 108.52 51.63 108.52 51.63 107.16 52.33 107.16 52.33 108.52 52.55 108.52 52.55 107.16 53.25 107.16 53.25 108.52 53.93 108.52 53.93 107.16 54.63 107.16 54.63 108.52 63.59 108.52 63.59 107.16 64.29 107.16 64.29 108.52 65.43 108.52 65.43 107.16 66.13 107.16 66.13 108.52 66.35 108.52 66.35 107.16 67.05 107.16 67.05 108.52 67.27 108.52 67.27 107.16 67.97 107.16 67.97 108.52 68.19 108.52 68.19 107.16 68.89 107.16 68.89 108.52 69.11 108.52 69.11 107.16 69.81 107.16 69.81 108.52 70.03 108.52 70.03 107.16 70.73 107.16 70.73 108.52 70.95 108.52 70.95 107.16 71.65 107.16 71.65 108.52 71.87 108.52 71.87 107.16 72.57 107.16 72.57 108.52 72.79 108.52 72.79 107.16 73.49 107.16 73.49 108.52 ;
    LAYER met4 ;
      POLYGON 84.24 108.4 84.24 0.4 72.46 0.4 72.46 1 71.06 1 71.06 0.4 69.55 0.4 69.55 1.76 68.45 1.76 68.45 0.4 59.43 0.4 59.43 1.76 58.33 1.76 58.33 0.4 57.74 0.4 57.74 1 56.34 1 56.34 0.4 50.23 0.4 50.23 1.76 49.13 1.76 49.13 0.4 48.39 0.4 48.39 1.76 47.29 1.76 47.29 0.4 46.55 0.4 46.55 1.76 45.45 1.76 45.45 0.4 44.71 0.4 44.71 1.76 43.61 1.76 43.61 0.4 43.02 0.4 43.02 1 41.62 1 41.62 0.4 29.99 0.4 29.99 1.76 28.89 1.76 28.89 0.4 28.3 0.4 28.3 1 26.9 1 26.9 0.4 26.31 0.4 26.31 1.76 25.21 1.76 25.21 0.4 24.47 0.4 24.47 1.76 23.37 1.76 23.37 0.4 22.63 0.4 22.63 1.76 21.53 1.76 21.53 0.4 20.79 0.4 20.79 1.76 19.69 1.76 19.69 0.4 15.27 0.4 15.27 1.76 14.17 1.76 14.17 0.4 13.58 0.4 13.58 1 12.18 1 12.18 0.4 9.75 0.4 9.75 1.76 8.65 1.76 8.65 0.4 7.91 0.4 7.91 1.76 6.81 1.76 6.81 0.4 6.07 0.4 6.07 1.76 4.97 1.76 4.97 0.4 0.4 0.4 0.4 108.4 12.18 108.4 12.18 107.8 13.58 107.8 13.58 108.4 23.37 108.4 23.37 107.04 24.47 107.04 24.47 108.4 25.21 108.4 25.21 107.04 26.31 107.04 26.31 108.4 26.9 108.4 26.9 107.8 28.3 107.8 28.3 108.4 41.62 108.4 41.62 107.8 43.02 107.8 43.02 108.4 45.45 108.4 45.45 107.04 46.55 107.04 46.55 108.4 47.29 108.4 47.29 107.04 48.39 107.04 48.39 108.4 49.13 108.4 49.13 107.04 50.23 107.04 50.23 108.4 56.34 108.4 56.34 107.8 57.74 107.8 57.74 108.4 71.06 108.4 71.06 107.8 72.46 107.8 72.46 108.4 ;
    LAYER met1 ;
      POLYGON 84.36 108.28 84.36 106.6 83.88 106.6 83.88 105.56 84.36 105.56 84.36 103.88 83.88 103.88 83.88 102.84 84.36 102.84 84.36 101.16 83.88 101.16 83.88 100.12 84.36 100.12 84.36 98.44 83.88 98.44 83.88 97.4 84.36 97.4 84.36 95.72 83.88 95.72 83.88 94.68 84.36 94.68 84.36 93 83.88 93 83.88 91.96 84.36 91.96 84.36 90.28 83.88 90.28 83.88 89.24 84.36 89.24 84.36 87.56 83.88 87.56 83.88 86.52 84.36 86.52 84.36 84.84 83.88 84.84 83.88 83.8 84.36 83.8 84.36 82.12 83.88 82.12 83.88 81.08 84.36 81.08 84.36 79.4 83.88 79.4 83.88 78.36 84.36 78.36 84.36 76.68 83.88 76.68 83.88 75.64 84.36 75.64 84.36 73.96 83.88 73.96 83.88 72.92 84.36 72.92 84.36 71.24 83.88 71.24 83.88 70.2 84.36 70.2 84.36 68.52 83.88 68.52 83.88 67.48 84.36 67.48 84.36 65.8 83.88 65.8 83.88 64.76 84.36 64.76 84.36 63.08 83.88 63.08 83.88 62.04 84.36 62.04 84.36 60.36 83.88 60.36 83.88 59.32 84.36 59.32 84.36 57.64 83.88 57.64 83.88 56.6 84.36 56.6 84.36 54.92 83.88 54.92 83.88 53.88 84.36 53.88 84.36 52.2 83.88 52.2 83.88 51.16 84.36 51.16 84.36 49.48 83.88 49.48 83.88 48.44 84.36 48.44 84.36 46.76 83.88 46.76 83.88 45.72 84.36 45.72 84.36 44.04 83.88 44.04 83.88 43 84.36 43 84.36 41.32 83.88 41.32 83.88 40.28 84.36 40.28 84.36 38.6 83.88 38.6 83.88 37.56 84.36 37.56 84.36 35.88 83.88 35.88 83.88 34.84 84.36 34.84 84.36 33.16 83.88 33.16 83.88 32.12 84.36 32.12 84.36 30.44 83.88 30.44 83.88 29.4 84.36 29.4 84.36 27.72 83.88 27.72 83.88 26.68 84.36 26.68 84.36 25 83.88 25 83.88 23.96 84.36 23.96 84.36 22.28 83.88 22.28 83.88 21.24 84.36 21.24 84.36 19.56 83.88 19.56 83.88 18.52 84.36 18.52 84.36 16.84 83.88 16.84 83.88 15.8 84.36 15.8 84.36 14.12 83.88 14.12 83.88 13.08 84.36 13.08 84.36 11.4 83.88 11.4 83.88 10.36 84.36 10.36 84.36 8.68 83.88 8.68 83.88 7.64 84.36 7.64 84.36 5.96 83.88 5.96 83.88 4.92 84.36 4.92 84.36 3.24 83.88 3.24 83.88 2.2 84.36 2.2 84.36 0.52 0.28 0.52 0.28 2.2 0.76 2.2 0.76 3.24 0.28 3.24 0.28 4.92 0.76 4.92 0.76 5.96 0.28 5.96 0.28 7.64 0.76 7.64 0.76 8.68 0.28 8.68 0.28 10.36 0.76 10.36 0.76 11.4 0.28 11.4 0.28 13.08 0.76 13.08 0.76 14.12 0.28 14.12 0.28 15.8 0.76 15.8 0.76 16.84 0.28 16.84 0.28 18.52 0.76 18.52 0.76 19.56 0.28 19.56 0.28 21.24 0.76 21.24 0.76 22.28 0.28 22.28 0.28 23.96 0.76 23.96 0.76 25 0.28 25 0.28 26.68 0.76 26.68 0.76 27.72 0.28 27.72 0.28 29.4 0.76 29.4 0.76 30.44 0.28 30.44 0.28 32.12 0.76 32.12 0.76 33.16 0.28 33.16 0.28 34.84 0.76 34.84 0.76 35.88 0.28 35.88 0.28 37.56 0.76 37.56 0.76 38.6 0.28 38.6 0.28 40.28 0.76 40.28 0.76 41.32 0.28 41.32 0.28 43 0.76 43 0.76 44.04 0.28 44.04 0.28 45.72 0.76 45.72 0.76 46.76 0.28 46.76 0.28 48.44 0.76 48.44 0.76 49.48 0.28 49.48 0.28 51.16 0.76 51.16 0.76 52.2 0.28 52.2 0.28 53.88 0.76 53.88 0.76 54.92 0.28 54.92 0.28 56.6 0.76 56.6 0.76 57.64 0.28 57.64 0.28 59.32 0.76 59.32 0.76 60.36 0.28 60.36 0.28 62.04 0.76 62.04 0.76 63.08 0.28 63.08 0.28 64.76 0.76 64.76 0.76 65.8 0.28 65.8 0.28 67.48 0.76 67.48 0.76 68.52 0.28 68.52 0.28 70.2 0.76 70.2 0.76 71.24 0.28 71.24 0.28 72.92 0.76 72.92 0.76 73.96 0.28 73.96 0.28 75.64 0.76 75.64 0.76 76.68 0.28 76.68 0.28 78.36 0.76 78.36 0.76 79.4 0.28 79.4 0.28 81.08 0.76 81.08 0.76 82.12 0.28 82.12 0.28 83.8 0.76 83.8 0.76 84.84 0.28 84.84 0.28 86.52 0.76 86.52 0.76 87.56 0.28 87.56 0.28 89.24 0.76 89.24 0.76 90.28 0.28 90.28 0.28 91.96 0.76 91.96 0.76 93 0.28 93 0.28 94.68 0.76 94.68 0.76 95.72 0.28 95.72 0.28 97.4 0.76 97.4 0.76 98.44 0.28 98.44 0.28 100.12 0.76 100.12 0.76 101.16 0.28 101.16 0.28 102.84 0.76 102.84 0.76 103.88 0.28 103.88 0.28 105.56 0.76 105.56 0.76 106.6 0.28 106.6 0.28 108.28 ;
    LAYER met5 ;
      RECT 6.4 103.8 78.24 107 ;
      RECT 6.4 1.8 78.24 5 ;
      POLYGON 78.24 105.6 78.24 100.6 81.44 100.6 81.44 89.8 78.24 89.8 78.24 80.2 81.44 80.2 81.44 69.4 78.24 69.4 78.24 59.8 81.44 59.8 81.44 49 78.24 49 78.24 39.4 81.44 39.4 81.44 28.6 78.24 28.6 78.24 19 81.44 19 81.44 8.2 78.24 8.2 78.24 3.2 6.4 3.2 6.4 8.2 3.2 8.2 3.2 19 6.4 19 6.4 28.6 3.2 28.6 3.2 39.4 6.4 39.4 6.4 49 3.2 49 3.2 59.8 6.4 59.8 6.4 69.4 3.2 69.4 3.2 80.2 6.4 80.2 6.4 89.8 3.2 89.8 3.2 100.6 6.4 100.6 6.4 105.6 ;
    LAYER li1 ;
      RECT 0.34 0.34 84.3 108.46 ;
    LAYER mcon ;
      RECT 84.325 108.715 84.495 108.885 ;
      RECT 83.865 108.715 84.035 108.885 ;
      RECT 83.405 108.715 83.575 108.885 ;
      RECT 82.945 108.715 83.115 108.885 ;
      RECT 82.485 108.715 82.655 108.885 ;
      RECT 82.025 108.715 82.195 108.885 ;
      RECT 81.565 108.715 81.735 108.885 ;
      RECT 81.105 108.715 81.275 108.885 ;
      RECT 80.645 108.715 80.815 108.885 ;
      RECT 80.185 108.715 80.355 108.885 ;
      RECT 79.725 108.715 79.895 108.885 ;
      RECT 79.265 108.715 79.435 108.885 ;
      RECT 78.805 108.715 78.975 108.885 ;
      RECT 78.345 108.715 78.515 108.885 ;
      RECT 77.885 108.715 78.055 108.885 ;
      RECT 77.425 108.715 77.595 108.885 ;
      RECT 76.965 108.715 77.135 108.885 ;
      RECT 76.505 108.715 76.675 108.885 ;
      RECT 76.045 108.715 76.215 108.885 ;
      RECT 75.585 108.715 75.755 108.885 ;
      RECT 75.125 108.715 75.295 108.885 ;
      RECT 74.665 108.715 74.835 108.885 ;
      RECT 74.205 108.715 74.375 108.885 ;
      RECT 73.745 108.715 73.915 108.885 ;
      RECT 73.285 108.715 73.455 108.885 ;
      RECT 72.825 108.715 72.995 108.885 ;
      RECT 72.365 108.715 72.535 108.885 ;
      RECT 71.905 108.715 72.075 108.885 ;
      RECT 71.445 108.715 71.615 108.885 ;
      RECT 70.985 108.715 71.155 108.885 ;
      RECT 70.525 108.715 70.695 108.885 ;
      RECT 70.065 108.715 70.235 108.885 ;
      RECT 69.605 108.715 69.775 108.885 ;
      RECT 69.145 108.715 69.315 108.885 ;
      RECT 68.685 108.715 68.855 108.885 ;
      RECT 68.225 108.715 68.395 108.885 ;
      RECT 67.765 108.715 67.935 108.885 ;
      RECT 67.305 108.715 67.475 108.885 ;
      RECT 66.845 108.715 67.015 108.885 ;
      RECT 66.385 108.715 66.555 108.885 ;
      RECT 65.925 108.715 66.095 108.885 ;
      RECT 65.465 108.715 65.635 108.885 ;
      RECT 65.005 108.715 65.175 108.885 ;
      RECT 64.545 108.715 64.715 108.885 ;
      RECT 64.085 108.715 64.255 108.885 ;
      RECT 63.625 108.715 63.795 108.885 ;
      RECT 63.165 108.715 63.335 108.885 ;
      RECT 62.705 108.715 62.875 108.885 ;
      RECT 62.245 108.715 62.415 108.885 ;
      RECT 61.785 108.715 61.955 108.885 ;
      RECT 61.325 108.715 61.495 108.885 ;
      RECT 60.865 108.715 61.035 108.885 ;
      RECT 60.405 108.715 60.575 108.885 ;
      RECT 59.945 108.715 60.115 108.885 ;
      RECT 59.485 108.715 59.655 108.885 ;
      RECT 59.025 108.715 59.195 108.885 ;
      RECT 58.565 108.715 58.735 108.885 ;
      RECT 58.105 108.715 58.275 108.885 ;
      RECT 57.645 108.715 57.815 108.885 ;
      RECT 57.185 108.715 57.355 108.885 ;
      RECT 56.725 108.715 56.895 108.885 ;
      RECT 56.265 108.715 56.435 108.885 ;
      RECT 55.805 108.715 55.975 108.885 ;
      RECT 55.345 108.715 55.515 108.885 ;
      RECT 54.885 108.715 55.055 108.885 ;
      RECT 54.425 108.715 54.595 108.885 ;
      RECT 53.965 108.715 54.135 108.885 ;
      RECT 53.505 108.715 53.675 108.885 ;
      RECT 53.045 108.715 53.215 108.885 ;
      RECT 52.585 108.715 52.755 108.885 ;
      RECT 52.125 108.715 52.295 108.885 ;
      RECT 51.665 108.715 51.835 108.885 ;
      RECT 51.205 108.715 51.375 108.885 ;
      RECT 50.745 108.715 50.915 108.885 ;
      RECT 50.285 108.715 50.455 108.885 ;
      RECT 49.825 108.715 49.995 108.885 ;
      RECT 49.365 108.715 49.535 108.885 ;
      RECT 48.905 108.715 49.075 108.885 ;
      RECT 48.445 108.715 48.615 108.885 ;
      RECT 47.985 108.715 48.155 108.885 ;
      RECT 47.525 108.715 47.695 108.885 ;
      RECT 47.065 108.715 47.235 108.885 ;
      RECT 46.605 108.715 46.775 108.885 ;
      RECT 46.145 108.715 46.315 108.885 ;
      RECT 45.685 108.715 45.855 108.885 ;
      RECT 45.225 108.715 45.395 108.885 ;
      RECT 44.765 108.715 44.935 108.885 ;
      RECT 44.305 108.715 44.475 108.885 ;
      RECT 43.845 108.715 44.015 108.885 ;
      RECT 43.385 108.715 43.555 108.885 ;
      RECT 42.925 108.715 43.095 108.885 ;
      RECT 42.465 108.715 42.635 108.885 ;
      RECT 42.005 108.715 42.175 108.885 ;
      RECT 41.545 108.715 41.715 108.885 ;
      RECT 41.085 108.715 41.255 108.885 ;
      RECT 40.625 108.715 40.795 108.885 ;
      RECT 40.165 108.715 40.335 108.885 ;
      RECT 39.705 108.715 39.875 108.885 ;
      RECT 39.245 108.715 39.415 108.885 ;
      RECT 38.785 108.715 38.955 108.885 ;
      RECT 38.325 108.715 38.495 108.885 ;
      RECT 37.865 108.715 38.035 108.885 ;
      RECT 37.405 108.715 37.575 108.885 ;
      RECT 36.945 108.715 37.115 108.885 ;
      RECT 36.485 108.715 36.655 108.885 ;
      RECT 36.025 108.715 36.195 108.885 ;
      RECT 35.565 108.715 35.735 108.885 ;
      RECT 35.105 108.715 35.275 108.885 ;
      RECT 34.645 108.715 34.815 108.885 ;
      RECT 34.185 108.715 34.355 108.885 ;
      RECT 33.725 108.715 33.895 108.885 ;
      RECT 33.265 108.715 33.435 108.885 ;
      RECT 32.805 108.715 32.975 108.885 ;
      RECT 32.345 108.715 32.515 108.885 ;
      RECT 31.885 108.715 32.055 108.885 ;
      RECT 31.425 108.715 31.595 108.885 ;
      RECT 30.965 108.715 31.135 108.885 ;
      RECT 30.505 108.715 30.675 108.885 ;
      RECT 30.045 108.715 30.215 108.885 ;
      RECT 29.585 108.715 29.755 108.885 ;
      RECT 29.125 108.715 29.295 108.885 ;
      RECT 28.665 108.715 28.835 108.885 ;
      RECT 28.205 108.715 28.375 108.885 ;
      RECT 27.745 108.715 27.915 108.885 ;
      RECT 27.285 108.715 27.455 108.885 ;
      RECT 26.825 108.715 26.995 108.885 ;
      RECT 26.365 108.715 26.535 108.885 ;
      RECT 25.905 108.715 26.075 108.885 ;
      RECT 25.445 108.715 25.615 108.885 ;
      RECT 24.985 108.715 25.155 108.885 ;
      RECT 24.525 108.715 24.695 108.885 ;
      RECT 24.065 108.715 24.235 108.885 ;
      RECT 23.605 108.715 23.775 108.885 ;
      RECT 23.145 108.715 23.315 108.885 ;
      RECT 22.685 108.715 22.855 108.885 ;
      RECT 22.225 108.715 22.395 108.885 ;
      RECT 21.765 108.715 21.935 108.885 ;
      RECT 21.305 108.715 21.475 108.885 ;
      RECT 20.845 108.715 21.015 108.885 ;
      RECT 20.385 108.715 20.555 108.885 ;
      RECT 19.925 108.715 20.095 108.885 ;
      RECT 19.465 108.715 19.635 108.885 ;
      RECT 19.005 108.715 19.175 108.885 ;
      RECT 18.545 108.715 18.715 108.885 ;
      RECT 18.085 108.715 18.255 108.885 ;
      RECT 17.625 108.715 17.795 108.885 ;
      RECT 17.165 108.715 17.335 108.885 ;
      RECT 16.705 108.715 16.875 108.885 ;
      RECT 16.245 108.715 16.415 108.885 ;
      RECT 15.785 108.715 15.955 108.885 ;
      RECT 15.325 108.715 15.495 108.885 ;
      RECT 14.865 108.715 15.035 108.885 ;
      RECT 14.405 108.715 14.575 108.885 ;
      RECT 13.945 108.715 14.115 108.885 ;
      RECT 13.485 108.715 13.655 108.885 ;
      RECT 13.025 108.715 13.195 108.885 ;
      RECT 12.565 108.715 12.735 108.885 ;
      RECT 12.105 108.715 12.275 108.885 ;
      RECT 11.645 108.715 11.815 108.885 ;
      RECT 11.185 108.715 11.355 108.885 ;
      RECT 10.725 108.715 10.895 108.885 ;
      RECT 10.265 108.715 10.435 108.885 ;
      RECT 9.805 108.715 9.975 108.885 ;
      RECT 9.345 108.715 9.515 108.885 ;
      RECT 8.885 108.715 9.055 108.885 ;
      RECT 8.425 108.715 8.595 108.885 ;
      RECT 7.965 108.715 8.135 108.885 ;
      RECT 7.505 108.715 7.675 108.885 ;
      RECT 7.045 108.715 7.215 108.885 ;
      RECT 6.585 108.715 6.755 108.885 ;
      RECT 6.125 108.715 6.295 108.885 ;
      RECT 5.665 108.715 5.835 108.885 ;
      RECT 5.205 108.715 5.375 108.885 ;
      RECT 4.745 108.715 4.915 108.885 ;
      RECT 4.285 108.715 4.455 108.885 ;
      RECT 3.825 108.715 3.995 108.885 ;
      RECT 3.365 108.715 3.535 108.885 ;
      RECT 2.905 108.715 3.075 108.885 ;
      RECT 2.445 108.715 2.615 108.885 ;
      RECT 1.985 108.715 2.155 108.885 ;
      RECT 1.525 108.715 1.695 108.885 ;
      RECT 1.065 108.715 1.235 108.885 ;
      RECT 0.605 108.715 0.775 108.885 ;
      RECT 0.145 108.715 0.315 108.885 ;
      RECT 84.325 105.995 84.495 106.165 ;
      RECT 83.865 105.995 84.035 106.165 ;
      RECT 0.605 105.995 0.775 106.165 ;
      RECT 0.145 105.995 0.315 106.165 ;
      RECT 84.325 103.275 84.495 103.445 ;
      RECT 83.865 103.275 84.035 103.445 ;
      RECT 0.605 103.275 0.775 103.445 ;
      RECT 0.145 103.275 0.315 103.445 ;
      RECT 84.325 100.555 84.495 100.725 ;
      RECT 83.865 100.555 84.035 100.725 ;
      RECT 0.605 100.555 0.775 100.725 ;
      RECT 0.145 100.555 0.315 100.725 ;
      RECT 84.325 97.835 84.495 98.005 ;
      RECT 83.865 97.835 84.035 98.005 ;
      RECT 0.605 97.835 0.775 98.005 ;
      RECT 0.145 97.835 0.315 98.005 ;
      RECT 84.325 95.115 84.495 95.285 ;
      RECT 83.865 95.115 84.035 95.285 ;
      RECT 0.605 95.115 0.775 95.285 ;
      RECT 0.145 95.115 0.315 95.285 ;
      RECT 84.325 92.395 84.495 92.565 ;
      RECT 83.865 92.395 84.035 92.565 ;
      RECT 0.605 92.395 0.775 92.565 ;
      RECT 0.145 92.395 0.315 92.565 ;
      RECT 84.325 89.675 84.495 89.845 ;
      RECT 83.865 89.675 84.035 89.845 ;
      RECT 0.605 89.675 0.775 89.845 ;
      RECT 0.145 89.675 0.315 89.845 ;
      RECT 84.325 86.955 84.495 87.125 ;
      RECT 83.865 86.955 84.035 87.125 ;
      RECT 0.605 86.955 0.775 87.125 ;
      RECT 0.145 86.955 0.315 87.125 ;
      RECT 84.325 84.235 84.495 84.405 ;
      RECT 83.865 84.235 84.035 84.405 ;
      RECT 0.605 84.235 0.775 84.405 ;
      RECT 0.145 84.235 0.315 84.405 ;
      RECT 84.325 81.515 84.495 81.685 ;
      RECT 83.865 81.515 84.035 81.685 ;
      RECT 0.605 81.515 0.775 81.685 ;
      RECT 0.145 81.515 0.315 81.685 ;
      RECT 84.325 78.795 84.495 78.965 ;
      RECT 83.865 78.795 84.035 78.965 ;
      RECT 0.605 78.795 0.775 78.965 ;
      RECT 0.145 78.795 0.315 78.965 ;
      RECT 84.325 76.075 84.495 76.245 ;
      RECT 83.865 76.075 84.035 76.245 ;
      RECT 0.605 76.075 0.775 76.245 ;
      RECT 0.145 76.075 0.315 76.245 ;
      RECT 84.325 73.355 84.495 73.525 ;
      RECT 83.865 73.355 84.035 73.525 ;
      RECT 0.605 73.355 0.775 73.525 ;
      RECT 0.145 73.355 0.315 73.525 ;
      RECT 84.325 70.635 84.495 70.805 ;
      RECT 83.865 70.635 84.035 70.805 ;
      RECT 0.605 70.635 0.775 70.805 ;
      RECT 0.145 70.635 0.315 70.805 ;
      RECT 84.325 67.915 84.495 68.085 ;
      RECT 83.865 67.915 84.035 68.085 ;
      RECT 0.605 67.915 0.775 68.085 ;
      RECT 0.145 67.915 0.315 68.085 ;
      RECT 84.325 65.195 84.495 65.365 ;
      RECT 83.865 65.195 84.035 65.365 ;
      RECT 0.605 65.195 0.775 65.365 ;
      RECT 0.145 65.195 0.315 65.365 ;
      RECT 84.325 62.475 84.495 62.645 ;
      RECT 83.865 62.475 84.035 62.645 ;
      RECT 0.605 62.475 0.775 62.645 ;
      RECT 0.145 62.475 0.315 62.645 ;
      RECT 84.325 59.755 84.495 59.925 ;
      RECT 83.865 59.755 84.035 59.925 ;
      RECT 0.605 59.755 0.775 59.925 ;
      RECT 0.145 59.755 0.315 59.925 ;
      RECT 84.325 57.035 84.495 57.205 ;
      RECT 83.865 57.035 84.035 57.205 ;
      RECT 0.605 57.035 0.775 57.205 ;
      RECT 0.145 57.035 0.315 57.205 ;
      RECT 84.325 54.315 84.495 54.485 ;
      RECT 83.865 54.315 84.035 54.485 ;
      RECT 0.605 54.315 0.775 54.485 ;
      RECT 0.145 54.315 0.315 54.485 ;
      RECT 84.325 51.595 84.495 51.765 ;
      RECT 83.865 51.595 84.035 51.765 ;
      RECT 0.605 51.595 0.775 51.765 ;
      RECT 0.145 51.595 0.315 51.765 ;
      RECT 84.325 48.875 84.495 49.045 ;
      RECT 83.865 48.875 84.035 49.045 ;
      RECT 0.605 48.875 0.775 49.045 ;
      RECT 0.145 48.875 0.315 49.045 ;
      RECT 84.325 46.155 84.495 46.325 ;
      RECT 83.865 46.155 84.035 46.325 ;
      RECT 0.605 46.155 0.775 46.325 ;
      RECT 0.145 46.155 0.315 46.325 ;
      RECT 84.325 43.435 84.495 43.605 ;
      RECT 83.865 43.435 84.035 43.605 ;
      RECT 0.605 43.435 0.775 43.605 ;
      RECT 0.145 43.435 0.315 43.605 ;
      RECT 84.325 40.715 84.495 40.885 ;
      RECT 83.865 40.715 84.035 40.885 ;
      RECT 0.605 40.715 0.775 40.885 ;
      RECT 0.145 40.715 0.315 40.885 ;
      RECT 84.325 37.995 84.495 38.165 ;
      RECT 83.865 37.995 84.035 38.165 ;
      RECT 0.605 37.995 0.775 38.165 ;
      RECT 0.145 37.995 0.315 38.165 ;
      RECT 84.325 35.275 84.495 35.445 ;
      RECT 83.865 35.275 84.035 35.445 ;
      RECT 0.605 35.275 0.775 35.445 ;
      RECT 0.145 35.275 0.315 35.445 ;
      RECT 84.325 32.555 84.495 32.725 ;
      RECT 83.865 32.555 84.035 32.725 ;
      RECT 0.605 32.555 0.775 32.725 ;
      RECT 0.145 32.555 0.315 32.725 ;
      RECT 84.325 29.835 84.495 30.005 ;
      RECT 83.865 29.835 84.035 30.005 ;
      RECT 0.605 29.835 0.775 30.005 ;
      RECT 0.145 29.835 0.315 30.005 ;
      RECT 84.325 27.115 84.495 27.285 ;
      RECT 83.865 27.115 84.035 27.285 ;
      RECT 0.605 27.115 0.775 27.285 ;
      RECT 0.145 27.115 0.315 27.285 ;
      RECT 84.325 24.395 84.495 24.565 ;
      RECT 83.865 24.395 84.035 24.565 ;
      RECT 0.605 24.395 0.775 24.565 ;
      RECT 0.145 24.395 0.315 24.565 ;
      RECT 84.325 21.675 84.495 21.845 ;
      RECT 83.865 21.675 84.035 21.845 ;
      RECT 0.605 21.675 0.775 21.845 ;
      RECT 0.145 21.675 0.315 21.845 ;
      RECT 84.325 18.955 84.495 19.125 ;
      RECT 83.865 18.955 84.035 19.125 ;
      RECT 0.605 18.955 0.775 19.125 ;
      RECT 0.145 18.955 0.315 19.125 ;
      RECT 84.325 16.235 84.495 16.405 ;
      RECT 83.865 16.235 84.035 16.405 ;
      RECT 0.605 16.235 0.775 16.405 ;
      RECT 0.145 16.235 0.315 16.405 ;
      RECT 84.325 13.515 84.495 13.685 ;
      RECT 83.865 13.515 84.035 13.685 ;
      RECT 0.605 13.515 0.775 13.685 ;
      RECT 0.145 13.515 0.315 13.685 ;
      RECT 84.325 10.795 84.495 10.965 ;
      RECT 83.865 10.795 84.035 10.965 ;
      RECT 0.605 10.795 0.775 10.965 ;
      RECT 0.145 10.795 0.315 10.965 ;
      RECT 84.325 8.075 84.495 8.245 ;
      RECT 83.865 8.075 84.035 8.245 ;
      RECT 0.605 8.075 0.775 8.245 ;
      RECT 0.145 8.075 0.315 8.245 ;
      RECT 84.325 5.355 84.495 5.525 ;
      RECT 83.865 5.355 84.035 5.525 ;
      RECT 0.605 5.355 0.775 5.525 ;
      RECT 0.145 5.355 0.315 5.525 ;
      RECT 84.325 2.635 84.495 2.805 ;
      RECT 83.865 2.635 84.035 2.805 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 84.325 -0.085 84.495 0.085 ;
      RECT 83.865 -0.085 84.035 0.085 ;
      RECT 83.405 -0.085 83.575 0.085 ;
      RECT 82.945 -0.085 83.115 0.085 ;
      RECT 82.485 -0.085 82.655 0.085 ;
      RECT 82.025 -0.085 82.195 0.085 ;
      RECT 81.565 -0.085 81.735 0.085 ;
      RECT 81.105 -0.085 81.275 0.085 ;
      RECT 80.645 -0.085 80.815 0.085 ;
      RECT 80.185 -0.085 80.355 0.085 ;
      RECT 79.725 -0.085 79.895 0.085 ;
      RECT 79.265 -0.085 79.435 0.085 ;
      RECT 78.805 -0.085 78.975 0.085 ;
      RECT 78.345 -0.085 78.515 0.085 ;
      RECT 77.885 -0.085 78.055 0.085 ;
      RECT 77.425 -0.085 77.595 0.085 ;
      RECT 76.965 -0.085 77.135 0.085 ;
      RECT 76.505 -0.085 76.675 0.085 ;
      RECT 76.045 -0.085 76.215 0.085 ;
      RECT 75.585 -0.085 75.755 0.085 ;
      RECT 75.125 -0.085 75.295 0.085 ;
      RECT 74.665 -0.085 74.835 0.085 ;
      RECT 74.205 -0.085 74.375 0.085 ;
      RECT 73.745 -0.085 73.915 0.085 ;
      RECT 73.285 -0.085 73.455 0.085 ;
      RECT 72.825 -0.085 72.995 0.085 ;
      RECT 72.365 -0.085 72.535 0.085 ;
      RECT 71.905 -0.085 72.075 0.085 ;
      RECT 71.445 -0.085 71.615 0.085 ;
      RECT 70.985 -0.085 71.155 0.085 ;
      RECT 70.525 -0.085 70.695 0.085 ;
      RECT 70.065 -0.085 70.235 0.085 ;
      RECT 69.605 -0.085 69.775 0.085 ;
      RECT 69.145 -0.085 69.315 0.085 ;
      RECT 68.685 -0.085 68.855 0.085 ;
      RECT 68.225 -0.085 68.395 0.085 ;
      RECT 67.765 -0.085 67.935 0.085 ;
      RECT 67.305 -0.085 67.475 0.085 ;
      RECT 66.845 -0.085 67.015 0.085 ;
      RECT 66.385 -0.085 66.555 0.085 ;
      RECT 65.925 -0.085 66.095 0.085 ;
      RECT 65.465 -0.085 65.635 0.085 ;
      RECT 65.005 -0.085 65.175 0.085 ;
      RECT 64.545 -0.085 64.715 0.085 ;
      RECT 64.085 -0.085 64.255 0.085 ;
      RECT 63.625 -0.085 63.795 0.085 ;
      RECT 63.165 -0.085 63.335 0.085 ;
      RECT 62.705 -0.085 62.875 0.085 ;
      RECT 62.245 -0.085 62.415 0.085 ;
      RECT 61.785 -0.085 61.955 0.085 ;
      RECT 61.325 -0.085 61.495 0.085 ;
      RECT 60.865 -0.085 61.035 0.085 ;
      RECT 60.405 -0.085 60.575 0.085 ;
      RECT 59.945 -0.085 60.115 0.085 ;
      RECT 59.485 -0.085 59.655 0.085 ;
      RECT 59.025 -0.085 59.195 0.085 ;
      RECT 58.565 -0.085 58.735 0.085 ;
      RECT 58.105 -0.085 58.275 0.085 ;
      RECT 57.645 -0.085 57.815 0.085 ;
      RECT 57.185 -0.085 57.355 0.085 ;
      RECT 56.725 -0.085 56.895 0.085 ;
      RECT 56.265 -0.085 56.435 0.085 ;
      RECT 55.805 -0.085 55.975 0.085 ;
      RECT 55.345 -0.085 55.515 0.085 ;
      RECT 54.885 -0.085 55.055 0.085 ;
      RECT 54.425 -0.085 54.595 0.085 ;
      RECT 53.965 -0.085 54.135 0.085 ;
      RECT 53.505 -0.085 53.675 0.085 ;
      RECT 53.045 -0.085 53.215 0.085 ;
      RECT 52.585 -0.085 52.755 0.085 ;
      RECT 52.125 -0.085 52.295 0.085 ;
      RECT 51.665 -0.085 51.835 0.085 ;
      RECT 51.205 -0.085 51.375 0.085 ;
      RECT 50.745 -0.085 50.915 0.085 ;
      RECT 50.285 -0.085 50.455 0.085 ;
      RECT 49.825 -0.085 49.995 0.085 ;
      RECT 49.365 -0.085 49.535 0.085 ;
      RECT 48.905 -0.085 49.075 0.085 ;
      RECT 48.445 -0.085 48.615 0.085 ;
      RECT 47.985 -0.085 48.155 0.085 ;
      RECT 47.525 -0.085 47.695 0.085 ;
      RECT 47.065 -0.085 47.235 0.085 ;
      RECT 46.605 -0.085 46.775 0.085 ;
      RECT 46.145 -0.085 46.315 0.085 ;
      RECT 45.685 -0.085 45.855 0.085 ;
      RECT 45.225 -0.085 45.395 0.085 ;
      RECT 44.765 -0.085 44.935 0.085 ;
      RECT 44.305 -0.085 44.475 0.085 ;
      RECT 43.845 -0.085 44.015 0.085 ;
      RECT 43.385 -0.085 43.555 0.085 ;
      RECT 42.925 -0.085 43.095 0.085 ;
      RECT 42.465 -0.085 42.635 0.085 ;
      RECT 42.005 -0.085 42.175 0.085 ;
      RECT 41.545 -0.085 41.715 0.085 ;
      RECT 41.085 -0.085 41.255 0.085 ;
      RECT 40.625 -0.085 40.795 0.085 ;
      RECT 40.165 -0.085 40.335 0.085 ;
      RECT 39.705 -0.085 39.875 0.085 ;
      RECT 39.245 -0.085 39.415 0.085 ;
      RECT 38.785 -0.085 38.955 0.085 ;
      RECT 38.325 -0.085 38.495 0.085 ;
      RECT 37.865 -0.085 38.035 0.085 ;
      RECT 37.405 -0.085 37.575 0.085 ;
      RECT 36.945 -0.085 37.115 0.085 ;
      RECT 36.485 -0.085 36.655 0.085 ;
      RECT 36.025 -0.085 36.195 0.085 ;
      RECT 35.565 -0.085 35.735 0.085 ;
      RECT 35.105 -0.085 35.275 0.085 ;
      RECT 34.645 -0.085 34.815 0.085 ;
      RECT 34.185 -0.085 34.355 0.085 ;
      RECT 33.725 -0.085 33.895 0.085 ;
      RECT 33.265 -0.085 33.435 0.085 ;
      RECT 32.805 -0.085 32.975 0.085 ;
      RECT 32.345 -0.085 32.515 0.085 ;
      RECT 31.885 -0.085 32.055 0.085 ;
      RECT 31.425 -0.085 31.595 0.085 ;
      RECT 30.965 -0.085 31.135 0.085 ;
      RECT 30.505 -0.085 30.675 0.085 ;
      RECT 30.045 -0.085 30.215 0.085 ;
      RECT 29.585 -0.085 29.755 0.085 ;
      RECT 29.125 -0.085 29.295 0.085 ;
      RECT 28.665 -0.085 28.835 0.085 ;
      RECT 28.205 -0.085 28.375 0.085 ;
      RECT 27.745 -0.085 27.915 0.085 ;
      RECT 27.285 -0.085 27.455 0.085 ;
      RECT 26.825 -0.085 26.995 0.085 ;
      RECT 26.365 -0.085 26.535 0.085 ;
      RECT 25.905 -0.085 26.075 0.085 ;
      RECT 25.445 -0.085 25.615 0.085 ;
      RECT 24.985 -0.085 25.155 0.085 ;
      RECT 24.525 -0.085 24.695 0.085 ;
      RECT 24.065 -0.085 24.235 0.085 ;
      RECT 23.605 -0.085 23.775 0.085 ;
      RECT 23.145 -0.085 23.315 0.085 ;
      RECT 22.685 -0.085 22.855 0.085 ;
      RECT 22.225 -0.085 22.395 0.085 ;
      RECT 21.765 -0.085 21.935 0.085 ;
      RECT 21.305 -0.085 21.475 0.085 ;
      RECT 20.845 -0.085 21.015 0.085 ;
      RECT 20.385 -0.085 20.555 0.085 ;
      RECT 19.925 -0.085 20.095 0.085 ;
      RECT 19.465 -0.085 19.635 0.085 ;
      RECT 19.005 -0.085 19.175 0.085 ;
      RECT 18.545 -0.085 18.715 0.085 ;
      RECT 18.085 -0.085 18.255 0.085 ;
      RECT 17.625 -0.085 17.795 0.085 ;
      RECT 17.165 -0.085 17.335 0.085 ;
      RECT 16.705 -0.085 16.875 0.085 ;
      RECT 16.245 -0.085 16.415 0.085 ;
      RECT 15.785 -0.085 15.955 0.085 ;
      RECT 15.325 -0.085 15.495 0.085 ;
      RECT 14.865 -0.085 15.035 0.085 ;
      RECT 14.405 -0.085 14.575 0.085 ;
      RECT 13.945 -0.085 14.115 0.085 ;
      RECT 13.485 -0.085 13.655 0.085 ;
      RECT 13.025 -0.085 13.195 0.085 ;
      RECT 12.565 -0.085 12.735 0.085 ;
      RECT 12.105 -0.085 12.275 0.085 ;
      RECT 11.645 -0.085 11.815 0.085 ;
      RECT 11.185 -0.085 11.355 0.085 ;
      RECT 10.725 -0.085 10.895 0.085 ;
      RECT 10.265 -0.085 10.435 0.085 ;
      RECT 9.805 -0.085 9.975 0.085 ;
      RECT 9.345 -0.085 9.515 0.085 ;
      RECT 8.885 -0.085 9.055 0.085 ;
      RECT 8.425 -0.085 8.595 0.085 ;
      RECT 7.965 -0.085 8.135 0.085 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.145 -0.085 0.315 0.085 ;
    LAYER via ;
      RECT 56.965 108.725 57.115 108.875 ;
      RECT 27.525 108.725 27.675 108.875 ;
      RECT 30.745 107.025 30.895 107.175 ;
      RECT 13.725 107.025 13.875 107.175 ;
      RECT 72.145 1.625 72.295 1.775 ;
      RECT 62.025 1.625 62.175 1.775 ;
      RECT 51.905 1.625 52.055 1.775 ;
      RECT 56.965 -0.075 57.115 0.075 ;
      RECT 27.525 -0.075 27.675 0.075 ;
    LAYER via2 ;
      RECT 56.94 108.7 57.14 108.9 ;
      RECT 27.5 108.7 27.7 108.9 ;
      RECT 56.94 -0.1 57.14 0.1 ;
      RECT 27.5 -0.1 27.7 0.1 ;
    LAYER via3 ;
      RECT 56.94 108.7 57.14 108.9 ;
      RECT 27.5 108.7 27.7 108.9 ;
      RECT 1.74 3.3 1.94 3.5 ;
      RECT 56.94 -0.1 57.14 0.1 ;
      RECT 27.5 -0.1 27.7 0.1 ;
    LAYER via4 ;
      RECT 71.36 105.8 72.16 106.6 ;
      RECT 41.92 105.8 42.72 106.6 ;
      RECT 12.48 105.8 13.28 106.6 ;
      RECT 56.64 2.2 57.44 3 ;
      RECT 27.2 2.2 28 3 ;
    LAYER fieldpoly ;
      RECT 0.14 0.14 84.5 108.66 ;
    LAYER diff ;
      RECT 0 0 84.64 108.8 ;
    LAYER nwell ;
      POLYGON 84.83 107.495 84.83 104.665 83.99 104.665 83.99 105.89 80.77 105.89 80.77 107.495 ;
      RECT -0.19 104.665 3.87 107.495 ;
      POLYGON 84.83 102.055 84.83 99.225 83.99 99.225 83.99 100.45 83.53 100.45 83.53 102.055 ;
      RECT -0.19 99.225 3.87 102.055 ;
      RECT 83.99 93.785 84.83 96.615 ;
      RECT -0.19 93.785 3.87 96.615 ;
      RECT 83.99 88.345 84.83 91.175 ;
      RECT -0.19 88.345 3.87 91.175 ;
      POLYGON 84.83 85.735 84.83 82.905 83.53 82.905 83.53 84.51 83.99 84.51 83.99 85.735 ;
      RECT -0.19 82.905 2.03 85.735 ;
      RECT 83.53 77.465 84.83 80.295 ;
      POLYGON 2.03 80.295 2.03 79.07 3.87 79.07 3.87 77.465 -0.19 77.465 -0.19 80.295 ;
      POLYGON 84.83 74.855 84.83 72.025 82.61 72.025 82.61 73.25 80.77 73.25 80.77 74.855 ;
      RECT -0.19 72.025 3.87 74.855 ;
      POLYGON 84.83 69.415 84.83 66.585 83.53 66.585 83.53 67.81 82.61 67.81 82.61 69.415 ;
      RECT -0.19 66.585 3.87 69.415 ;
      POLYGON 84.83 63.975 84.83 61.145 83.53 61.145 83.53 62.75 83.99 62.75 83.99 63.975 ;
      RECT -0.19 61.145 3.87 63.975 ;
      POLYGON 84.83 58.535 84.83 55.705 80.77 55.705 80.77 57.31 83.53 57.31 83.53 58.535 ;
      RECT -0.19 55.705 3.87 58.535 ;
      POLYGON 84.83 53.095 84.83 50.265 80.77 50.265 80.77 51.87 83.53 51.87 83.53 53.095 ;
      RECT -0.19 50.265 3.87 53.095 ;
      RECT 80.77 44.825 84.83 47.655 ;
      RECT -0.19 44.825 3.87 47.655 ;
      RECT 80.77 39.385 84.83 42.215 ;
      RECT -0.19 39.385 3.87 42.215 ;
      RECT 80.77 33.945 84.83 36.775 ;
      RECT -0.19 33.945 3.87 36.775 ;
      RECT 80.77 28.505 84.83 31.335 ;
      RECT -0.19 28.505 3.87 31.335 ;
      POLYGON 84.83 25.895 84.83 23.065 82.61 23.065 82.61 24.67 83.53 24.67 83.53 25.895 ;
      RECT -0.19 23.065 3.87 25.895 ;
      POLYGON 84.83 20.455 84.83 17.625 82.61 17.625 82.61 19.23 83.99 19.23 83.99 20.455 ;
      RECT -0.19 17.625 3.87 20.455 ;
      RECT 83.99 12.185 84.83 15.015 ;
      RECT -0.19 12.185 3.87 15.015 ;
      POLYGON 84.83 9.575 84.83 6.745 83.53 6.745 83.53 8.35 83.99 8.35 83.99 9.575 ;
      RECT -0.19 6.745 3.87 9.575 ;
      RECT 80.77 1.305 84.83 4.135 ;
      RECT -0.19 1.305 3.87 4.135 ;
      RECT 0 0 84.64 108.8 ;
    LAYER pwell ;
      RECT 81.09 108.75 81.31 108.92 ;
      RECT 77.41 108.75 77.63 108.92 ;
      RECT 73.73 108.75 73.95 108.92 ;
      RECT 70.05 108.75 70.27 108.92 ;
      RECT 66.37 108.75 66.59 108.92 ;
      RECT 62.69 108.75 62.91 108.92 ;
      RECT 59.01 108.75 59.23 108.92 ;
      RECT 55.33 108.75 55.55 108.92 ;
      RECT 51.65 108.75 51.87 108.92 ;
      RECT 47.97 108.75 48.19 108.92 ;
      RECT 44.29 108.75 44.51 108.92 ;
      RECT 40.61 108.75 40.83 108.92 ;
      RECT 36.93 108.75 37.15 108.92 ;
      RECT 33.25 108.75 33.47 108.92 ;
      RECT 29.57 108.75 29.79 108.92 ;
      RECT 25.89 108.75 26.11 108.92 ;
      RECT 22.21 108.75 22.43 108.92 ;
      RECT 18.53 108.75 18.75 108.92 ;
      RECT 14.85 108.75 15.07 108.92 ;
      RECT 11.17 108.75 11.39 108.92 ;
      RECT 7.49 108.75 7.71 108.92 ;
      RECT 3.81 108.75 4.03 108.92 ;
      RECT 0.13 108.75 0.35 108.92 ;
      RECT 81.09 -0.12 81.31 0.05 ;
      RECT 77.41 -0.12 77.63 0.05 ;
      RECT 73.73 -0.12 73.95 0.05 ;
      RECT 70.05 -0.12 70.27 0.05 ;
      RECT 66.37 -0.12 66.59 0.05 ;
      RECT 62.69 -0.12 62.91 0.05 ;
      RECT 59.01 -0.12 59.23 0.05 ;
      RECT 55.33 -0.12 55.55 0.05 ;
      RECT 51.65 -0.12 51.87 0.05 ;
      RECT 47.97 -0.12 48.19 0.05 ;
      RECT 44.29 -0.12 44.51 0.05 ;
      RECT 40.61 -0.12 40.83 0.05 ;
      RECT 36.93 -0.12 37.15 0.05 ;
      RECT 33.25 -0.12 33.47 0.05 ;
      RECT 29.57 -0.12 29.79 0.05 ;
      RECT 25.89 -0.12 26.11 0.05 ;
      RECT 22.21 -0.12 22.43 0.05 ;
      RECT 18.53 -0.12 18.75 0.05 ;
      RECT 14.85 -0.12 15.07 0.05 ;
      RECT 11.17 -0.12 11.39 0.05 ;
      RECT 7.49 -0.12 7.71 0.05 ;
      RECT 3.81 -0.12 4.03 0.05 ;
      RECT 0.13 -0.12 0.35 0.05 ;
      RECT 0 0 84.64 108.8 ;
    LAYER OVERLAP ;
      POLYGON 0 0 0 108.8 84.64 108.8 84.64 0 ;
  END
END cby_0__1_

END LIBRARY
