//Generated from netlist by SpyDrNet
//netlist name: FPGA88_SOFA_A
module sky130_fd_sc_hd__mux2_1_wrapper
(
    A0,
    A1,
    S,
    X
);

    input A0;
    input A1;
    input S;
    output X;

    wire A0;
    wire A1;
    wire S;
    wire X;

endmodule

