VERSION 5.7 ;
BUSBITCHARS "[]" ;

UNITS
  DATABASE MICRONS 1000 ;
END UNITS

MANUFACTURINGGRID 0.005 ;

LAYER li1
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.46 ;
  WIDTH 0.17 ;
END li1

LAYER mcon
  TYPE CUT ;
END mcon

LAYER met1
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.34 ;
  WIDTH 0.14 ;
END met1

LAYER via
  TYPE CUT ;
END via

LAYER met2
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.46 ;
  WIDTH 0.14 ;
END met2

LAYER via2
  TYPE CUT ;
END via2

LAYER met3
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.68 ;
  WIDTH 0.3 ;
END met3

LAYER via3
  TYPE CUT ;
END via3

LAYER met4
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.92 ;
  WIDTH 0.3 ;
END met4

LAYER via4
  TYPE CUT ;
END via4

LAYER met5
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 3.4 ;
  WIDTH 1.6 ;
END met5

LAYER nwell
  TYPE MASTERSLICE ;
END nwell

LAYER pwell
  TYPE MASTERSLICE ;
END pwell

LAYER OVERLAP
  TYPE OVERLAP ;
END OVERLAP

VIA L1M1_PR
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.145 -0.115 0.145 0.115 ;
END L1M1_PR

VIA L1M1_PR_R
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.115 -0.145 0.115 0.145 ;
END L1M1_PR_R

VIA L1M1_PR_M
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.115 -0.145 0.115 0.145 ;
END L1M1_PR_M

VIA L1M1_PR_MR
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.145 -0.115 0.145 0.115 ;
END L1M1_PR_MR

VIA L1M1_PR_C
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.145 -0.145 0.145 0.145 ;
END L1M1_PR_C

VIA M1M2_PR
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR

VIA M1M2_PR_Enc
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_Enc

VIA M1M2_PR_R
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_R

VIA M1M2_PR_R_Enc
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR_R_Enc

VIA M1M2_PR_M
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_M

VIA M1M2_PR_M_Enc
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR_M_Enc

VIA M1M2_PR_MR
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR_MR

VIA M1M2_PR_MR_Enc
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_MR_Enc

VIA M1M2_PR_C
  LAYER met1 ;
    RECT -0.16 -0.16 0.16 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.16 0.16 0.16 ;
END M1M2_PR_C

VIA M2M3_PR
  LAYER met2 ;
    RECT -0.14 -0.185 0.14 0.185 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR

VIA M2M3_PR_R
  LAYER met2 ;
    RECT -0.185 -0.14 0.185 0.14 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_R

VIA M2M3_PR_M
  LAYER met2 ;
    RECT -0.14 -0.185 0.14 0.185 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_M

VIA M2M3_PR_MR
  LAYER met2 ;
    RECT -0.185 -0.14 0.185 0.14 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_MR

VIA M2M3_PR_C
  LAYER met2 ;
    RECT -0.185 -0.185 0.185 0.185 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_C

VIA M3M4_PR
  LAYER met3 ;
    RECT -0.19 -0.16 0.19 0.16 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR

VIA M3M4_PR_R
  LAYER met3 ;
    RECT -0.16 -0.19 0.16 0.19 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_R

VIA M3M4_PR_M
  LAYER met3 ;
    RECT -0.19 -0.16 0.19 0.16 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_M

VIA M3M4_PR_MR
  LAYER met3 ;
    RECT -0.16 -0.19 0.16 0.19 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_MR

VIA M3M4_PR_C
  LAYER met3 ;
    RECT -0.19 -0.19 0.19 0.19 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_C

VIA M4M5_PR
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR

VIA M4M5_PR_R
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_R

VIA M4M5_PR_M
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_M

VIA M4M5_PR_MR
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_MR

VIA M4M5_PR_C
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_C

SITE unit
  CLASS CORE ;
  SYMMETRY Y ;
  SIZE 0.46 BY 2.72 ;
END unit

SITE unithddbl
  CLASS CORE ;
  SIZE 0.46 BY 5.44 ;
END unithddbl

MACRO sb_0__1_
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  SIZE 95.68 BY 108.8 ;
  SYMMETRY X Y ;
  PIN prog_clk[0]
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER met2 ;
        RECT 83.65 10.88 83.79 12.24 ;
    END
  END prog_clk[0]
  PIN chany_top_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.33 107.44 41.47 108.8 ;
    END
  END chany_top_in[0]
  PIN chany_top_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.11 107.44 61.25 108.8 ;
    END
  END chany_top_in[1]
  PIN chany_top_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.37 107.44 52.51 108.8 ;
    END
  END chany_top_in[2]
  PIN chany_top_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.19 107.44 60.33 108.8 ;
    END
  END chany_top_in[3]
  PIN chany_top_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.55 107.44 44.69 108.8 ;
    END
  END chany_top_in[4]
  PIN chany_top_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.03 107.44 62.17 108.8 ;
    END
  END chany_top_in[5]
  PIN chany_top_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.33 107.44 18.47 108.8 ;
    END
  END chany_top_in[6]
  PIN chany_top_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.41 107.44 40.55 108.8 ;
    END
  END chany_top_in[7]
  PIN chany_top_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.49 107.44 39.63 108.8 ;
    END
  END chany_top_in[8]
  PIN chany_top_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 17.33 107.44 17.63 108.8 ;
    END
  END chany_top_in[9]
  PIN chany_top_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 54.13 107.44 54.43 108.8 ;
    END
  END chany_top_in[10]
  PIN chany_top_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.43 107.44 57.57 108.8 ;
    END
  END chany_top_in[11]
  PIN chany_top_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.21 107.44 54.35 108.8 ;
    END
  END chany_top_in[12]
  PIN chany_top_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.95 107.44 63.09 108.8 ;
    END
  END chany_top_in[13]
  PIN chany_top_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.73 107.44 13.87 108.8 ;
    END
  END chany_top_in[14]
  PIN chany_top_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.41 107.44 17.55 108.8 ;
    END
  END chany_top_in[15]
  PIN chany_top_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.97 107.44 34.11 108.8 ;
    END
  END chany_top_in[16]
  PIN chany_top_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 63.33 107.44 63.63 108.8 ;
    END
  END chany_top_in[17]
  PIN chany_top_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 33.89 107.44 34.19 108.8 ;
    END
  END chany_top_in[18]
  PIN chany_top_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.89 107.44 35.03 108.8 ;
    END
  END chany_top_in[19]
  PIN top_left_grid_pin_1_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.45 107.44 51.59 108.8 ;
    END
  END top_left_grid_pin_1_[0]
  PIN chanx_right_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 94.3 37.25 95.68 37.55 ;
    END
  END chanx_right_in[0]
  PIN chanx_right_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 94.3 71.25 95.68 71.55 ;
    END
  END chanx_right_in[1]
  PIN chanx_right_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 94.3 92.33 95.68 92.63 ;
    END
  END chanx_right_in[2]
  PIN chanx_right_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 94.3 84.85 95.68 85.15 ;
    END
  END chanx_right_in[3]
  PIN chanx_right_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 94.3 73.97 95.68 74.27 ;
    END
  END chanx_right_in[4]
  PIN chanx_right_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 94.3 76.69 95.68 76.99 ;
    END
  END chanx_right_in[5]
  PIN chanx_right_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 94.3 67.17 95.68 67.47 ;
    END
  END chanx_right_in[6]
  PIN chanx_right_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 94.3 39.97 95.68 40.27 ;
    END
  END chanx_right_in[7]
  PIN chanx_right_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 94.3 55.61 95.68 55.91 ;
    END
  END chanx_right_in[8]
  PIN chanx_right_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 94.3 75.33 95.68 75.63 ;
    END
  END chanx_right_in[9]
  PIN chanx_right_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 94.3 59.69 95.68 59.99 ;
    END
  END chanx_right_in[10]
  PIN chanx_right_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 94.3 72.61 95.68 72.91 ;
    END
  END chanx_right_in[11]
  PIN chanx_right_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 94.3 78.05 95.68 78.35 ;
    END
  END chanx_right_in[12]
  PIN chanx_right_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 94.3 35.89 95.68 36.19 ;
    END
  END chanx_right_in[13]
  PIN chanx_right_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 94.3 31.81 95.68 32.11 ;
    END
  END chanx_right_in[14]
  PIN chanx_right_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 94.3 41.33 95.68 41.63 ;
    END
  END chanx_right_in[15]
  PIN chanx_right_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 94.3 89.61 95.68 89.91 ;
    END
  END chanx_right_in[16]
  PIN chanx_right_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 94.3 44.05 95.68 44.35 ;
    END
  END chanx_right_in[17]
  PIN chanx_right_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 94.3 80.77 95.68 81.07 ;
    END
  END chanx_right_in[18]
  PIN chanx_right_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 94.3 38.61 95.68 38.91 ;
    END
  END chanx_right_in[19]
  PIN right_bottom_grid_pin_34_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.33 10.88 87.47 12.24 ;
    END
  END right_bottom_grid_pin_34_[0]
  PIN right_bottom_grid_pin_35_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.25 10.88 88.39 12.24 ;
    END
  END right_bottom_grid_pin_35_[0]
  PIN right_bottom_grid_pin_36_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.27 10.88 82.41 12.24 ;
    END
  END right_bottom_grid_pin_36_[0]
  PIN right_bottom_grid_pin_37_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.03 10.88 85.17 12.24 ;
    END
  END right_bottom_grid_pin_37_[0]
  PIN right_bottom_grid_pin_38_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.01 10.88 91.15 12.24 ;
    END
  END right_bottom_grid_pin_38_[0]
  PIN right_bottom_grid_pin_39_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.17 10.88 89.31 12.24 ;
    END
  END right_bottom_grid_pin_39_[0]
  PIN right_bottom_grid_pin_40_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.09 10.88 90.23 12.24 ;
    END
  END right_bottom_grid_pin_40_[0]
  PIN right_bottom_grid_pin_41_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.41 10.88 86.55 12.24 ;
    END
  END right_bottom_grid_pin_41_[0]
  PIN chany_bottom_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.91 0 52.05 1.36 ;
    END
  END chany_bottom_in[0]
  PIN chany_bottom_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.23 0 48.37 1.36 ;
    END
  END chany_bottom_in[1]
  PIN chany_bottom_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.87 0 64.01 1.36 ;
    END
  END chany_bottom_in[2]
  PIN chany_bottom_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.03 0 62.17 1.36 ;
    END
  END chany_bottom_in[3]
  PIN chany_bottom_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.39 0 46.53 1.36 ;
    END
  END chany_bottom_in[4]
  PIN chany_bottom_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.55 0 44.69 1.36 ;
    END
  END chany_bottom_in[5]
  PIN chany_bottom_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.25 0 19.39 1.36 ;
    END
  END chany_bottom_in[6]
  PIN chany_bottom_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.43 0 34.57 1.36 ;
    END
  END chany_bottom_in[7]
  PIN chany_bottom_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.81 0 12.95 1.36 ;
    END
  END chany_bottom_in[8]
  PIN chany_bottom_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.33 0 18.47 1.36 ;
    END
  END chany_bottom_in[9]
  PIN chany_bottom_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.77 0 24.91 1.36 ;
    END
  END chany_bottom_in[10]
  PIN chany_bottom_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.59 0 32.73 1.36 ;
    END
  END chany_bottom_in[11]
  PIN chany_bottom_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.47 0 45.61 1.36 ;
    END
  END chany_bottom_in[12]
  PIN chany_bottom_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.51 0 33.65 1.36 ;
    END
  END chany_bottom_in[13]
  PIN chany_bottom_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.87 0 41.01 1.36 ;
    END
  END chany_bottom_in[14]
  PIN chany_bottom_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.73 0 13.87 1.36 ;
    END
  END chany_bottom_in[15]
  PIN chany_bottom_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.69 0 25.83 1.36 ;
    END
  END chany_bottom_in[16]
  PIN chany_bottom_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.97 0 11.11 1.36 ;
    END
  END chany_bottom_in[17]
  PIN chany_bottom_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.89 0 12.03 1.36 ;
    END
  END chany_bottom_in[18]
  PIN chany_bottom_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.05 0 10.19 1.36 ;
    END
  END chany_bottom_in[19]
  PIN bottom_left_grid_pin_1_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.99 0 51.13 1.36 ;
    END
  END bottom_left_grid_pin_1_[0]
  PIN ccff_head[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 94.3 86.89 95.68 87.19 ;
    END
  END ccff_head[0]
  PIN chany_top_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.29 107.44 53.43 108.8 ;
    END
  END chany_top_out[0]
  PIN chany_top_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.65 107.44 14.79 108.8 ;
    END
  END chany_top_out[1]
  PIN chany_top_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.71 107.44 65.85 108.8 ;
    END
  END chany_top_out[2]
  PIN chany_top_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.49 107.44 16.63 108.8 ;
    END
  END chany_top_out[3]
  PIN chany_top_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.33 107.44 64.47 108.8 ;
    END
  END chany_top_out[4]
  PIN chany_top_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.81 107.44 35.95 108.8 ;
    END
  END chany_top_out[5]
  PIN chany_top_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.57 107.44 38.71 108.8 ;
    END
  END chany_top_out[6]
  PIN chany_top_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.73 107.44 36.87 108.8 ;
    END
  END chany_top_out[7]
  PIN chany_top_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.57 107.44 15.71 108.8 ;
    END
  END chany_top_out[8]
  PIN chany_top_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.65 107.44 37.79 108.8 ;
    END
  END chany_top_out[9]
  PIN chany_top_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.13 107.44 55.27 108.8 ;
    END
  END chany_top_out[10]
  PIN chany_top_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 61.49 107.44 61.79 108.8 ;
    END
  END chany_top_out[11]
  PIN chany_top_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.35 107.44 58.49 108.8 ;
    END
  END chany_top_out[12]
  PIN chany_top_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 39.41 107.44 39.71 108.8 ;
    END
  END chany_top_out[13]
  PIN chany_top_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 15.49 107.44 15.79 108.8 ;
    END
  END chany_top_out[14]
  PIN chany_top_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 35.73 107.44 36.03 108.8 ;
    END
  END chany_top_out[15]
  PIN chany_top_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.27 107.44 59.41 108.8 ;
    END
  END chany_top_out[16]
  PIN chany_top_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 59.65 107.44 59.95 108.8 ;
    END
  END chany_top_out[17]
  PIN chany_top_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 57.81 107.44 58.11 108.8 ;
    END
  END chany_top_out[18]
  PIN chany_top_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 37.57 107.44 37.87 108.8 ;
    END
  END chany_top_out[19]
  PIN chanx_right_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 94.3 83.49 95.68 83.79 ;
    END
  END chanx_right_out[0]
  PIN chanx_right_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 94.3 90.97 95.68 91.27 ;
    END
  END chanx_right_out[1]
  PIN chanx_right_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 94.3 48.13 95.68 48.43 ;
    END
  END chanx_right_out[2]
  PIN chanx_right_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 94.3 61.05 95.68 61.35 ;
    END
  END chanx_right_out[3]
  PIN chanx_right_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 94.3 82.13 95.68 82.43 ;
    END
  END chanx_right_out[4]
  PIN chanx_right_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 94.3 79.41 95.68 79.71 ;
    END
  END chanx_right_out[5]
  PIN chanx_right_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 94.3 54.25 95.68 54.55 ;
    END
  END chanx_right_out[6]
  PIN chanx_right_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 94.3 64.45 95.68 64.75 ;
    END
  END chanx_right_out[7]
  PIN chanx_right_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 94.3 56.97 95.68 57.27 ;
    END
  END chanx_right_out[8]
  PIN chanx_right_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 94.3 50.85 95.68 51.15 ;
    END
  END chanx_right_out[9]
  PIN chanx_right_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 94.3 49.49 95.68 49.79 ;
    END
  END chanx_right_out[10]
  PIN chanx_right_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 94.3 65.81 95.68 66.11 ;
    END
  END chanx_right_out[11]
  PIN chanx_right_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 94.3 45.41 95.68 45.71 ;
    END
  END chanx_right_out[12]
  PIN chanx_right_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 94.3 88.25 95.68 88.55 ;
    END
  END chanx_right_out[13]
  PIN chanx_right_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 94.3 46.77 95.68 47.07 ;
    END
  END chanx_right_out[14]
  PIN chanx_right_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 94.3 42.69 95.68 42.99 ;
    END
  END chanx_right_out[15]
  PIN chanx_right_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 94.3 58.33 95.68 58.63 ;
    END
  END chanx_right_out[16]
  PIN chanx_right_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 94.3 52.89 95.68 53.19 ;
    END
  END chanx_right_out[17]
  PIN chanx_right_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 94.3 62.41 95.68 62.71 ;
    END
  END chanx_right_out[18]
  PIN chanx_right_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 94.3 69.21 95.68 69.51 ;
    END
  END chanx_right_out[19]
  PIN chany_bottom_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.75 0 53.89 1.36 ;
    END
  END chany_bottom_out[0]
  PIN chany_bottom_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.13 0 55.27 1.36 ;
    END
  END chany_bottom_out[1]
  PIN chany_bottom_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.25 0 65.39 1.36 ;
    END
  END chany_bottom_out[2]
  PIN chany_bottom_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.11 0 61.25 1.36 ;
    END
  END chany_bottom_out[3]
  PIN chany_bottom_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.83 0 52.97 1.36 ;
    END
  END chany_bottom_out[4]
  PIN chany_bottom_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.41 0 17.55 1.36 ;
    END
  END chany_bottom_out[5]
  PIN chany_bottom_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.95 0 40.09 1.36 ;
    END
  END chany_bottom_out[6]
  PIN chany_bottom_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.19 0 60.33 1.36 ;
    END
  END chany_bottom_out[7]
  PIN chany_bottom_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.27 0 59.41 1.36 ;
    END
  END chany_bottom_out[8]
  PIN chany_bottom_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.35 0 35.49 1.36 ;
    END
  END chany_bottom_out[9]
  PIN chany_bottom_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.95 0 63.09 1.36 ;
    END
  END chany_bottom_out[10]
  PIN chany_bottom_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.03 0 39.17 1.36 ;
    END
  END chany_bottom_out[11]
  PIN chany_bottom_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.79 0 41.93 1.36 ;
    END
  END chany_bottom_out[12]
  PIN chany_bottom_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.65 0 14.79 1.36 ;
    END
  END chany_bottom_out[13]
  PIN chany_bottom_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.49 0 16.63 1.36 ;
    END
  END chany_bottom_out[14]
  PIN chany_bottom_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.27 0 36.41 1.36 ;
    END
  END chany_bottom_out[15]
  PIN chany_bottom_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.63 0 43.77 1.36 ;
    END
  END chany_bottom_out[16]
  PIN chany_bottom_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.43 0 57.57 1.36 ;
    END
  END chany_bottom_out[17]
  PIN chany_bottom_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.57 0 15.71 1.36 ;
    END
  END chany_bottom_out[18]
  PIN chany_bottom_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.35 0 58.49 1.36 ;
    END
  END chany_bottom_out[19]
  PIN ccff_tail[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.71 0 42.85 1.36 ;
    END
  END ccff_tail[0]
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0 2.48 0.48 2.96 ;
        RECT 67.6 2.48 68.08 2.96 ;
        RECT 0 7.92 0.48 8.4 ;
        RECT 67.6 7.92 68.08 8.4 ;
        RECT 0 13.36 0.48 13.84 ;
        RECT 95.2 13.36 95.68 13.84 ;
        RECT 0 18.8 0.48 19.28 ;
        RECT 95.2 18.8 95.68 19.28 ;
        RECT 0 24.24 0.48 24.72 ;
        RECT 95.2 24.24 95.68 24.72 ;
        RECT 0 29.68 0.48 30.16 ;
        RECT 95.2 29.68 95.68 30.16 ;
        RECT 0 35.12 0.48 35.6 ;
        RECT 95.2 35.12 95.68 35.6 ;
        RECT 0 40.56 0.48 41.04 ;
        RECT 95.2 40.56 95.68 41.04 ;
        RECT 0 46 0.48 46.48 ;
        RECT 95.2 46 95.68 46.48 ;
        RECT 0 51.44 0.48 51.92 ;
        RECT 95.2 51.44 95.68 51.92 ;
        RECT 0 56.88 0.48 57.36 ;
        RECT 95.2 56.88 95.68 57.36 ;
        RECT 0 62.32 0.48 62.8 ;
        RECT 95.2 62.32 95.68 62.8 ;
        RECT 0 67.76 0.48 68.24 ;
        RECT 95.2 67.76 95.68 68.24 ;
        RECT 0 73.2 0.48 73.68 ;
        RECT 95.2 73.2 95.68 73.68 ;
        RECT 0 78.64 0.48 79.12 ;
        RECT 95.2 78.64 95.68 79.12 ;
        RECT 0 84.08 0.48 84.56 ;
        RECT 95.2 84.08 95.68 84.56 ;
        RECT 0 89.52 0.48 90 ;
        RECT 95.2 89.52 95.68 90 ;
        RECT 0 94.96 0.48 95.44 ;
        RECT 95.2 94.96 95.68 95.44 ;
        RECT 0 100.4 0.48 100.88 ;
        RECT 67.6 100.4 68.08 100.88 ;
        RECT 0 105.84 0.48 106.32 ;
        RECT 67.6 105.84 68.08 106.32 ;
      LAYER met4 ;
        RECT 11.66 0 12.26 0.6 ;
        RECT 41.1 0 41.7 0.6 ;
        RECT 85.26 10.88 85.86 11.48 ;
        RECT 85.26 97.32 85.86 97.92 ;
        RECT 11.66 108.2 12.26 108.8 ;
        RECT 41.1 108.2 41.7 108.8 ;
      LAYER met5 ;
        RECT 0 22.2 3.2 25.4 ;
        RECT 92.48 22.2 95.68 25.4 ;
        RECT 0 63 3.2 66.2 ;
        RECT 92.48 63 95.68 66.2 ;
    END
  END VDD
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0 0 68.08 0.24 ;
        RECT 0 5.2 0.48 5.68 ;
        RECT 67.6 5.2 68.08 5.68 ;
        RECT 0 10.64 95.68 11.12 ;
        RECT 0 16.08 0.48 16.56 ;
        RECT 95.2 16.08 95.68 16.56 ;
        RECT 0 21.52 0.48 22 ;
        RECT 95.2 21.52 95.68 22 ;
        RECT 0 26.96 0.48 27.44 ;
        RECT 95.2 26.96 95.68 27.44 ;
        RECT 0 32.4 0.48 32.88 ;
        RECT 95.2 32.4 95.68 32.88 ;
        RECT 0 37.84 0.48 38.32 ;
        RECT 95.2 37.84 95.68 38.32 ;
        RECT 0 43.28 0.48 43.76 ;
        RECT 95.2 43.28 95.68 43.76 ;
        RECT 0 48.72 0.48 49.2 ;
        RECT 95.2 48.72 95.68 49.2 ;
        RECT 0 54.16 0.48 54.64 ;
        RECT 95.2 54.16 95.68 54.64 ;
        RECT 0 59.6 0.48 60.08 ;
        RECT 95.2 59.6 95.68 60.08 ;
        RECT 0 65.04 0.48 65.52 ;
        RECT 95.2 65.04 95.68 65.52 ;
        RECT 0 70.48 0.48 70.96 ;
        RECT 95.2 70.48 95.68 70.96 ;
        RECT 0 75.92 0.48 76.4 ;
        RECT 95.2 75.92 95.68 76.4 ;
        RECT 0 81.36 0.48 81.84 ;
        RECT 95.2 81.36 95.68 81.84 ;
        RECT 0 86.8 0.48 87.28 ;
        RECT 95.2 86.8 95.68 87.28 ;
        RECT 0 92.24 0.48 92.72 ;
        RECT 95.2 92.24 95.68 92.72 ;
        RECT 0 97.68 95.68 98.16 ;
        RECT 0 103.12 0.48 103.6 ;
        RECT 67.6 103.12 68.08 103.6 ;
        RECT 0 108.56 68.08 108.8 ;
      LAYER met4 ;
        RECT 26.38 0 26.98 0.6 ;
        RECT 55.82 0 56.42 0.6 ;
        RECT 26.38 108.2 26.98 108.8 ;
        RECT 55.82 108.2 56.42 108.8 ;
      LAYER met5 ;
        RECT 0 42.6 3.2 45.8 ;
        RECT 92.48 42.6 95.68 45.8 ;
        RECT 0 83.4 3.2 86.6 ;
        RECT 92.48 83.4 95.68 86.6 ;
    END
  END VSS
  PIN prog_clk__FEEDTHRU_1[0]
    DIRECTION OUTPUT ;
    USE CLOCK ;
    PORT
      LAYER met2 ;
        RECT 75.37 96.56 75.51 97.92 ;
    END
  END prog_clk__FEEDTHRU_1[0]
  OBS
    LAYER li1 ;
      RECT 0 108.715 68.08 108.885 ;
      RECT 67.16 105.995 68.08 106.165 ;
      RECT 0 105.995 3.68 106.165 ;
      RECT 67.16 103.275 68.08 103.445 ;
      RECT 0 103.275 3.68 103.445 ;
      RECT 67.16 100.555 68.08 100.725 ;
      RECT 0 100.555 3.68 100.725 ;
      RECT 65.32 97.835 95.68 98.005 ;
      RECT 0 97.835 3.68 98.005 ;
      RECT 95.22 95.115 95.68 95.285 ;
      RECT 0 95.115 3.68 95.285 ;
      RECT 95.22 92.395 95.68 92.565 ;
      RECT 0 92.395 3.68 92.565 ;
      RECT 95.22 89.675 95.68 89.845 ;
      RECT 0 89.675 3.68 89.845 ;
      RECT 94.76 86.955 95.68 87.125 ;
      RECT 0 86.955 3.68 87.125 ;
      RECT 94.76 84.235 95.68 84.405 ;
      RECT 0 84.235 3.68 84.405 ;
      RECT 94.76 81.515 95.68 81.685 ;
      RECT 0 81.515 3.68 81.685 ;
      RECT 94.76 78.795 95.68 78.965 ;
      RECT 0 78.795 3.68 78.965 ;
      RECT 94.76 76.075 95.68 76.245 ;
      RECT 0 76.075 3.68 76.245 ;
      RECT 94.76 73.355 95.68 73.525 ;
      RECT 0 73.355 3.68 73.525 ;
      RECT 94.76 70.635 95.68 70.805 ;
      RECT 0 70.635 3.68 70.805 ;
      RECT 95.22 67.915 95.68 68.085 ;
      RECT 0 67.915 3.68 68.085 ;
      RECT 94.76 65.195 95.68 65.365 ;
      RECT 0 65.195 3.68 65.365 ;
      RECT 94.76 62.475 95.68 62.645 ;
      RECT 0 62.475 3.68 62.645 ;
      RECT 94.76 59.755 95.68 59.925 ;
      RECT 0 59.755 3.68 59.925 ;
      RECT 94.76 57.035 95.68 57.205 ;
      RECT 0 57.035 3.68 57.205 ;
      RECT 94.76 54.315 95.68 54.485 ;
      RECT 0 54.315 3.68 54.485 ;
      RECT 94.76 51.595 95.68 51.765 ;
      RECT 0 51.595 3.68 51.765 ;
      RECT 94.76 48.875 95.68 49.045 ;
      RECT 0 48.875 3.68 49.045 ;
      RECT 94.76 46.155 95.68 46.325 ;
      RECT 0 46.155 3.68 46.325 ;
      RECT 94.76 43.435 95.68 43.605 ;
      RECT 0 43.435 3.68 43.605 ;
      RECT 94.76 40.715 95.68 40.885 ;
      RECT 0 40.715 3.68 40.885 ;
      RECT 95.22 37.995 95.68 38.165 ;
      RECT 0 37.995 3.68 38.165 ;
      RECT 95.22 35.275 95.68 35.445 ;
      RECT 0 35.275 3.68 35.445 ;
      RECT 95.22 32.555 95.68 32.725 ;
      RECT 0 32.555 3.68 32.725 ;
      RECT 95.22 29.835 95.68 30.005 ;
      RECT 0 29.835 3.68 30.005 ;
      RECT 95.22 27.115 95.68 27.285 ;
      RECT 0 27.115 3.68 27.285 ;
      RECT 92 24.395 95.68 24.565 ;
      RECT 0 24.395 3.68 24.565 ;
      RECT 92 21.675 95.68 21.845 ;
      RECT 0 21.675 3.68 21.845 ;
      RECT 92 18.955 95.68 19.125 ;
      RECT 0 18.955 3.68 19.125 ;
      RECT 92 16.235 95.68 16.405 ;
      RECT 0 16.235 3.68 16.405 ;
      RECT 94.76 13.515 95.68 13.685 ;
      RECT 0 13.515 3.68 13.685 ;
      RECT 65.32 10.795 95.68 10.965 ;
      RECT 0 10.795 3.68 10.965 ;
      RECT 67.16 8.075 68.08 8.245 ;
      RECT 0 8.075 3.68 8.245 ;
      RECT 67.16 5.355 68.08 5.525 ;
      RECT 0 5.355 3.68 5.525 ;
      RECT 67.16 2.635 68.08 2.805 ;
      RECT 0 2.635 3.68 2.805 ;
      RECT 0 -0.085 68.08 0.085 ;
    LAYER met2 ;
      RECT 55.98 108.615 56.26 108.985 ;
      RECT 26.54 108.615 26.82 108.985 ;
      RECT 58.75 106.94 59.01 107.26 ;
      RECT 51.85 106.94 52.11 107.26 ;
      RECT 64.73 1.54 64.99 1.86 ;
      RECT 56.91 1.54 57.17 1.86 ;
      RECT 48.63 1.54 48.89 1.86 ;
      RECT 55.98 -0.185 56.26 0.185 ;
      RECT 26.54 -0.185 26.82 0.185 ;
      POLYGON 67.8 108.52 67.8 97.64 75.09 97.64 75.09 96.28 75.79 96.28 75.79 97.64 95.4 97.64 95.4 11.16 91.43 11.16 91.43 12.52 90.73 12.52 90.73 11.16 90.51 11.16 90.51 12.52 89.81 12.52 89.81 11.16 89.59 11.16 89.59 12.52 88.89 12.52 88.89 11.16 88.67 11.16 88.67 12.52 87.97 12.52 87.97 11.16 87.75 11.16 87.75 12.52 87.05 12.52 87.05 11.16 86.83 11.16 86.83 12.52 86.13 12.52 86.13 11.16 85.45 11.16 85.45 12.52 84.75 12.52 84.75 11.16 84.07 11.16 84.07 12.52 83.37 12.52 83.37 11.16 82.69 11.16 82.69 12.52 81.99 12.52 81.99 11.16 67.8 11.16 67.8 0.28 65.67 0.28 65.67 1.64 64.97 1.64 64.97 0.28 64.29 0.28 64.29 1.64 63.59 1.64 63.59 0.28 63.37 0.28 63.37 1.64 62.67 1.64 62.67 0.28 62.45 0.28 62.45 1.64 61.75 1.64 61.75 0.28 61.53 0.28 61.53 1.64 60.83 1.64 60.83 0.28 60.61 0.28 60.61 1.64 59.91 1.64 59.91 0.28 59.69 0.28 59.69 1.64 58.99 1.64 58.99 0.28 58.77 0.28 58.77 1.64 58.07 1.64 58.07 0.28 57.85 0.28 57.85 1.64 57.15 1.64 57.15 0.28 55.55 0.28 55.55 1.64 54.85 1.64 54.85 0.28 54.17 0.28 54.17 1.64 53.47 1.64 53.47 0.28 53.25 0.28 53.25 1.64 52.55 1.64 52.55 0.28 52.33 0.28 52.33 1.64 51.63 1.64 51.63 0.28 51.41 0.28 51.41 1.64 50.71 1.64 50.71 0.28 48.65 0.28 48.65 1.64 47.95 1.64 47.95 0.28 46.81 0.28 46.81 1.64 46.11 1.64 46.11 0.28 45.89 0.28 45.89 1.64 45.19 1.64 45.19 0.28 44.97 0.28 44.97 1.64 44.27 1.64 44.27 0.28 44.05 0.28 44.05 1.64 43.35 1.64 43.35 0.28 43.13 0.28 43.13 1.64 42.43 1.64 42.43 0.28 42.21 0.28 42.21 1.64 41.51 1.64 41.51 0.28 41.29 0.28 41.29 1.64 40.59 1.64 40.59 0.28 40.37 0.28 40.37 1.64 39.67 1.64 39.67 0.28 39.45 0.28 39.45 1.64 38.75 1.64 38.75 0.28 36.69 0.28 36.69 1.64 35.99 1.64 35.99 0.28 35.77 0.28 35.77 1.64 35.07 1.64 35.07 0.28 34.85 0.28 34.85 1.64 34.15 1.64 34.15 0.28 33.93 0.28 33.93 1.64 33.23 1.64 33.23 0.28 33.01 0.28 33.01 1.64 32.31 1.64 32.31 0.28 26.11 0.28 26.11 1.64 25.41 1.64 25.41 0.28 25.19 0.28 25.19 1.64 24.49 1.64 24.49 0.28 19.67 0.28 19.67 1.64 18.97 1.64 18.97 0.28 18.75 0.28 18.75 1.64 18.05 1.64 18.05 0.28 17.83 0.28 17.83 1.64 17.13 1.64 17.13 0.28 16.91 0.28 16.91 1.64 16.21 1.64 16.21 0.28 15.99 0.28 15.99 1.64 15.29 1.64 15.29 0.28 15.07 0.28 15.07 1.64 14.37 1.64 14.37 0.28 14.15 0.28 14.15 1.64 13.45 1.64 13.45 0.28 13.23 0.28 13.23 1.64 12.53 1.64 12.53 0.28 12.31 0.28 12.31 1.64 11.61 1.64 11.61 0.28 11.39 0.28 11.39 1.64 10.69 1.64 10.69 0.28 10.47 0.28 10.47 1.64 9.77 1.64 9.77 0.28 0.28 0.28 0.28 108.52 13.45 108.52 13.45 107.16 14.15 107.16 14.15 108.52 14.37 108.52 14.37 107.16 15.07 107.16 15.07 108.52 15.29 108.52 15.29 107.16 15.99 107.16 15.99 108.52 16.21 108.52 16.21 107.16 16.91 107.16 16.91 108.52 17.13 108.52 17.13 107.16 17.83 107.16 17.83 108.52 18.05 108.52 18.05 107.16 18.75 107.16 18.75 108.52 33.69 108.52 33.69 107.16 34.39 107.16 34.39 108.52 34.61 108.52 34.61 107.16 35.31 107.16 35.31 108.52 35.53 108.52 35.53 107.16 36.23 107.16 36.23 108.52 36.45 108.52 36.45 107.16 37.15 107.16 37.15 108.52 37.37 108.52 37.37 107.16 38.07 107.16 38.07 108.52 38.29 108.52 38.29 107.16 38.99 107.16 38.99 108.52 39.21 108.52 39.21 107.16 39.91 107.16 39.91 108.52 40.13 108.52 40.13 107.16 40.83 107.16 40.83 108.52 41.05 108.52 41.05 107.16 41.75 107.16 41.75 108.52 44.27 108.52 44.27 107.16 44.97 107.16 44.97 108.52 51.17 108.52 51.17 107.16 51.87 107.16 51.87 108.52 52.09 108.52 52.09 107.16 52.79 107.16 52.79 108.52 53.01 108.52 53.01 107.16 53.71 107.16 53.71 108.52 53.93 108.52 53.93 107.16 54.63 107.16 54.63 108.52 54.85 108.52 54.85 107.16 55.55 107.16 55.55 108.52 57.15 108.52 57.15 107.16 57.85 107.16 57.85 108.52 58.07 108.52 58.07 107.16 58.77 107.16 58.77 108.52 58.99 108.52 58.99 107.16 59.69 107.16 59.69 108.52 59.91 108.52 59.91 107.16 60.61 107.16 60.61 108.52 60.83 108.52 60.83 107.16 61.53 107.16 61.53 108.52 61.75 108.52 61.75 107.16 62.45 107.16 62.45 108.52 62.67 108.52 62.67 107.16 63.37 107.16 63.37 108.52 64.05 108.52 64.05 107.16 64.75 107.16 64.75 108.52 65.43 108.52 65.43 107.16 66.13 107.16 66.13 108.52 ;
    LAYER met4 ;
      POLYGON 67.68 108.4 67.68 97.52 84.86 97.52 84.86 96.92 86.26 96.92 86.26 97.52 95.28 97.52 95.28 11.28 86.26 11.28 86.26 11.88 84.86 11.88 84.86 11.28 67.68 11.28 67.68 0.4 56.82 0.4 56.82 1 55.42 1 55.42 0.4 42.1 0.4 42.1 1 40.7 1 40.7 0.4 27.38 0.4 27.38 1 25.98 1 25.98 0.4 12.66 0.4 12.66 1 11.26 1 11.26 0.4 0.4 0.4 0.4 108.4 11.26 108.4 11.26 107.8 12.66 107.8 12.66 108.4 15.09 108.4 15.09 107.04 16.19 107.04 16.19 108.4 16.93 108.4 16.93 107.04 18.03 107.04 18.03 108.4 25.98 108.4 25.98 107.8 27.38 107.8 27.38 108.4 33.49 108.4 33.49 107.04 34.59 107.04 34.59 108.4 35.33 108.4 35.33 107.04 36.43 107.04 36.43 108.4 37.17 108.4 37.17 107.04 38.27 107.04 38.27 108.4 39.01 108.4 39.01 107.04 40.11 107.04 40.11 108.4 40.7 108.4 40.7 107.8 42.1 107.8 42.1 108.4 53.73 108.4 53.73 107.04 54.83 107.04 54.83 108.4 55.42 108.4 55.42 107.8 56.82 107.8 56.82 108.4 57.41 108.4 57.41 107.04 58.51 107.04 58.51 108.4 59.25 108.4 59.25 107.04 60.35 107.04 60.35 108.4 61.09 108.4 61.09 107.04 62.19 107.04 62.19 108.4 62.93 108.4 62.93 107.04 64.03 107.04 64.03 108.4 ;
    LAYER met3 ;
      POLYGON 56.285 108.965 56.285 108.96 56.5 108.96 56.5 108.64 56.285 108.64 56.285 108.635 55.955 108.635 55.955 108.64 55.74 108.64 55.74 108.96 55.955 108.96 55.955 108.965 ;
      POLYGON 26.845 108.965 26.845 108.96 27.06 108.96 27.06 108.64 26.845 108.64 26.845 108.635 26.515 108.635 26.515 108.64 26.3 108.64 26.3 108.96 26.515 108.96 26.515 108.965 ;
      POLYGON 56.285 0.165 56.285 0.16 56.5 0.16 56.5 -0.16 56.285 -0.16 56.285 -0.165 55.955 -0.165 55.955 -0.16 55.74 -0.16 55.74 0.16 55.955 0.16 55.955 0.165 ;
      POLYGON 26.845 0.165 26.845 0.16 27.06 0.16 27.06 -0.16 26.845 -0.16 26.845 -0.165 26.515 -0.165 26.515 -0.16 26.3 -0.16 26.3 0.16 26.515 0.16 26.515 0.165 ;
      POLYGON 67.68 108.4 67.68 97.52 95.28 97.52 95.28 93.03 93.9 93.03 93.9 91.93 95.28 91.93 95.28 91.67 93.9 91.67 93.9 90.57 95.28 90.57 95.28 90.31 93.9 90.31 93.9 89.21 95.28 89.21 95.28 88.95 93.9 88.95 93.9 87.85 95.28 87.85 95.28 87.59 93.9 87.59 93.9 86.49 95.28 86.49 95.28 85.55 93.9 85.55 93.9 84.45 95.28 84.45 95.28 84.19 93.9 84.19 93.9 83.09 95.28 83.09 95.28 82.83 93.9 82.83 93.9 81.73 95.28 81.73 95.28 81.47 93.9 81.47 93.9 80.37 95.28 80.37 95.28 80.11 93.9 80.11 93.9 79.01 95.28 79.01 95.28 78.75 93.9 78.75 93.9 77.65 95.28 77.65 95.28 77.39 93.9 77.39 93.9 76.29 95.28 76.29 95.28 76.03 93.9 76.03 93.9 74.93 95.28 74.93 95.28 74.67 93.9 74.67 93.9 73.57 95.28 73.57 95.28 73.31 93.9 73.31 93.9 72.21 95.28 72.21 95.28 71.95 93.9 71.95 93.9 70.85 95.28 70.85 95.28 69.91 93.9 69.91 93.9 68.81 95.28 68.81 95.28 67.87 93.9 67.87 93.9 66.77 95.28 66.77 95.28 66.51 93.9 66.51 93.9 65.41 95.28 65.41 95.28 65.15 93.9 65.15 93.9 64.05 95.28 64.05 95.28 63.11 93.9 63.11 93.9 62.01 95.28 62.01 95.28 61.75 93.9 61.75 93.9 60.65 95.28 60.65 95.28 60.39 93.9 60.39 93.9 59.29 95.28 59.29 95.28 59.03 93.9 59.03 93.9 57.93 95.28 57.93 95.28 57.67 93.9 57.67 93.9 56.57 95.28 56.57 95.28 56.31 93.9 56.31 93.9 55.21 95.28 55.21 95.28 54.95 93.9 54.95 93.9 53.85 95.28 53.85 95.28 53.59 93.9 53.59 93.9 52.49 95.28 52.49 95.28 51.55 93.9 51.55 93.9 50.45 95.28 50.45 95.28 50.19 93.9 50.19 93.9 49.09 95.28 49.09 95.28 48.83 93.9 48.83 93.9 47.73 95.28 47.73 95.28 47.47 93.9 47.47 93.9 46.37 95.28 46.37 95.28 46.11 93.9 46.11 93.9 45.01 95.28 45.01 95.28 44.75 93.9 44.75 93.9 43.65 95.28 43.65 95.28 43.39 93.9 43.39 93.9 42.29 95.28 42.29 95.28 42.03 93.9 42.03 93.9 40.93 95.28 40.93 95.28 40.67 93.9 40.67 93.9 39.57 95.28 39.57 95.28 39.31 93.9 39.31 93.9 38.21 95.28 38.21 95.28 37.95 93.9 37.95 93.9 36.85 95.28 36.85 95.28 36.59 93.9 36.59 93.9 35.49 95.28 35.49 95.28 32.51 93.9 32.51 93.9 31.41 95.28 31.41 95.28 11.28 67.68 11.28 67.68 0.4 0.4 0.4 0.4 108.4 ;
    LAYER met5 ;
      POLYGON 66.48 107.2 66.48 96.32 94.08 96.32 94.08 88.2 90.88 88.2 90.88 81.8 94.08 81.8 94.08 67.8 90.88 67.8 90.88 61.4 94.08 61.4 94.08 47.4 90.88 47.4 90.88 41 94.08 41 94.08 27 90.88 27 90.88 20.6 94.08 20.6 94.08 12.48 66.48 12.48 66.48 1.6 1.6 1.6 1.6 20.6 4.8 20.6 4.8 27 1.6 27 1.6 41 4.8 41 4.8 47.4 1.6 47.4 1.6 61.4 4.8 61.4 4.8 67.8 1.6 67.8 1.6 81.8 4.8 81.8 4.8 88.2 1.6 88.2 1.6 107.2 ;
    LAYER met1 ;
      POLYGON 67.8 108.28 67.8 106.6 67.32 106.6 67.32 105.56 67.8 105.56 67.8 103.88 67.32 103.88 67.32 102.84 67.8 102.84 67.8 101.16 67.32 101.16 67.32 100.12 67.8 100.12 67.8 98.44 0.28 98.44 0.28 100.12 0.76 100.12 0.76 101.16 0.28 101.16 0.28 102.84 0.76 102.84 0.76 103.88 0.28 103.88 0.28 105.56 0.76 105.56 0.76 106.6 0.28 106.6 0.28 108.28 ;
      POLYGON 95.4 97.4 95.4 95.72 94.92 95.72 94.92 94.68 95.4 94.68 95.4 93 94.92 93 94.92 91.96 95.4 91.96 95.4 90.28 94.92 90.28 94.92 89.24 95.4 89.24 95.4 87.56 94.92 87.56 94.92 86.52 95.4 86.52 95.4 84.84 94.92 84.84 94.92 83.8 95.4 83.8 95.4 82.12 94.92 82.12 94.92 81.08 95.4 81.08 95.4 79.4 94.92 79.4 94.92 78.36 95.4 78.36 95.4 76.68 94.92 76.68 94.92 75.64 95.4 75.64 95.4 73.96 94.92 73.96 94.92 72.92 95.4 72.92 95.4 71.24 94.92 71.24 94.92 70.2 95.4 70.2 95.4 68.52 94.92 68.52 94.92 67.48 95.4 67.48 95.4 65.8 94.92 65.8 94.92 64.76 95.4 64.76 95.4 63.08 94.92 63.08 94.92 62.04 95.4 62.04 95.4 60.36 94.92 60.36 94.92 59.32 95.4 59.32 95.4 57.64 94.92 57.64 94.92 56.6 95.4 56.6 95.4 54.92 94.92 54.92 94.92 53.88 95.4 53.88 95.4 52.2 94.92 52.2 94.92 51.16 95.4 51.16 95.4 49.48 94.92 49.48 94.92 48.44 95.4 48.44 95.4 46.76 94.92 46.76 94.92 45.72 95.4 45.72 95.4 44.04 94.92 44.04 94.92 43 95.4 43 95.4 41.32 94.92 41.32 94.92 40.28 95.4 40.28 95.4 38.6 94.92 38.6 94.92 37.56 95.4 37.56 95.4 35.88 94.92 35.88 94.92 34.84 95.4 34.84 95.4 33.16 94.92 33.16 94.92 32.12 95.4 32.12 95.4 30.44 94.92 30.44 94.92 29.4 95.4 29.4 95.4 27.72 94.92 27.72 94.92 26.68 95.4 26.68 95.4 25 94.92 25 94.92 23.96 95.4 23.96 95.4 22.28 94.92 22.28 94.92 21.24 95.4 21.24 95.4 19.56 94.92 19.56 94.92 18.52 95.4 18.52 95.4 16.84 94.92 16.84 94.92 15.8 95.4 15.8 95.4 14.12 94.92 14.12 94.92 13.08 95.4 13.08 95.4 11.4 0.28 11.4 0.28 13.08 0.76 13.08 0.76 14.12 0.28 14.12 0.28 15.8 0.76 15.8 0.76 16.84 0.28 16.84 0.28 18.52 0.76 18.52 0.76 19.56 0.28 19.56 0.28 21.24 0.76 21.24 0.76 22.28 0.28 22.28 0.28 23.96 0.76 23.96 0.76 25 0.28 25 0.28 26.68 0.76 26.68 0.76 27.72 0.28 27.72 0.28 29.4 0.76 29.4 0.76 30.44 0.28 30.44 0.28 32.12 0.76 32.12 0.76 33.16 0.28 33.16 0.28 34.84 0.76 34.84 0.76 35.88 0.28 35.88 0.28 37.56 0.76 37.56 0.76 38.6 0.28 38.6 0.28 40.28 0.76 40.28 0.76 41.32 0.28 41.32 0.28 43 0.76 43 0.76 44.04 0.28 44.04 0.28 45.72 0.76 45.72 0.76 46.76 0.28 46.76 0.28 48.44 0.76 48.44 0.76 49.48 0.28 49.48 0.28 51.16 0.76 51.16 0.76 52.2 0.28 52.2 0.28 53.88 0.76 53.88 0.76 54.92 0.28 54.92 0.28 56.6 0.76 56.6 0.76 57.64 0.28 57.64 0.28 59.32 0.76 59.32 0.76 60.36 0.28 60.36 0.28 62.04 0.76 62.04 0.76 63.08 0.28 63.08 0.28 64.76 0.76 64.76 0.76 65.8 0.28 65.8 0.28 67.48 0.76 67.48 0.76 68.52 0.28 68.52 0.28 70.2 0.76 70.2 0.76 71.24 0.28 71.24 0.28 72.92 0.76 72.92 0.76 73.96 0.28 73.96 0.28 75.64 0.76 75.64 0.76 76.68 0.28 76.68 0.28 78.36 0.76 78.36 0.76 79.4 0.28 79.4 0.28 81.08 0.76 81.08 0.76 82.12 0.28 82.12 0.28 83.8 0.76 83.8 0.76 84.84 0.28 84.84 0.28 86.52 0.76 86.52 0.76 87.56 0.28 87.56 0.28 89.24 0.76 89.24 0.76 90.28 0.28 90.28 0.28 91.96 0.76 91.96 0.76 93 0.28 93 0.28 94.68 0.76 94.68 0.76 95.72 0.28 95.72 0.28 97.4 ;
      POLYGON 67.8 10.36 67.8 8.68 67.32 8.68 67.32 7.64 67.8 7.64 67.8 5.96 67.32 5.96 67.32 4.92 67.8 4.92 67.8 3.24 67.32 3.24 67.32 2.2 67.8 2.2 67.8 0.52 0.28 0.52 0.28 2.2 0.76 2.2 0.76 3.24 0.28 3.24 0.28 4.92 0.76 4.92 0.76 5.96 0.28 5.96 0.28 7.64 0.76 7.64 0.76 8.68 0.28 8.68 0.28 10.36 ;
    LAYER li1 ;
      POLYGON 67.91 108.63 67.91 97.75 95.51 97.75 95.51 11.05 67.91 11.05 67.91 0.17 0.17 0.17 0.17 108.63 ;
    LAYER mcon ;
      RECT 67.765 108.715 67.935 108.885 ;
      RECT 67.305 108.715 67.475 108.885 ;
      RECT 66.845 108.715 67.015 108.885 ;
      RECT 66.385 108.715 66.555 108.885 ;
      RECT 65.925 108.715 66.095 108.885 ;
      RECT 65.465 108.715 65.635 108.885 ;
      RECT 65.005 108.715 65.175 108.885 ;
      RECT 64.545 108.715 64.715 108.885 ;
      RECT 64.085 108.715 64.255 108.885 ;
      RECT 63.625 108.715 63.795 108.885 ;
      RECT 63.165 108.715 63.335 108.885 ;
      RECT 62.705 108.715 62.875 108.885 ;
      RECT 62.245 108.715 62.415 108.885 ;
      RECT 61.785 108.715 61.955 108.885 ;
      RECT 61.325 108.715 61.495 108.885 ;
      RECT 60.865 108.715 61.035 108.885 ;
      RECT 60.405 108.715 60.575 108.885 ;
      RECT 59.945 108.715 60.115 108.885 ;
      RECT 59.485 108.715 59.655 108.885 ;
      RECT 59.025 108.715 59.195 108.885 ;
      RECT 58.565 108.715 58.735 108.885 ;
      RECT 58.105 108.715 58.275 108.885 ;
      RECT 57.645 108.715 57.815 108.885 ;
      RECT 57.185 108.715 57.355 108.885 ;
      RECT 56.725 108.715 56.895 108.885 ;
      RECT 56.265 108.715 56.435 108.885 ;
      RECT 55.805 108.715 55.975 108.885 ;
      RECT 55.345 108.715 55.515 108.885 ;
      RECT 54.885 108.715 55.055 108.885 ;
      RECT 54.425 108.715 54.595 108.885 ;
      RECT 53.965 108.715 54.135 108.885 ;
      RECT 53.505 108.715 53.675 108.885 ;
      RECT 53.045 108.715 53.215 108.885 ;
      RECT 52.585 108.715 52.755 108.885 ;
      RECT 52.125 108.715 52.295 108.885 ;
      RECT 51.665 108.715 51.835 108.885 ;
      RECT 51.205 108.715 51.375 108.885 ;
      RECT 50.745 108.715 50.915 108.885 ;
      RECT 50.285 108.715 50.455 108.885 ;
      RECT 49.825 108.715 49.995 108.885 ;
      RECT 49.365 108.715 49.535 108.885 ;
      RECT 48.905 108.715 49.075 108.885 ;
      RECT 48.445 108.715 48.615 108.885 ;
      RECT 47.985 108.715 48.155 108.885 ;
      RECT 47.525 108.715 47.695 108.885 ;
      RECT 47.065 108.715 47.235 108.885 ;
      RECT 46.605 108.715 46.775 108.885 ;
      RECT 46.145 108.715 46.315 108.885 ;
      RECT 45.685 108.715 45.855 108.885 ;
      RECT 45.225 108.715 45.395 108.885 ;
      RECT 44.765 108.715 44.935 108.885 ;
      RECT 44.305 108.715 44.475 108.885 ;
      RECT 43.845 108.715 44.015 108.885 ;
      RECT 43.385 108.715 43.555 108.885 ;
      RECT 42.925 108.715 43.095 108.885 ;
      RECT 42.465 108.715 42.635 108.885 ;
      RECT 42.005 108.715 42.175 108.885 ;
      RECT 41.545 108.715 41.715 108.885 ;
      RECT 41.085 108.715 41.255 108.885 ;
      RECT 40.625 108.715 40.795 108.885 ;
      RECT 40.165 108.715 40.335 108.885 ;
      RECT 39.705 108.715 39.875 108.885 ;
      RECT 39.245 108.715 39.415 108.885 ;
      RECT 38.785 108.715 38.955 108.885 ;
      RECT 38.325 108.715 38.495 108.885 ;
      RECT 37.865 108.715 38.035 108.885 ;
      RECT 37.405 108.715 37.575 108.885 ;
      RECT 36.945 108.715 37.115 108.885 ;
      RECT 36.485 108.715 36.655 108.885 ;
      RECT 36.025 108.715 36.195 108.885 ;
      RECT 35.565 108.715 35.735 108.885 ;
      RECT 35.105 108.715 35.275 108.885 ;
      RECT 34.645 108.715 34.815 108.885 ;
      RECT 34.185 108.715 34.355 108.885 ;
      RECT 33.725 108.715 33.895 108.885 ;
      RECT 33.265 108.715 33.435 108.885 ;
      RECT 32.805 108.715 32.975 108.885 ;
      RECT 32.345 108.715 32.515 108.885 ;
      RECT 31.885 108.715 32.055 108.885 ;
      RECT 31.425 108.715 31.595 108.885 ;
      RECT 30.965 108.715 31.135 108.885 ;
      RECT 30.505 108.715 30.675 108.885 ;
      RECT 30.045 108.715 30.215 108.885 ;
      RECT 29.585 108.715 29.755 108.885 ;
      RECT 29.125 108.715 29.295 108.885 ;
      RECT 28.665 108.715 28.835 108.885 ;
      RECT 28.205 108.715 28.375 108.885 ;
      RECT 27.745 108.715 27.915 108.885 ;
      RECT 27.285 108.715 27.455 108.885 ;
      RECT 26.825 108.715 26.995 108.885 ;
      RECT 26.365 108.715 26.535 108.885 ;
      RECT 25.905 108.715 26.075 108.885 ;
      RECT 25.445 108.715 25.615 108.885 ;
      RECT 24.985 108.715 25.155 108.885 ;
      RECT 24.525 108.715 24.695 108.885 ;
      RECT 24.065 108.715 24.235 108.885 ;
      RECT 23.605 108.715 23.775 108.885 ;
      RECT 23.145 108.715 23.315 108.885 ;
      RECT 22.685 108.715 22.855 108.885 ;
      RECT 22.225 108.715 22.395 108.885 ;
      RECT 21.765 108.715 21.935 108.885 ;
      RECT 21.305 108.715 21.475 108.885 ;
      RECT 20.845 108.715 21.015 108.885 ;
      RECT 20.385 108.715 20.555 108.885 ;
      RECT 19.925 108.715 20.095 108.885 ;
      RECT 19.465 108.715 19.635 108.885 ;
      RECT 19.005 108.715 19.175 108.885 ;
      RECT 18.545 108.715 18.715 108.885 ;
      RECT 18.085 108.715 18.255 108.885 ;
      RECT 17.625 108.715 17.795 108.885 ;
      RECT 17.165 108.715 17.335 108.885 ;
      RECT 16.705 108.715 16.875 108.885 ;
      RECT 16.245 108.715 16.415 108.885 ;
      RECT 15.785 108.715 15.955 108.885 ;
      RECT 15.325 108.715 15.495 108.885 ;
      RECT 14.865 108.715 15.035 108.885 ;
      RECT 14.405 108.715 14.575 108.885 ;
      RECT 13.945 108.715 14.115 108.885 ;
      RECT 13.485 108.715 13.655 108.885 ;
      RECT 13.025 108.715 13.195 108.885 ;
      RECT 12.565 108.715 12.735 108.885 ;
      RECT 12.105 108.715 12.275 108.885 ;
      RECT 11.645 108.715 11.815 108.885 ;
      RECT 11.185 108.715 11.355 108.885 ;
      RECT 10.725 108.715 10.895 108.885 ;
      RECT 10.265 108.715 10.435 108.885 ;
      RECT 9.805 108.715 9.975 108.885 ;
      RECT 9.345 108.715 9.515 108.885 ;
      RECT 8.885 108.715 9.055 108.885 ;
      RECT 8.425 108.715 8.595 108.885 ;
      RECT 7.965 108.715 8.135 108.885 ;
      RECT 7.505 108.715 7.675 108.885 ;
      RECT 7.045 108.715 7.215 108.885 ;
      RECT 6.585 108.715 6.755 108.885 ;
      RECT 6.125 108.715 6.295 108.885 ;
      RECT 5.665 108.715 5.835 108.885 ;
      RECT 5.205 108.715 5.375 108.885 ;
      RECT 4.745 108.715 4.915 108.885 ;
      RECT 4.285 108.715 4.455 108.885 ;
      RECT 3.825 108.715 3.995 108.885 ;
      RECT 3.365 108.715 3.535 108.885 ;
      RECT 2.905 108.715 3.075 108.885 ;
      RECT 2.445 108.715 2.615 108.885 ;
      RECT 1.985 108.715 2.155 108.885 ;
      RECT 1.525 108.715 1.695 108.885 ;
      RECT 1.065 108.715 1.235 108.885 ;
      RECT 0.605 108.715 0.775 108.885 ;
      RECT 0.145 108.715 0.315 108.885 ;
      RECT 67.765 105.995 67.935 106.165 ;
      RECT 67.305 105.995 67.475 106.165 ;
      RECT 0.605 105.995 0.775 106.165 ;
      RECT 0.145 105.995 0.315 106.165 ;
      RECT 67.765 103.275 67.935 103.445 ;
      RECT 67.305 103.275 67.475 103.445 ;
      RECT 0.605 103.275 0.775 103.445 ;
      RECT 0.145 103.275 0.315 103.445 ;
      RECT 67.765 100.555 67.935 100.725 ;
      RECT 67.305 100.555 67.475 100.725 ;
      RECT 0.605 100.555 0.775 100.725 ;
      RECT 0.145 100.555 0.315 100.725 ;
      RECT 95.365 97.835 95.535 98.005 ;
      RECT 94.905 97.835 95.075 98.005 ;
      RECT 94.445 97.835 94.615 98.005 ;
      RECT 93.985 97.835 94.155 98.005 ;
      RECT 93.525 97.835 93.695 98.005 ;
      RECT 93.065 97.835 93.235 98.005 ;
      RECT 92.605 97.835 92.775 98.005 ;
      RECT 92.145 97.835 92.315 98.005 ;
      RECT 91.685 97.835 91.855 98.005 ;
      RECT 91.225 97.835 91.395 98.005 ;
      RECT 90.765 97.835 90.935 98.005 ;
      RECT 90.305 97.835 90.475 98.005 ;
      RECT 89.845 97.835 90.015 98.005 ;
      RECT 89.385 97.835 89.555 98.005 ;
      RECT 88.925 97.835 89.095 98.005 ;
      RECT 88.465 97.835 88.635 98.005 ;
      RECT 88.005 97.835 88.175 98.005 ;
      RECT 87.545 97.835 87.715 98.005 ;
      RECT 87.085 97.835 87.255 98.005 ;
      RECT 86.625 97.835 86.795 98.005 ;
      RECT 86.165 97.835 86.335 98.005 ;
      RECT 85.705 97.835 85.875 98.005 ;
      RECT 85.245 97.835 85.415 98.005 ;
      RECT 84.785 97.835 84.955 98.005 ;
      RECT 84.325 97.835 84.495 98.005 ;
      RECT 83.865 97.835 84.035 98.005 ;
      RECT 83.405 97.835 83.575 98.005 ;
      RECT 82.945 97.835 83.115 98.005 ;
      RECT 82.485 97.835 82.655 98.005 ;
      RECT 82.025 97.835 82.195 98.005 ;
      RECT 81.565 97.835 81.735 98.005 ;
      RECT 81.105 97.835 81.275 98.005 ;
      RECT 80.645 97.835 80.815 98.005 ;
      RECT 80.185 97.835 80.355 98.005 ;
      RECT 79.725 97.835 79.895 98.005 ;
      RECT 79.265 97.835 79.435 98.005 ;
      RECT 78.805 97.835 78.975 98.005 ;
      RECT 78.345 97.835 78.515 98.005 ;
      RECT 77.885 97.835 78.055 98.005 ;
      RECT 77.425 97.835 77.595 98.005 ;
      RECT 76.965 97.835 77.135 98.005 ;
      RECT 76.505 97.835 76.675 98.005 ;
      RECT 76.045 97.835 76.215 98.005 ;
      RECT 75.585 97.835 75.755 98.005 ;
      RECT 75.125 97.835 75.295 98.005 ;
      RECT 74.665 97.835 74.835 98.005 ;
      RECT 74.205 97.835 74.375 98.005 ;
      RECT 73.745 97.835 73.915 98.005 ;
      RECT 73.285 97.835 73.455 98.005 ;
      RECT 72.825 97.835 72.995 98.005 ;
      RECT 72.365 97.835 72.535 98.005 ;
      RECT 71.905 97.835 72.075 98.005 ;
      RECT 71.445 97.835 71.615 98.005 ;
      RECT 70.985 97.835 71.155 98.005 ;
      RECT 70.525 97.835 70.695 98.005 ;
      RECT 70.065 97.835 70.235 98.005 ;
      RECT 69.605 97.835 69.775 98.005 ;
      RECT 69.145 97.835 69.315 98.005 ;
      RECT 68.685 97.835 68.855 98.005 ;
      RECT 68.225 97.835 68.395 98.005 ;
      RECT 67.765 97.835 67.935 98.005 ;
      RECT 67.305 97.835 67.475 98.005 ;
      RECT 66.845 97.835 67.015 98.005 ;
      RECT 66.385 97.835 66.555 98.005 ;
      RECT 65.925 97.835 66.095 98.005 ;
      RECT 65.465 97.835 65.635 98.005 ;
      RECT 65.005 97.835 65.175 98.005 ;
      RECT 64.545 97.835 64.715 98.005 ;
      RECT 64.085 97.835 64.255 98.005 ;
      RECT 63.625 97.835 63.795 98.005 ;
      RECT 63.165 97.835 63.335 98.005 ;
      RECT 62.705 97.835 62.875 98.005 ;
      RECT 62.245 97.835 62.415 98.005 ;
      RECT 61.785 97.835 61.955 98.005 ;
      RECT 61.325 97.835 61.495 98.005 ;
      RECT 60.865 97.835 61.035 98.005 ;
      RECT 60.405 97.835 60.575 98.005 ;
      RECT 59.945 97.835 60.115 98.005 ;
      RECT 59.485 97.835 59.655 98.005 ;
      RECT 59.025 97.835 59.195 98.005 ;
      RECT 58.565 97.835 58.735 98.005 ;
      RECT 58.105 97.835 58.275 98.005 ;
      RECT 57.645 97.835 57.815 98.005 ;
      RECT 57.185 97.835 57.355 98.005 ;
      RECT 56.725 97.835 56.895 98.005 ;
      RECT 56.265 97.835 56.435 98.005 ;
      RECT 55.805 97.835 55.975 98.005 ;
      RECT 55.345 97.835 55.515 98.005 ;
      RECT 54.885 97.835 55.055 98.005 ;
      RECT 54.425 97.835 54.595 98.005 ;
      RECT 53.965 97.835 54.135 98.005 ;
      RECT 53.505 97.835 53.675 98.005 ;
      RECT 53.045 97.835 53.215 98.005 ;
      RECT 52.585 97.835 52.755 98.005 ;
      RECT 52.125 97.835 52.295 98.005 ;
      RECT 51.665 97.835 51.835 98.005 ;
      RECT 51.205 97.835 51.375 98.005 ;
      RECT 50.745 97.835 50.915 98.005 ;
      RECT 50.285 97.835 50.455 98.005 ;
      RECT 49.825 97.835 49.995 98.005 ;
      RECT 49.365 97.835 49.535 98.005 ;
      RECT 48.905 97.835 49.075 98.005 ;
      RECT 48.445 97.835 48.615 98.005 ;
      RECT 47.985 97.835 48.155 98.005 ;
      RECT 47.525 97.835 47.695 98.005 ;
      RECT 47.065 97.835 47.235 98.005 ;
      RECT 46.605 97.835 46.775 98.005 ;
      RECT 46.145 97.835 46.315 98.005 ;
      RECT 45.685 97.835 45.855 98.005 ;
      RECT 45.225 97.835 45.395 98.005 ;
      RECT 44.765 97.835 44.935 98.005 ;
      RECT 44.305 97.835 44.475 98.005 ;
      RECT 43.845 97.835 44.015 98.005 ;
      RECT 43.385 97.835 43.555 98.005 ;
      RECT 42.925 97.835 43.095 98.005 ;
      RECT 42.465 97.835 42.635 98.005 ;
      RECT 42.005 97.835 42.175 98.005 ;
      RECT 41.545 97.835 41.715 98.005 ;
      RECT 41.085 97.835 41.255 98.005 ;
      RECT 40.625 97.835 40.795 98.005 ;
      RECT 40.165 97.835 40.335 98.005 ;
      RECT 39.705 97.835 39.875 98.005 ;
      RECT 39.245 97.835 39.415 98.005 ;
      RECT 38.785 97.835 38.955 98.005 ;
      RECT 38.325 97.835 38.495 98.005 ;
      RECT 37.865 97.835 38.035 98.005 ;
      RECT 37.405 97.835 37.575 98.005 ;
      RECT 36.945 97.835 37.115 98.005 ;
      RECT 36.485 97.835 36.655 98.005 ;
      RECT 36.025 97.835 36.195 98.005 ;
      RECT 35.565 97.835 35.735 98.005 ;
      RECT 35.105 97.835 35.275 98.005 ;
      RECT 34.645 97.835 34.815 98.005 ;
      RECT 34.185 97.835 34.355 98.005 ;
      RECT 33.725 97.835 33.895 98.005 ;
      RECT 33.265 97.835 33.435 98.005 ;
      RECT 32.805 97.835 32.975 98.005 ;
      RECT 32.345 97.835 32.515 98.005 ;
      RECT 31.885 97.835 32.055 98.005 ;
      RECT 31.425 97.835 31.595 98.005 ;
      RECT 30.965 97.835 31.135 98.005 ;
      RECT 30.505 97.835 30.675 98.005 ;
      RECT 30.045 97.835 30.215 98.005 ;
      RECT 29.585 97.835 29.755 98.005 ;
      RECT 29.125 97.835 29.295 98.005 ;
      RECT 28.665 97.835 28.835 98.005 ;
      RECT 28.205 97.835 28.375 98.005 ;
      RECT 27.745 97.835 27.915 98.005 ;
      RECT 27.285 97.835 27.455 98.005 ;
      RECT 26.825 97.835 26.995 98.005 ;
      RECT 26.365 97.835 26.535 98.005 ;
      RECT 25.905 97.835 26.075 98.005 ;
      RECT 25.445 97.835 25.615 98.005 ;
      RECT 24.985 97.835 25.155 98.005 ;
      RECT 24.525 97.835 24.695 98.005 ;
      RECT 24.065 97.835 24.235 98.005 ;
      RECT 23.605 97.835 23.775 98.005 ;
      RECT 23.145 97.835 23.315 98.005 ;
      RECT 22.685 97.835 22.855 98.005 ;
      RECT 22.225 97.835 22.395 98.005 ;
      RECT 21.765 97.835 21.935 98.005 ;
      RECT 21.305 97.835 21.475 98.005 ;
      RECT 20.845 97.835 21.015 98.005 ;
      RECT 20.385 97.835 20.555 98.005 ;
      RECT 19.925 97.835 20.095 98.005 ;
      RECT 19.465 97.835 19.635 98.005 ;
      RECT 19.005 97.835 19.175 98.005 ;
      RECT 18.545 97.835 18.715 98.005 ;
      RECT 18.085 97.835 18.255 98.005 ;
      RECT 17.625 97.835 17.795 98.005 ;
      RECT 17.165 97.835 17.335 98.005 ;
      RECT 16.705 97.835 16.875 98.005 ;
      RECT 16.245 97.835 16.415 98.005 ;
      RECT 15.785 97.835 15.955 98.005 ;
      RECT 15.325 97.835 15.495 98.005 ;
      RECT 14.865 97.835 15.035 98.005 ;
      RECT 14.405 97.835 14.575 98.005 ;
      RECT 13.945 97.835 14.115 98.005 ;
      RECT 13.485 97.835 13.655 98.005 ;
      RECT 13.025 97.835 13.195 98.005 ;
      RECT 12.565 97.835 12.735 98.005 ;
      RECT 12.105 97.835 12.275 98.005 ;
      RECT 11.645 97.835 11.815 98.005 ;
      RECT 11.185 97.835 11.355 98.005 ;
      RECT 10.725 97.835 10.895 98.005 ;
      RECT 10.265 97.835 10.435 98.005 ;
      RECT 9.805 97.835 9.975 98.005 ;
      RECT 9.345 97.835 9.515 98.005 ;
      RECT 8.885 97.835 9.055 98.005 ;
      RECT 8.425 97.835 8.595 98.005 ;
      RECT 7.965 97.835 8.135 98.005 ;
      RECT 7.505 97.835 7.675 98.005 ;
      RECT 7.045 97.835 7.215 98.005 ;
      RECT 6.585 97.835 6.755 98.005 ;
      RECT 6.125 97.835 6.295 98.005 ;
      RECT 5.665 97.835 5.835 98.005 ;
      RECT 5.205 97.835 5.375 98.005 ;
      RECT 4.745 97.835 4.915 98.005 ;
      RECT 4.285 97.835 4.455 98.005 ;
      RECT 3.825 97.835 3.995 98.005 ;
      RECT 3.365 97.835 3.535 98.005 ;
      RECT 2.905 97.835 3.075 98.005 ;
      RECT 2.445 97.835 2.615 98.005 ;
      RECT 1.985 97.835 2.155 98.005 ;
      RECT 1.525 97.835 1.695 98.005 ;
      RECT 1.065 97.835 1.235 98.005 ;
      RECT 0.605 97.835 0.775 98.005 ;
      RECT 0.145 97.835 0.315 98.005 ;
      RECT 95.365 95.115 95.535 95.285 ;
      RECT 94.905 95.115 95.075 95.285 ;
      RECT 0.605 95.115 0.775 95.285 ;
      RECT 0.145 95.115 0.315 95.285 ;
      RECT 95.365 92.395 95.535 92.565 ;
      RECT 94.905 92.395 95.075 92.565 ;
      RECT 0.605 92.395 0.775 92.565 ;
      RECT 0.145 92.395 0.315 92.565 ;
      RECT 95.365 89.675 95.535 89.845 ;
      RECT 94.905 89.675 95.075 89.845 ;
      RECT 0.605 89.675 0.775 89.845 ;
      RECT 0.145 89.675 0.315 89.845 ;
      RECT 95.365 86.955 95.535 87.125 ;
      RECT 94.905 86.955 95.075 87.125 ;
      RECT 0.605 86.955 0.775 87.125 ;
      RECT 0.145 86.955 0.315 87.125 ;
      RECT 95.365 84.235 95.535 84.405 ;
      RECT 94.905 84.235 95.075 84.405 ;
      RECT 0.605 84.235 0.775 84.405 ;
      RECT 0.145 84.235 0.315 84.405 ;
      RECT 95.365 81.515 95.535 81.685 ;
      RECT 94.905 81.515 95.075 81.685 ;
      RECT 0.605 81.515 0.775 81.685 ;
      RECT 0.145 81.515 0.315 81.685 ;
      RECT 95.365 78.795 95.535 78.965 ;
      RECT 94.905 78.795 95.075 78.965 ;
      RECT 0.605 78.795 0.775 78.965 ;
      RECT 0.145 78.795 0.315 78.965 ;
      RECT 95.365 76.075 95.535 76.245 ;
      RECT 94.905 76.075 95.075 76.245 ;
      RECT 0.605 76.075 0.775 76.245 ;
      RECT 0.145 76.075 0.315 76.245 ;
      RECT 95.365 73.355 95.535 73.525 ;
      RECT 94.905 73.355 95.075 73.525 ;
      RECT 0.605 73.355 0.775 73.525 ;
      RECT 0.145 73.355 0.315 73.525 ;
      RECT 95.365 70.635 95.535 70.805 ;
      RECT 94.905 70.635 95.075 70.805 ;
      RECT 0.605 70.635 0.775 70.805 ;
      RECT 0.145 70.635 0.315 70.805 ;
      RECT 95.365 67.915 95.535 68.085 ;
      RECT 94.905 67.915 95.075 68.085 ;
      RECT 0.605 67.915 0.775 68.085 ;
      RECT 0.145 67.915 0.315 68.085 ;
      RECT 95.365 65.195 95.535 65.365 ;
      RECT 94.905 65.195 95.075 65.365 ;
      RECT 0.605 65.195 0.775 65.365 ;
      RECT 0.145 65.195 0.315 65.365 ;
      RECT 95.365 62.475 95.535 62.645 ;
      RECT 94.905 62.475 95.075 62.645 ;
      RECT 0.605 62.475 0.775 62.645 ;
      RECT 0.145 62.475 0.315 62.645 ;
      RECT 95.365 59.755 95.535 59.925 ;
      RECT 94.905 59.755 95.075 59.925 ;
      RECT 0.605 59.755 0.775 59.925 ;
      RECT 0.145 59.755 0.315 59.925 ;
      RECT 95.365 57.035 95.535 57.205 ;
      RECT 94.905 57.035 95.075 57.205 ;
      RECT 0.605 57.035 0.775 57.205 ;
      RECT 0.145 57.035 0.315 57.205 ;
      RECT 95.365 54.315 95.535 54.485 ;
      RECT 94.905 54.315 95.075 54.485 ;
      RECT 0.605 54.315 0.775 54.485 ;
      RECT 0.145 54.315 0.315 54.485 ;
      RECT 95.365 51.595 95.535 51.765 ;
      RECT 94.905 51.595 95.075 51.765 ;
      RECT 0.605 51.595 0.775 51.765 ;
      RECT 0.145 51.595 0.315 51.765 ;
      RECT 95.365 48.875 95.535 49.045 ;
      RECT 94.905 48.875 95.075 49.045 ;
      RECT 0.605 48.875 0.775 49.045 ;
      RECT 0.145 48.875 0.315 49.045 ;
      RECT 95.365 46.155 95.535 46.325 ;
      RECT 94.905 46.155 95.075 46.325 ;
      RECT 0.605 46.155 0.775 46.325 ;
      RECT 0.145 46.155 0.315 46.325 ;
      RECT 95.365 43.435 95.535 43.605 ;
      RECT 94.905 43.435 95.075 43.605 ;
      RECT 0.605 43.435 0.775 43.605 ;
      RECT 0.145 43.435 0.315 43.605 ;
      RECT 95.365 40.715 95.535 40.885 ;
      RECT 94.905 40.715 95.075 40.885 ;
      RECT 0.605 40.715 0.775 40.885 ;
      RECT 0.145 40.715 0.315 40.885 ;
      RECT 95.365 37.995 95.535 38.165 ;
      RECT 94.905 37.995 95.075 38.165 ;
      RECT 0.605 37.995 0.775 38.165 ;
      RECT 0.145 37.995 0.315 38.165 ;
      RECT 95.365 35.275 95.535 35.445 ;
      RECT 94.905 35.275 95.075 35.445 ;
      RECT 0.605 35.275 0.775 35.445 ;
      RECT 0.145 35.275 0.315 35.445 ;
      RECT 95.365 32.555 95.535 32.725 ;
      RECT 94.905 32.555 95.075 32.725 ;
      RECT 0.605 32.555 0.775 32.725 ;
      RECT 0.145 32.555 0.315 32.725 ;
      RECT 95.365 29.835 95.535 30.005 ;
      RECT 94.905 29.835 95.075 30.005 ;
      RECT 0.605 29.835 0.775 30.005 ;
      RECT 0.145 29.835 0.315 30.005 ;
      RECT 95.365 27.115 95.535 27.285 ;
      RECT 94.905 27.115 95.075 27.285 ;
      RECT 0.605 27.115 0.775 27.285 ;
      RECT 0.145 27.115 0.315 27.285 ;
      RECT 95.365 24.395 95.535 24.565 ;
      RECT 94.905 24.395 95.075 24.565 ;
      RECT 0.605 24.395 0.775 24.565 ;
      RECT 0.145 24.395 0.315 24.565 ;
      RECT 95.365 21.675 95.535 21.845 ;
      RECT 94.905 21.675 95.075 21.845 ;
      RECT 0.605 21.675 0.775 21.845 ;
      RECT 0.145 21.675 0.315 21.845 ;
      RECT 95.365 18.955 95.535 19.125 ;
      RECT 94.905 18.955 95.075 19.125 ;
      RECT 0.605 18.955 0.775 19.125 ;
      RECT 0.145 18.955 0.315 19.125 ;
      RECT 95.365 16.235 95.535 16.405 ;
      RECT 94.905 16.235 95.075 16.405 ;
      RECT 0.605 16.235 0.775 16.405 ;
      RECT 0.145 16.235 0.315 16.405 ;
      RECT 95.365 13.515 95.535 13.685 ;
      RECT 94.905 13.515 95.075 13.685 ;
      RECT 0.605 13.515 0.775 13.685 ;
      RECT 0.145 13.515 0.315 13.685 ;
      RECT 95.365 10.795 95.535 10.965 ;
      RECT 94.905 10.795 95.075 10.965 ;
      RECT 94.445 10.795 94.615 10.965 ;
      RECT 93.985 10.795 94.155 10.965 ;
      RECT 93.525 10.795 93.695 10.965 ;
      RECT 93.065 10.795 93.235 10.965 ;
      RECT 92.605 10.795 92.775 10.965 ;
      RECT 92.145 10.795 92.315 10.965 ;
      RECT 91.685 10.795 91.855 10.965 ;
      RECT 91.225 10.795 91.395 10.965 ;
      RECT 90.765 10.795 90.935 10.965 ;
      RECT 90.305 10.795 90.475 10.965 ;
      RECT 89.845 10.795 90.015 10.965 ;
      RECT 89.385 10.795 89.555 10.965 ;
      RECT 88.925 10.795 89.095 10.965 ;
      RECT 88.465 10.795 88.635 10.965 ;
      RECT 88.005 10.795 88.175 10.965 ;
      RECT 87.545 10.795 87.715 10.965 ;
      RECT 87.085 10.795 87.255 10.965 ;
      RECT 86.625 10.795 86.795 10.965 ;
      RECT 86.165 10.795 86.335 10.965 ;
      RECT 85.705 10.795 85.875 10.965 ;
      RECT 85.245 10.795 85.415 10.965 ;
      RECT 84.785 10.795 84.955 10.965 ;
      RECT 84.325 10.795 84.495 10.965 ;
      RECT 83.865 10.795 84.035 10.965 ;
      RECT 83.405 10.795 83.575 10.965 ;
      RECT 82.945 10.795 83.115 10.965 ;
      RECT 82.485 10.795 82.655 10.965 ;
      RECT 82.025 10.795 82.195 10.965 ;
      RECT 81.565 10.795 81.735 10.965 ;
      RECT 81.105 10.795 81.275 10.965 ;
      RECT 80.645 10.795 80.815 10.965 ;
      RECT 80.185 10.795 80.355 10.965 ;
      RECT 79.725 10.795 79.895 10.965 ;
      RECT 79.265 10.795 79.435 10.965 ;
      RECT 78.805 10.795 78.975 10.965 ;
      RECT 78.345 10.795 78.515 10.965 ;
      RECT 77.885 10.795 78.055 10.965 ;
      RECT 77.425 10.795 77.595 10.965 ;
      RECT 76.965 10.795 77.135 10.965 ;
      RECT 76.505 10.795 76.675 10.965 ;
      RECT 76.045 10.795 76.215 10.965 ;
      RECT 75.585 10.795 75.755 10.965 ;
      RECT 75.125 10.795 75.295 10.965 ;
      RECT 74.665 10.795 74.835 10.965 ;
      RECT 74.205 10.795 74.375 10.965 ;
      RECT 73.745 10.795 73.915 10.965 ;
      RECT 73.285 10.795 73.455 10.965 ;
      RECT 72.825 10.795 72.995 10.965 ;
      RECT 72.365 10.795 72.535 10.965 ;
      RECT 71.905 10.795 72.075 10.965 ;
      RECT 71.445 10.795 71.615 10.965 ;
      RECT 70.985 10.795 71.155 10.965 ;
      RECT 70.525 10.795 70.695 10.965 ;
      RECT 70.065 10.795 70.235 10.965 ;
      RECT 69.605 10.795 69.775 10.965 ;
      RECT 69.145 10.795 69.315 10.965 ;
      RECT 68.685 10.795 68.855 10.965 ;
      RECT 68.225 10.795 68.395 10.965 ;
      RECT 67.765 10.795 67.935 10.965 ;
      RECT 67.305 10.795 67.475 10.965 ;
      RECT 66.845 10.795 67.015 10.965 ;
      RECT 66.385 10.795 66.555 10.965 ;
      RECT 65.925 10.795 66.095 10.965 ;
      RECT 65.465 10.795 65.635 10.965 ;
      RECT 65.005 10.795 65.175 10.965 ;
      RECT 64.545 10.795 64.715 10.965 ;
      RECT 64.085 10.795 64.255 10.965 ;
      RECT 63.625 10.795 63.795 10.965 ;
      RECT 63.165 10.795 63.335 10.965 ;
      RECT 62.705 10.795 62.875 10.965 ;
      RECT 62.245 10.795 62.415 10.965 ;
      RECT 61.785 10.795 61.955 10.965 ;
      RECT 61.325 10.795 61.495 10.965 ;
      RECT 60.865 10.795 61.035 10.965 ;
      RECT 60.405 10.795 60.575 10.965 ;
      RECT 59.945 10.795 60.115 10.965 ;
      RECT 59.485 10.795 59.655 10.965 ;
      RECT 59.025 10.795 59.195 10.965 ;
      RECT 58.565 10.795 58.735 10.965 ;
      RECT 58.105 10.795 58.275 10.965 ;
      RECT 57.645 10.795 57.815 10.965 ;
      RECT 57.185 10.795 57.355 10.965 ;
      RECT 56.725 10.795 56.895 10.965 ;
      RECT 56.265 10.795 56.435 10.965 ;
      RECT 55.805 10.795 55.975 10.965 ;
      RECT 55.345 10.795 55.515 10.965 ;
      RECT 54.885 10.795 55.055 10.965 ;
      RECT 54.425 10.795 54.595 10.965 ;
      RECT 53.965 10.795 54.135 10.965 ;
      RECT 53.505 10.795 53.675 10.965 ;
      RECT 53.045 10.795 53.215 10.965 ;
      RECT 52.585 10.795 52.755 10.965 ;
      RECT 52.125 10.795 52.295 10.965 ;
      RECT 51.665 10.795 51.835 10.965 ;
      RECT 51.205 10.795 51.375 10.965 ;
      RECT 50.745 10.795 50.915 10.965 ;
      RECT 50.285 10.795 50.455 10.965 ;
      RECT 49.825 10.795 49.995 10.965 ;
      RECT 49.365 10.795 49.535 10.965 ;
      RECT 48.905 10.795 49.075 10.965 ;
      RECT 48.445 10.795 48.615 10.965 ;
      RECT 47.985 10.795 48.155 10.965 ;
      RECT 47.525 10.795 47.695 10.965 ;
      RECT 47.065 10.795 47.235 10.965 ;
      RECT 46.605 10.795 46.775 10.965 ;
      RECT 46.145 10.795 46.315 10.965 ;
      RECT 45.685 10.795 45.855 10.965 ;
      RECT 45.225 10.795 45.395 10.965 ;
      RECT 44.765 10.795 44.935 10.965 ;
      RECT 44.305 10.795 44.475 10.965 ;
      RECT 43.845 10.795 44.015 10.965 ;
      RECT 43.385 10.795 43.555 10.965 ;
      RECT 42.925 10.795 43.095 10.965 ;
      RECT 42.465 10.795 42.635 10.965 ;
      RECT 42.005 10.795 42.175 10.965 ;
      RECT 41.545 10.795 41.715 10.965 ;
      RECT 41.085 10.795 41.255 10.965 ;
      RECT 40.625 10.795 40.795 10.965 ;
      RECT 40.165 10.795 40.335 10.965 ;
      RECT 39.705 10.795 39.875 10.965 ;
      RECT 39.245 10.795 39.415 10.965 ;
      RECT 38.785 10.795 38.955 10.965 ;
      RECT 38.325 10.795 38.495 10.965 ;
      RECT 37.865 10.795 38.035 10.965 ;
      RECT 37.405 10.795 37.575 10.965 ;
      RECT 36.945 10.795 37.115 10.965 ;
      RECT 36.485 10.795 36.655 10.965 ;
      RECT 36.025 10.795 36.195 10.965 ;
      RECT 35.565 10.795 35.735 10.965 ;
      RECT 35.105 10.795 35.275 10.965 ;
      RECT 34.645 10.795 34.815 10.965 ;
      RECT 34.185 10.795 34.355 10.965 ;
      RECT 33.725 10.795 33.895 10.965 ;
      RECT 33.265 10.795 33.435 10.965 ;
      RECT 32.805 10.795 32.975 10.965 ;
      RECT 32.345 10.795 32.515 10.965 ;
      RECT 31.885 10.795 32.055 10.965 ;
      RECT 31.425 10.795 31.595 10.965 ;
      RECT 30.965 10.795 31.135 10.965 ;
      RECT 30.505 10.795 30.675 10.965 ;
      RECT 30.045 10.795 30.215 10.965 ;
      RECT 29.585 10.795 29.755 10.965 ;
      RECT 29.125 10.795 29.295 10.965 ;
      RECT 28.665 10.795 28.835 10.965 ;
      RECT 28.205 10.795 28.375 10.965 ;
      RECT 27.745 10.795 27.915 10.965 ;
      RECT 27.285 10.795 27.455 10.965 ;
      RECT 26.825 10.795 26.995 10.965 ;
      RECT 26.365 10.795 26.535 10.965 ;
      RECT 25.905 10.795 26.075 10.965 ;
      RECT 25.445 10.795 25.615 10.965 ;
      RECT 24.985 10.795 25.155 10.965 ;
      RECT 24.525 10.795 24.695 10.965 ;
      RECT 24.065 10.795 24.235 10.965 ;
      RECT 23.605 10.795 23.775 10.965 ;
      RECT 23.145 10.795 23.315 10.965 ;
      RECT 22.685 10.795 22.855 10.965 ;
      RECT 22.225 10.795 22.395 10.965 ;
      RECT 21.765 10.795 21.935 10.965 ;
      RECT 21.305 10.795 21.475 10.965 ;
      RECT 20.845 10.795 21.015 10.965 ;
      RECT 20.385 10.795 20.555 10.965 ;
      RECT 19.925 10.795 20.095 10.965 ;
      RECT 19.465 10.795 19.635 10.965 ;
      RECT 19.005 10.795 19.175 10.965 ;
      RECT 18.545 10.795 18.715 10.965 ;
      RECT 18.085 10.795 18.255 10.965 ;
      RECT 17.625 10.795 17.795 10.965 ;
      RECT 17.165 10.795 17.335 10.965 ;
      RECT 16.705 10.795 16.875 10.965 ;
      RECT 16.245 10.795 16.415 10.965 ;
      RECT 15.785 10.795 15.955 10.965 ;
      RECT 15.325 10.795 15.495 10.965 ;
      RECT 14.865 10.795 15.035 10.965 ;
      RECT 14.405 10.795 14.575 10.965 ;
      RECT 13.945 10.795 14.115 10.965 ;
      RECT 13.485 10.795 13.655 10.965 ;
      RECT 13.025 10.795 13.195 10.965 ;
      RECT 12.565 10.795 12.735 10.965 ;
      RECT 12.105 10.795 12.275 10.965 ;
      RECT 11.645 10.795 11.815 10.965 ;
      RECT 11.185 10.795 11.355 10.965 ;
      RECT 10.725 10.795 10.895 10.965 ;
      RECT 10.265 10.795 10.435 10.965 ;
      RECT 9.805 10.795 9.975 10.965 ;
      RECT 9.345 10.795 9.515 10.965 ;
      RECT 8.885 10.795 9.055 10.965 ;
      RECT 8.425 10.795 8.595 10.965 ;
      RECT 7.965 10.795 8.135 10.965 ;
      RECT 7.505 10.795 7.675 10.965 ;
      RECT 7.045 10.795 7.215 10.965 ;
      RECT 6.585 10.795 6.755 10.965 ;
      RECT 6.125 10.795 6.295 10.965 ;
      RECT 5.665 10.795 5.835 10.965 ;
      RECT 5.205 10.795 5.375 10.965 ;
      RECT 4.745 10.795 4.915 10.965 ;
      RECT 4.285 10.795 4.455 10.965 ;
      RECT 3.825 10.795 3.995 10.965 ;
      RECT 3.365 10.795 3.535 10.965 ;
      RECT 2.905 10.795 3.075 10.965 ;
      RECT 2.445 10.795 2.615 10.965 ;
      RECT 1.985 10.795 2.155 10.965 ;
      RECT 1.525 10.795 1.695 10.965 ;
      RECT 1.065 10.795 1.235 10.965 ;
      RECT 0.605 10.795 0.775 10.965 ;
      RECT 0.145 10.795 0.315 10.965 ;
      RECT 67.765 8.075 67.935 8.245 ;
      RECT 67.305 8.075 67.475 8.245 ;
      RECT 0.605 8.075 0.775 8.245 ;
      RECT 0.145 8.075 0.315 8.245 ;
      RECT 67.765 5.355 67.935 5.525 ;
      RECT 67.305 5.355 67.475 5.525 ;
      RECT 0.605 5.355 0.775 5.525 ;
      RECT 0.145 5.355 0.315 5.525 ;
      RECT 67.765 2.635 67.935 2.805 ;
      RECT 67.305 2.635 67.475 2.805 ;
      RECT 0.605 2.635 0.775 2.805 ;
      RECT 0.145 2.635 0.315 2.805 ;
      RECT 67.765 -0.085 67.935 0.085 ;
      RECT 67.305 -0.085 67.475 0.085 ;
      RECT 66.845 -0.085 67.015 0.085 ;
      RECT 66.385 -0.085 66.555 0.085 ;
      RECT 65.925 -0.085 66.095 0.085 ;
      RECT 65.465 -0.085 65.635 0.085 ;
      RECT 65.005 -0.085 65.175 0.085 ;
      RECT 64.545 -0.085 64.715 0.085 ;
      RECT 64.085 -0.085 64.255 0.085 ;
      RECT 63.625 -0.085 63.795 0.085 ;
      RECT 63.165 -0.085 63.335 0.085 ;
      RECT 62.705 -0.085 62.875 0.085 ;
      RECT 62.245 -0.085 62.415 0.085 ;
      RECT 61.785 -0.085 61.955 0.085 ;
      RECT 61.325 -0.085 61.495 0.085 ;
      RECT 60.865 -0.085 61.035 0.085 ;
      RECT 60.405 -0.085 60.575 0.085 ;
      RECT 59.945 -0.085 60.115 0.085 ;
      RECT 59.485 -0.085 59.655 0.085 ;
      RECT 59.025 -0.085 59.195 0.085 ;
      RECT 58.565 -0.085 58.735 0.085 ;
      RECT 58.105 -0.085 58.275 0.085 ;
      RECT 57.645 -0.085 57.815 0.085 ;
      RECT 57.185 -0.085 57.355 0.085 ;
      RECT 56.725 -0.085 56.895 0.085 ;
      RECT 56.265 -0.085 56.435 0.085 ;
      RECT 55.805 -0.085 55.975 0.085 ;
      RECT 55.345 -0.085 55.515 0.085 ;
      RECT 54.885 -0.085 55.055 0.085 ;
      RECT 54.425 -0.085 54.595 0.085 ;
      RECT 53.965 -0.085 54.135 0.085 ;
      RECT 53.505 -0.085 53.675 0.085 ;
      RECT 53.045 -0.085 53.215 0.085 ;
      RECT 52.585 -0.085 52.755 0.085 ;
      RECT 52.125 -0.085 52.295 0.085 ;
      RECT 51.665 -0.085 51.835 0.085 ;
      RECT 51.205 -0.085 51.375 0.085 ;
      RECT 50.745 -0.085 50.915 0.085 ;
      RECT 50.285 -0.085 50.455 0.085 ;
      RECT 49.825 -0.085 49.995 0.085 ;
      RECT 49.365 -0.085 49.535 0.085 ;
      RECT 48.905 -0.085 49.075 0.085 ;
      RECT 48.445 -0.085 48.615 0.085 ;
      RECT 47.985 -0.085 48.155 0.085 ;
      RECT 47.525 -0.085 47.695 0.085 ;
      RECT 47.065 -0.085 47.235 0.085 ;
      RECT 46.605 -0.085 46.775 0.085 ;
      RECT 46.145 -0.085 46.315 0.085 ;
      RECT 45.685 -0.085 45.855 0.085 ;
      RECT 45.225 -0.085 45.395 0.085 ;
      RECT 44.765 -0.085 44.935 0.085 ;
      RECT 44.305 -0.085 44.475 0.085 ;
      RECT 43.845 -0.085 44.015 0.085 ;
      RECT 43.385 -0.085 43.555 0.085 ;
      RECT 42.925 -0.085 43.095 0.085 ;
      RECT 42.465 -0.085 42.635 0.085 ;
      RECT 42.005 -0.085 42.175 0.085 ;
      RECT 41.545 -0.085 41.715 0.085 ;
      RECT 41.085 -0.085 41.255 0.085 ;
      RECT 40.625 -0.085 40.795 0.085 ;
      RECT 40.165 -0.085 40.335 0.085 ;
      RECT 39.705 -0.085 39.875 0.085 ;
      RECT 39.245 -0.085 39.415 0.085 ;
      RECT 38.785 -0.085 38.955 0.085 ;
      RECT 38.325 -0.085 38.495 0.085 ;
      RECT 37.865 -0.085 38.035 0.085 ;
      RECT 37.405 -0.085 37.575 0.085 ;
      RECT 36.945 -0.085 37.115 0.085 ;
      RECT 36.485 -0.085 36.655 0.085 ;
      RECT 36.025 -0.085 36.195 0.085 ;
      RECT 35.565 -0.085 35.735 0.085 ;
      RECT 35.105 -0.085 35.275 0.085 ;
      RECT 34.645 -0.085 34.815 0.085 ;
      RECT 34.185 -0.085 34.355 0.085 ;
      RECT 33.725 -0.085 33.895 0.085 ;
      RECT 33.265 -0.085 33.435 0.085 ;
      RECT 32.805 -0.085 32.975 0.085 ;
      RECT 32.345 -0.085 32.515 0.085 ;
      RECT 31.885 -0.085 32.055 0.085 ;
      RECT 31.425 -0.085 31.595 0.085 ;
      RECT 30.965 -0.085 31.135 0.085 ;
      RECT 30.505 -0.085 30.675 0.085 ;
      RECT 30.045 -0.085 30.215 0.085 ;
      RECT 29.585 -0.085 29.755 0.085 ;
      RECT 29.125 -0.085 29.295 0.085 ;
      RECT 28.665 -0.085 28.835 0.085 ;
      RECT 28.205 -0.085 28.375 0.085 ;
      RECT 27.745 -0.085 27.915 0.085 ;
      RECT 27.285 -0.085 27.455 0.085 ;
      RECT 26.825 -0.085 26.995 0.085 ;
      RECT 26.365 -0.085 26.535 0.085 ;
      RECT 25.905 -0.085 26.075 0.085 ;
      RECT 25.445 -0.085 25.615 0.085 ;
      RECT 24.985 -0.085 25.155 0.085 ;
      RECT 24.525 -0.085 24.695 0.085 ;
      RECT 24.065 -0.085 24.235 0.085 ;
      RECT 23.605 -0.085 23.775 0.085 ;
      RECT 23.145 -0.085 23.315 0.085 ;
      RECT 22.685 -0.085 22.855 0.085 ;
      RECT 22.225 -0.085 22.395 0.085 ;
      RECT 21.765 -0.085 21.935 0.085 ;
      RECT 21.305 -0.085 21.475 0.085 ;
      RECT 20.845 -0.085 21.015 0.085 ;
      RECT 20.385 -0.085 20.555 0.085 ;
      RECT 19.925 -0.085 20.095 0.085 ;
      RECT 19.465 -0.085 19.635 0.085 ;
      RECT 19.005 -0.085 19.175 0.085 ;
      RECT 18.545 -0.085 18.715 0.085 ;
      RECT 18.085 -0.085 18.255 0.085 ;
      RECT 17.625 -0.085 17.795 0.085 ;
      RECT 17.165 -0.085 17.335 0.085 ;
      RECT 16.705 -0.085 16.875 0.085 ;
      RECT 16.245 -0.085 16.415 0.085 ;
      RECT 15.785 -0.085 15.955 0.085 ;
      RECT 15.325 -0.085 15.495 0.085 ;
      RECT 14.865 -0.085 15.035 0.085 ;
      RECT 14.405 -0.085 14.575 0.085 ;
      RECT 13.945 -0.085 14.115 0.085 ;
      RECT 13.485 -0.085 13.655 0.085 ;
      RECT 13.025 -0.085 13.195 0.085 ;
      RECT 12.565 -0.085 12.735 0.085 ;
      RECT 12.105 -0.085 12.275 0.085 ;
      RECT 11.645 -0.085 11.815 0.085 ;
      RECT 11.185 -0.085 11.355 0.085 ;
      RECT 10.725 -0.085 10.895 0.085 ;
      RECT 10.265 -0.085 10.435 0.085 ;
      RECT 9.805 -0.085 9.975 0.085 ;
      RECT 9.345 -0.085 9.515 0.085 ;
      RECT 8.885 -0.085 9.055 0.085 ;
      RECT 8.425 -0.085 8.595 0.085 ;
      RECT 7.965 -0.085 8.135 0.085 ;
      RECT 7.505 -0.085 7.675 0.085 ;
      RECT 7.045 -0.085 7.215 0.085 ;
      RECT 6.585 -0.085 6.755 0.085 ;
      RECT 6.125 -0.085 6.295 0.085 ;
      RECT 5.665 -0.085 5.835 0.085 ;
      RECT 5.205 -0.085 5.375 0.085 ;
      RECT 4.745 -0.085 4.915 0.085 ;
      RECT 4.285 -0.085 4.455 0.085 ;
      RECT 3.825 -0.085 3.995 0.085 ;
      RECT 3.365 -0.085 3.535 0.085 ;
      RECT 2.905 -0.085 3.075 0.085 ;
      RECT 2.445 -0.085 2.615 0.085 ;
      RECT 1.985 -0.085 2.155 0.085 ;
      RECT 1.525 -0.085 1.695 0.085 ;
      RECT 1.065 -0.085 1.235 0.085 ;
      RECT 0.605 -0.085 0.775 0.085 ;
      RECT 0.145 -0.085 0.315 0.085 ;
    LAYER via ;
      RECT 56.045 108.725 56.195 108.875 ;
      RECT 26.605 108.725 26.755 108.875 ;
      RECT 61.105 107.025 61.255 107.175 ;
      RECT 38.565 107.025 38.715 107.175 ;
      RECT 56.045 97.845 56.195 97.995 ;
      RECT 26.605 97.845 26.755 97.995 ;
      RECT 56.045 10.805 56.195 10.955 ;
      RECT 26.605 10.805 26.755 10.955 ;
      RECT 61.105 1.625 61.255 1.775 ;
      RECT 42.705 1.625 42.855 1.775 ;
      RECT 56.045 -0.075 56.195 0.075 ;
      RECT 26.605 -0.075 26.755 0.075 ;
    LAYER via2 ;
      RECT 56.02 108.7 56.22 108.9 ;
      RECT 26.58 108.7 26.78 108.9 ;
      RECT 94.2 88.3 94.4 88.5 ;
      RECT 94.2 86.94 94.4 87.14 ;
      RECT 94.2 65.86 94.4 66.06 ;
      RECT 94.2 49.54 94.4 49.74 ;
      RECT 94.2 45.46 94.4 45.66 ;
      RECT 94.2 37.3 94.4 37.5 ;
      RECT 56.02 -0.1 56.22 0.1 ;
      RECT 26.58 -0.1 26.78 0.1 ;
    LAYER via3 ;
      RECT 56.02 108.7 56.22 108.9 ;
      RECT 26.58 108.7 26.78 108.9 ;
      RECT 56.02 -0.1 56.22 0.1 ;
      RECT 26.58 -0.1 26.78 0.1 ;
    LAYER OVERLAP ;
      POLYGON 0 0 0 108.8 68.08 108.8 68.08 97.92 95.68 97.92 95.68 10.88 68.08 10.88 68.08 0 ;
  END
END sb_0__1_

END LIBRARY
