//
//
//
//
//
//
module direct_interc_5 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_6__5 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_4 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_5__4 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_3 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_4__3 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_2 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_3__2 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_1 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_2__1 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module direct_interc_0 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

sky130_fd_sc_hd__dlygate4sd3_1 FTB_1__0 ( .A ( in[0] ) , .X ( out[0] ) ) ;
endmodule


module mux_tree_tapbuf_size8_mem_3_2 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd1_1 FTB_17__56 ( .A ( mem_out[3] ) , 
    .X ( net_aps_56 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_RR_88 ( .A ( net_aps_56 ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size8_mem_2_3 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd1_1 FTB_16__55 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size8_mem_1_4 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd1_1 FTB_15__54 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size8_mem_0_4 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd1_1 FTB_14__53 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size8_mem_9 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd1_1 FTB_13__52 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size8_mem_6_2 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd1_1 FTB_12__51 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size8_mem_5_2 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd1_1 FTB_11__50 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size8_mem_4_2 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd1_1 FTB_10__49 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_44 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size8_3_2 ( in , sram , sram_inv , out , p0 ) ;
input  [0:7] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;

const1_44 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( in[2] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[4] ) , .A1 ( in[3] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[6] ) , .A1 ( in[5] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
endmodule


module const1_15_10 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size8_2_3 ( in , sram , sram_inv , out , p0 ) ;
input  [0:7] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;

const1_15_10 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( in[2] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[4] ) , .A1 ( in[3] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[6] ) , .A1 ( in[5] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
endmodule


module const1_14_11 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size8_1_4 ( in , sram , sram_inv , out , p0 ) ;
input  [0:7] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;

const1_14_11 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( in[2] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[4] ) , .A1 ( in[3] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[6] ) , .A1 ( in[5] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
endmodule


module const1_13_11 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size8_0_4 ( in , sram , sram_inv , out , p0 ) ;
input  [0:7] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;

const1_13_11 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( in[2] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[4] ) , .A1 ( in[3] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[6] ) , .A1 ( in[5] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_2 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[3] ) , .X ( out[0] ) ) ;
endmodule


module const1_12_11 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size8_9 ( in , sram , sram_inv , out , p0 ) ;
input  [0:7] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;

const1_12_11 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( in[2] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[4] ) , .A1 ( in[3] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[6] ) , .A1 ( in[5] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
endmodule


module const1_11_11 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size8_6_2 ( in , sram , sram_inv , out , p0 ) ;
input  [0:7] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;

const1_11_11 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( in[2] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[4] ) , .A1 ( in[3] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[6] ) , .A1 ( in[5] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
endmodule


module const1_10_11 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size8_5_2 ( in , sram , sram_inv , out , p0 ) ;
input  [0:7] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;

const1_10_11 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( in[2] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[4] ) , .A1 ( in[3] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[6] ) , .A1 ( in[5] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
endmodule


module const1_9_11 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size8_4_2 ( in , sram , sram_inv , out , p0 ) ;
input  [0:7] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;

const1_9_11 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( in[2] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[4] ) , .A1 ( in[3] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[6] ) , .A1 ( in[5] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
endmodule


module mux_tree_tapbuf_size10_mem_4_3 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd1_1 FTB_9__48 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size10_mem_3_3 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd1_1 FTB_8__47 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size10_mem_16 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd1_1 FTB_7__46 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size10_mem_7_2 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd1_1 FTB_6__45 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size10_mem_6_3 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd1_1 FTB_5__44 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size10_mem_5_3 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd1_1 FTB_4__43 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size10_mem_2_3 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd1_1 FTB_3__42 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size10_mem_1_3 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd1_1 FTB_2__41 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size10_mem_0_5 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd1_1 FTB_1__40 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_8_11 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size10_4_3 ( in , sram , sram_inv , out , p0 ) ;
input  [0:9] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

const1_8_11 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[6] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[8] ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[9] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
endmodule


module const1_7_11 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size10_3_3 ( in , sram , sram_inv , out , p0 ) ;
input  [0:9] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

const1_7_11 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[6] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[8] ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[9] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
endmodule


module const1_6_12 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size10_16 ( in , sram , sram_inv , out , p0 ) ;
input  [0:9] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

const1_6_12 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[6] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[8] ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[9] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
endmodule


module const1_5_12 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size10_7_2 ( in , sram , sram_inv , out , p0 ) ;
input  [0:9] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

const1_5_12 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[6] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[8] ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[9] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
endmodule


module const1_4_12 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size10_6_3 ( in , sram , sram_inv , out , p0 ) ;
input  [0:9] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

const1_4_12 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[6] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[8] ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[9] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
endmodule


module const1_3_12 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size10_5_3 ( in , sram , sram_inv , out , p0 ) ;
input  [0:9] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

const1_3_12 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[6] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[8] ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[9] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
endmodule


module const1_2_12 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size10_2_3 ( in , sram , sram_inv , out , p0 ) ;
input  [0:9] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

const1_2_12 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[6] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[8] ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[9] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
endmodule


module const1_1_12 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size10_1_3 ( in , sram , sram_inv , out , p0 ) ;
input  [0:9] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

const1_1_12 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[6] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[8] ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[9] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
endmodule


module const1_0_13 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size10_0_5 ( in , sram , sram_inv , out , p0 ) ;
input  [0:9] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

const1_0_13 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[6] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[8] ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[9] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
endmodule


module cby_1__1_ ( prog_clk , chany_bottom_in , chany_top_in , ccff_head , 
    chany_bottom_out , chany_top_out , right_grid_pin_52_ , left_grid_pin_0_ , 
    left_grid_pin_1_ , left_grid_pin_2_ , left_grid_pin_3_ , 
    left_grid_pin_4_ , left_grid_pin_5_ , left_grid_pin_6_ , 
    left_grid_pin_7_ , left_grid_pin_8_ , left_grid_pin_9_ , 
    left_grid_pin_10_ , left_grid_pin_11_ , left_grid_pin_12_ , 
    left_grid_pin_13_ , left_grid_pin_14_ , left_grid_pin_15_ , ccff_tail ) ;
input  [0:0] prog_clk ;
input  [0:19] chany_bottom_in ;
input  [0:19] chany_top_in ;
input  [0:0] ccff_head ;
output [0:19] chany_bottom_out ;
output [0:19] chany_top_out ;
output [0:0] right_grid_pin_52_ ;
output [0:0] left_grid_pin_0_ ;
output [0:0] left_grid_pin_1_ ;
output [0:0] left_grid_pin_2_ ;
output [0:0] left_grid_pin_3_ ;
output [0:0] left_grid_pin_4_ ;
output [0:0] left_grid_pin_5_ ;
output [0:0] left_grid_pin_6_ ;
output [0:0] left_grid_pin_7_ ;
output [0:0] left_grid_pin_8_ ;
output [0:0] left_grid_pin_9_ ;
output [0:0] left_grid_pin_10_ ;
output [0:0] left_grid_pin_11_ ;
output [0:0] left_grid_pin_12_ ;
output [0:0] left_grid_pin_13_ ;
output [0:0] left_grid_pin_14_ ;
output [0:0] left_grid_pin_15_ ;
output [0:0] ccff_tail ;

wire [0:3] mux_tree_tapbuf_size10_0_sram ;
wire [0:3] mux_tree_tapbuf_size10_0_sram_inv ;
wire [0:3] mux_tree_tapbuf_size10_1_sram ;
wire [0:3] mux_tree_tapbuf_size10_1_sram_inv ;
wire [0:3] mux_tree_tapbuf_size10_2_sram ;
wire [0:3] mux_tree_tapbuf_size10_2_sram_inv ;
wire [0:3] mux_tree_tapbuf_size10_3_sram ;
wire [0:3] mux_tree_tapbuf_size10_3_sram_inv ;
wire [0:3] mux_tree_tapbuf_size10_4_sram ;
wire [0:3] mux_tree_tapbuf_size10_4_sram_inv ;
wire [0:3] mux_tree_tapbuf_size10_5_sram ;
wire [0:3] mux_tree_tapbuf_size10_5_sram_inv ;
wire [0:3] mux_tree_tapbuf_size10_6_sram ;
wire [0:3] mux_tree_tapbuf_size10_6_sram_inv ;
wire [0:3] mux_tree_tapbuf_size10_7_sram ;
wire [0:3] mux_tree_tapbuf_size10_7_sram_inv ;
wire [0:3] mux_tree_tapbuf_size10_8_sram ;
wire [0:3] mux_tree_tapbuf_size10_8_sram_inv ;
wire [0:0] mux_tree_tapbuf_size10_mem_0_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size10_mem_1_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size10_mem_2_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size10_mem_3_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size10_mem_4_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size10_mem_5_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size10_mem_6_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size10_mem_7_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size10_mem_8_ccff_tail ;
wire [0:3] mux_tree_tapbuf_size8_0_sram ;
wire [0:3] mux_tree_tapbuf_size8_0_sram_inv ;
wire [0:3] mux_tree_tapbuf_size8_1_sram ;
wire [0:3] mux_tree_tapbuf_size8_1_sram_inv ;
wire [0:3] mux_tree_tapbuf_size8_2_sram ;
wire [0:3] mux_tree_tapbuf_size8_2_sram_inv ;
wire [0:3] mux_tree_tapbuf_size8_3_sram ;
wire [0:3] mux_tree_tapbuf_size8_3_sram_inv ;
wire [0:3] mux_tree_tapbuf_size8_4_sram ;
wire [0:3] mux_tree_tapbuf_size8_4_sram_inv ;
wire [0:3] mux_tree_tapbuf_size8_5_sram ;
wire [0:3] mux_tree_tapbuf_size8_5_sram_inv ;
wire [0:3] mux_tree_tapbuf_size8_6_sram ;
wire [0:3] mux_tree_tapbuf_size8_6_sram_inv ;
wire [0:3] mux_tree_tapbuf_size8_7_sram ;
wire [0:3] mux_tree_tapbuf_size8_7_sram_inv ;
wire [0:0] mux_tree_tapbuf_size8_mem_0_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size8_mem_1_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size8_mem_2_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size8_mem_3_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size8_mem_4_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size8_mem_5_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size8_mem_6_ccff_tail ;

mux_tree_tapbuf_size10_0_5 mux_left_ipin_0 (
    .in ( { chany_bottom_in[0] , chany_top_in[0] , chany_bottom_in[2] , 
        chany_top_in[2] , chany_bottom_in[4] , chany_top_in[4] , 
        chany_bottom_in[10] , chany_top_in[10] , chany_bottom_in[16] , 
        chany_top_in[16] } ) ,
    .sram ( mux_tree_tapbuf_size10_0_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size10_0_sram_inv ) , 
    .out ( right_grid_pin_52_ ) , .p0 ( optlc_net_112 ) ) ;
mux_tree_tapbuf_size10_1_3 mux_right_ipin_0 (
    .in ( { chany_bottom_in[1] , chany_top_in[1] , chany_bottom_in[3] , 
        chany_top_in[3] , chany_bottom_in[5] , chany_top_in[5] , 
        chany_bottom_in[11] , chany_top_in[11] , chany_bottom_in[17] , 
        chany_top_in[17] } ) ,
    .sram ( mux_tree_tapbuf_size10_1_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size10_1_sram_inv ) , 
    .out ( left_grid_pin_0_ ) , .p0 ( optlc_net_111 ) ) ;
mux_tree_tapbuf_size10_2_3 mux_right_ipin_1 (
    .in ( { chany_bottom_in[0] , chany_top_in[0] , chany_bottom_in[2] , 
        chany_top_in[2] , chany_bottom_in[6] , chany_top_in[6] , 
        chany_bottom_in[12] , chany_top_in[12] , chany_bottom_in[18] , 
        chany_top_in[18] } ) ,
    .sram ( mux_tree_tapbuf_size10_2_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size10_2_sram_inv ) , 
    .out ( left_grid_pin_1_ ) , .p0 ( optlc_net_111 ) ) ;
mux_tree_tapbuf_size10_5_3 mux_right_ipin_4 (
    .in ( { chany_bottom_in[1] , chany_top_in[1] , chany_bottom_in[3] , 
        chany_top_in[3] , chany_bottom_in[5] , chany_top_in[5] , 
        chany_bottom_in[9] , chany_top_in[9] , chany_bottom_in[15] , 
        chany_top_in[15] } ) ,
    .sram ( mux_tree_tapbuf_size10_3_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size10_3_sram_inv ) , 
    .out ( left_grid_pin_4_ ) , .p0 ( optlc_net_111 ) ) ;
mux_tree_tapbuf_size10_6_3 mux_right_ipin_5 (
    .in ( { chany_bottom_in[0] , chany_top_in[0] , chany_bottom_in[2] , 
        chany_top_in[2] , chany_bottom_in[6] , chany_top_in[6] , 
        chany_bottom_in[10] , chany_top_in[10] , chany_bottom_in[16] , 
        chany_top_in[16] } ) ,
    .sram ( mux_tree_tapbuf_size10_4_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size10_4_sram_inv ) , 
    .out ( left_grid_pin_5_ ) , .p0 ( optlc_net_109 ) ) ;
mux_tree_tapbuf_size10_7_2 mux_right_ipin_8 (
    .in ( { chany_bottom_in[1] , chany_top_in[1] , chany_bottom_in[3] , 
        chany_top_in[3] , chany_bottom_in[9] , chany_top_in[9] , 
        chany_bottom_in[13] , chany_top_in[13] , chany_bottom_in[19] , 
        chany_top_in[19] } ) ,
    .sram ( mux_tree_tapbuf_size10_5_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size10_5_sram_inv ) , 
    .out ( left_grid_pin_8_ ) , .p0 ( optlc_net_111 ) ) ;
mux_tree_tapbuf_size10_16 mux_right_ipin_9 (
    .in ( { chany_bottom_in[0] , chany_top_in[0] , chany_bottom_in[2] , 
        chany_top_in[2] , chany_bottom_in[4] , chany_top_in[4] , 
        chany_bottom_in[10] , chany_top_in[10] , chany_bottom_in[14] , 
        chany_top_in[14] } ) ,
    .sram ( mux_tree_tapbuf_size10_6_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size10_6_sram_inv ) , 
    .out ( left_grid_pin_9_ ) , .p0 ( optlc_net_109 ) ) ;
mux_tree_tapbuf_size10_3_3 mux_right_ipin_12 (
    .in ( { chany_bottom_in[1] , chany_top_in[1] , chany_bottom_in[3] , 
        chany_top_in[3] , chany_bottom_in[7] , chany_top_in[7] , 
        chany_bottom_in[13] , chany_top_in[13] , chany_bottom_in[17] , 
        chany_top_in[17] } ) ,
    .sram ( mux_tree_tapbuf_size10_7_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size10_7_sram_inv ) , 
    .out ( left_grid_pin_12_ ) , .p0 ( optlc_net_110 ) ) ;
mux_tree_tapbuf_size10_4_3 mux_right_ipin_13 (
    .in ( { chany_bottom_in[0] , chany_top_in[0] , chany_bottom_in[2] , 
        chany_top_in[2] , chany_bottom_in[8] , chany_top_in[8] , 
        chany_bottom_in[14] , chany_top_in[14] , chany_bottom_in[18] , 
        chany_top_in[18] } ) ,
    .sram ( mux_tree_tapbuf_size10_8_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size10_8_sram_inv ) , 
    .out ( left_grid_pin_13_ ) , .p0 ( optlc_net_109 ) ) ;
mux_tree_tapbuf_size10_mem_0_5 mem_left_ipin_0 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( ccff_head ) , 
    .ccff_tail ( mux_tree_tapbuf_size10_mem_0_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size10_0_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size10_0_sram_inv ) ) ;
mux_tree_tapbuf_size10_mem_1_3 mem_right_ipin_0 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size10_mem_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size10_mem_1_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size10_1_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size10_1_sram_inv ) ) ;
mux_tree_tapbuf_size10_mem_2_3 mem_right_ipin_1 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size10_mem_1_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size10_mem_2_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size10_2_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size10_2_sram_inv ) ) ;
mux_tree_tapbuf_size10_mem_5_3 mem_right_ipin_4 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size8_mem_1_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size10_mem_3_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size10_3_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size10_3_sram_inv ) ) ;
mux_tree_tapbuf_size10_mem_6_3 mem_right_ipin_5 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size10_mem_3_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size10_mem_4_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size10_4_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size10_4_sram_inv ) ) ;
mux_tree_tapbuf_size10_mem_7_2 mem_right_ipin_8 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size8_mem_3_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size10_mem_5_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size10_5_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size10_5_sram_inv ) ) ;
mux_tree_tapbuf_size10_mem_16 mem_right_ipin_9 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size10_mem_5_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size10_mem_6_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size10_6_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size10_6_sram_inv ) ) ;
mux_tree_tapbuf_size10_mem_3_3 mem_right_ipin_12 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size8_mem_5_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size10_mem_7_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size10_7_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size10_7_sram_inv ) ) ;
mux_tree_tapbuf_size10_mem_4_3 mem_right_ipin_13 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size10_mem_7_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size10_mem_8_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size10_8_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size10_8_sram_inv ) ) ;
mux_tree_tapbuf_size8_4_2 mux_right_ipin_2 (
    .in ( { chany_bottom_in[1] , chany_top_in[1] , chany_bottom_in[3] , 
        chany_top_in[3] , chany_bottom_in[7] , chany_top_in[7] , 
        chany_bottom_in[15] , chany_top_in[15] } ) ,
    .sram ( mux_tree_tapbuf_size8_0_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size8_0_sram_inv ) , 
    .out ( left_grid_pin_2_ ) , .p0 ( optlc_net_111 ) ) ;
mux_tree_tapbuf_size8_5_2 mux_right_ipin_3 (
    .in ( { chany_bottom_in[0] , chany_top_in[0] , chany_bottom_in[2] , 
        chany_top_in[2] , chany_bottom_in[8] , chany_top_in[8] , 
        chany_bottom_in[16] , chany_top_in[16] } ) ,
    .sram ( mux_tree_tapbuf_size8_1_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size8_1_sram_inv ) , 
    .out ( left_grid_pin_3_ ) , .p0 ( optlc_net_112 ) ) ;
mux_tree_tapbuf_size8_6_2 mux_right_ipin_6 (
    .in ( { chany_bottom_in[1] , chany_top_in[1] , chany_bottom_in[3] , 
        chany_top_in[3] , chany_bottom_in[11] , chany_top_in[11] , 
        chany_bottom_in[19] , chany_top_in[19] } ) ,
    .sram ( mux_tree_tapbuf_size8_2_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size8_2_sram_inv ) , 
    .out ( left_grid_pin_6_ ) , .p0 ( optlc_net_110 ) ) ;
mux_tree_tapbuf_size8_9 mux_right_ipin_7 (
    .in ( { chany_bottom_in[0] , chany_top_in[0] , chany_bottom_in[2] , 
        chany_top_in[2] , chany_bottom_in[4] , chany_top_in[4] , 
        chany_bottom_in[12] , chany_top_in[12] } ) ,
    .sram ( mux_tree_tapbuf_size8_3_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size8_3_sram_inv ) , 
    .out ( left_grid_pin_7_ ) , .p0 ( optlc_net_112 ) ) ;
mux_tree_tapbuf_size8_0_4 mux_right_ipin_10 (
    .in ( { chany_bottom_in[1] , chany_top_in[1] , chany_bottom_in[3] , 
        chany_top_in[3] , chany_bottom_in[7] , chany_top_in[7] , 
        chany_bottom_in[15] , chany_top_in[15] } ) ,
    .sram ( mux_tree_tapbuf_size8_4_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size8_4_sram_inv ) , 
    .out ( left_grid_pin_10_ ) , .p0 ( optlc_net_109 ) ) ;
mux_tree_tapbuf_size8_1_4 mux_right_ipin_11 (
    .in ( { chany_bottom_in[0] , chany_top_in[0] , chany_bottom_in[2] , 
        chany_top_in[2] , chany_bottom_in[8] , chany_top_in[8] , 
        chany_bottom_in[16] , chany_top_in[16] } ) ,
    .sram ( mux_tree_tapbuf_size8_5_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size8_5_sram_inv ) , 
    .out ( left_grid_pin_11_ ) , .p0 ( optlc_net_109 ) ) ;
mux_tree_tapbuf_size8_2_3 mux_right_ipin_14 (
    .in ( { chany_bottom_in[1] , chany_top_in[1] , chany_bottom_in[3] , 
        chany_top_in[3] , chany_bottom_in[11] , chany_top_in[11] , 
        chany_bottom_in[19] , chany_top_in[19] } ) ,
    .sram ( mux_tree_tapbuf_size8_6_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size8_6_sram_inv ) , 
    .out ( left_grid_pin_14_ ) , .p0 ( optlc_net_110 ) ) ;
mux_tree_tapbuf_size8_3_2 mux_right_ipin_15 (
    .in ( { chany_bottom_in[0] , chany_top_in[0] , chany_bottom_in[2] , 
        chany_top_in[2] , chany_bottom_in[4] , chany_top_in[4] , 
        chany_bottom_in[12] , chany_top_in[12] } ) ,
    .sram ( mux_tree_tapbuf_size8_7_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size8_7_sram_inv ) , 
    .out ( left_grid_pin_15_ ) , .p0 ( optlc_net_112 ) ) ;
mux_tree_tapbuf_size8_mem_4_2 mem_right_ipin_2 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size10_mem_2_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size8_mem_0_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size8_0_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size8_0_sram_inv ) ) ;
mux_tree_tapbuf_size8_mem_5_2 mem_right_ipin_3 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size8_mem_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size8_mem_1_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size8_1_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size8_1_sram_inv ) ) ;
mux_tree_tapbuf_size8_mem_6_2 mem_right_ipin_6 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size10_mem_4_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size8_mem_2_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size8_2_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size8_2_sram_inv ) ) ;
mux_tree_tapbuf_size8_mem_9 mem_right_ipin_7 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size8_mem_2_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size8_mem_3_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size8_3_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size8_3_sram_inv ) ) ;
mux_tree_tapbuf_size8_mem_0_4 mem_right_ipin_10 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size10_mem_6_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size8_mem_4_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size8_4_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size8_4_sram_inv ) ) ;
mux_tree_tapbuf_size8_mem_1_4 mem_right_ipin_11 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size8_mem_4_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size8_mem_5_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size8_5_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size8_5_sram_inv ) ) ;
mux_tree_tapbuf_size8_mem_2_3 mem_right_ipin_14 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size10_mem_8_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size8_mem_6_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size8_6_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size8_6_sram_inv ) ) ;
mux_tree_tapbuf_size8_mem_3_2 mem_right_ipin_15 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size8_mem_6_ccff_tail ) , 
    .ccff_tail ( ccff_tail ) , .mem_out ( mux_tree_tapbuf_size8_7_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size8_7_sram_inv ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_689 ( .A ( ropt_net_113 ) , 
    .X ( chany_top_out[11] ) ) ;
sky130_fd_sc_hd__dlygate4sd1_1 FTB_2__1 ( .A ( chany_bottom_in[1] ) , 
    .X ( chany_top_out[1] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_3__2 ( .A ( chany_bottom_in[2] ) , 
    .X ( chany_top_out[2] ) ) ;
sky130_fd_sc_hd__conb_1 optlc_104 ( .LO ( SYNOPSYS_UNCONNECTED_1 ) , 
    .HI ( optlc_net_109 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_5__4 ( .A ( chany_bottom_in[4] ) , 
    .X ( chany_top_out[4] ) ) ;
sky130_fd_sc_hd__dlygate4sd1_1 FTB_6__5 ( .A ( chany_bottom_in[5] ) , 
    .X ( chany_top_out[5] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_7__6 ( .A ( chany_bottom_in[6] ) , 
    .X ( chany_top_out[6] ) ) ;
sky130_fd_sc_hd__conb_1 optlc_106 ( .LO ( SYNOPSYS_UNCONNECTED_2 ) , 
    .HI ( optlc_net_110 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_9__8 ( .A ( chany_bottom_in[8] ) , 
    .X ( chany_top_out[8] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_10__9 ( .A ( chany_bottom_in[9] ) , 
    .X ( aps_rename_1_ ) ) ;
sky130_fd_sc_hd__conb_1 optlc_108 ( .LO ( SYNOPSYS_UNCONNECTED_3 ) , 
    .HI ( optlc_net_111 ) ) ;
sky130_fd_sc_hd__dlygate4sd1_1 FTB_12__11 ( .A ( chany_bottom_in[11] ) , 
    .X ( ropt_net_113 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_110 ( .LO ( SYNOPSYS_UNCONNECTED_4 ) , 
    .HI ( optlc_net_112 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_14__13 ( .A ( chany_bottom_in[13] ) , 
    .X ( aps_rename_2_ ) ) ;
sky130_fd_sc_hd__dlygate4sd1_1 FTB_16__15 ( .A ( chany_bottom_in[15] ) , 
    .X ( chany_top_out[15] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_17__16 ( .A ( chany_bottom_in[16] ) , 
    .X ( aps_rename_4_ ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_18__17 ( .A ( chany_bottom_in[17] ) , 
    .X ( aps_rename_5_ ) ) ;
sky130_fd_sc_hd__dlygate4sd1_1 FTB_21__20 ( .A ( chany_top_in[0] ) , 
    .X ( chany_bottom_out[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd1_1 FTB_22__21 ( .A ( chany_top_in[1] ) , 
    .X ( chany_bottom_out[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd1_1 FTB_23__22 ( .A ( chany_top_in[2] ) , 
    .X ( chany_bottom_out[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd1_1 FTB_24__23 ( .A ( chany_top_in[3] ) , 
    .X ( chany_bottom_out[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd1_1 FTB_25__24 ( .A ( chany_top_in[4] ) , 
    .X ( chany_bottom_out[4] ) ) ;
sky130_fd_sc_hd__dlygate4sd1_1 FTB_27__26 ( .A ( chany_top_in[6] ) , 
    .X ( chany_bottom_out[6] ) ) ;
sky130_fd_sc_hd__dlygate4sd1_1 FTB_28__27 ( .A ( chany_top_in[7] ) , 
    .X ( chany_bottom_out[7] ) ) ;
sky130_fd_sc_hd__dlygate4sd1_1 FTB_29__28 ( .A ( chany_top_in[8] ) , 
    .X ( chany_bottom_out[8] ) ) ;
sky130_fd_sc_hd__dlygate4sd1_1 FTB_33__32 ( .A ( chany_top_in[12] ) , 
    .X ( chany_bottom_out[12] ) ) ;
sky130_fd_sc_hd__dlygate4sd1_1 FTB_34__33 ( .A ( chany_top_in[13] ) , 
    .X ( chany_bottom_out[13] ) ) ;
sky130_fd_sc_hd__dlygate4sd1_1 FTB_35__34 ( .A ( chany_top_in[14] ) , 
    .X ( chany_bottom_out[14] ) ) ;
sky130_fd_sc_hd__dlygate4sd1_1 FTB_36__35 ( .A ( chany_top_in[15] ) , 
    .X ( chany_bottom_out[15] ) ) ;
sky130_fd_sc_hd__dlygate4sd1_1 FTB_38__37 ( .A ( chany_top_in[17] ) , 
    .X ( chany_bottom_out[17] ) ) ;
sky130_fd_sc_hd__dlygate4sd1_1 FTB_40__39 ( .A ( chany_top_in[19] ) , 
    .X ( chany_bottom_out[19] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_RR_61 ( .A ( chany_bottom_in[3] ) , 
    .X ( chany_top_out[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_68 ( .A ( chany_bottom_in[19] ) , 
    .X ( BUF_net_68 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_71 ( .A ( chany_top_in[16] ) , 
    .X ( BUF_net_71 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_RR_73 ( .A ( chany_bottom_in[7] ) , 
    .X ( chany_top_out[7] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_RR_74 ( .A ( chany_bottom_in[10] ) , 
    .X ( chany_top_out[10] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_RR_77 ( .A ( chany_bottom_in[0] ) , 
    .X ( chany_top_out[0] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 BUFT_RR_78 ( .A ( aps_rename_1_ ) , 
    .X ( chany_top_out[9] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 BUFT_RR_79 ( .A ( aps_rename_2_ ) , 
    .X ( chany_top_out[13] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_RR_80 ( .A ( chany_bottom_in[14] ) , 
    .X ( chany_top_out[14] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 BUFT_RR_81 ( .A ( aps_rename_4_ ) , 
    .X ( chany_top_out[16] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 BUFT_RR_82 ( .A ( aps_rename_5_ ) , 
    .X ( chany_top_out[17] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_RR_86 ( .A ( chany_top_in[9] ) , 
    .X ( chany_bottom_out[9] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_P_93 ( .A ( chany_bottom_in[12] ) , 
    .X ( chany_top_out[12] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_P_94 ( .A ( chany_top_in[10] ) , 
    .X ( chany_bottom_out[10] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_P_95 ( .A ( chany_top_in[11] ) , 
    .X ( chany_bottom_out[11] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_P_96 ( .A ( chany_top_in[18] ) , 
    .X ( chany_bottom_out[18] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_P_97 ( .A ( chany_bottom_in[18] ) , 
    .X ( chany_top_out[18] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 BUFT_P_98 ( .A ( BUF_net_68 ) , 
    .X ( chany_top_out[19] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_P_99 ( .A ( chany_top_in[5] ) , 
    .X ( chany_bottom_out[5] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 BUFT_P_101 ( .A ( BUF_net_71 ) , 
    .X ( chany_bottom_out[16] ) ) ;
endmodule


module mux_tree_tapbuf_size10_mem_15 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_2__41 ( .A ( mem_out[3] ) , 
    .X ( net_net_76 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 BUFT_RR_114 ( .A ( net_net_76 ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size10_mem_0_4 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_1__40 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_43 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size10_15 ( in , sram , sram_inv , out , p0 ) ;
input  [0:9] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

const1_43 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[6] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[8] ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[9] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
endmodule


module const1_0_12 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size10_0_4 ( in , sram , sram_inv , out , p0 ) ;
input  [0:9] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

const1_0_12 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[6] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[8] ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[9] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
endmodule


module cby_0__1_ ( prog_clk , chany_bottom_in , chany_top_in , ccff_head , 
    chany_bottom_out , chany_top_out , right_grid_pin_52_ , left_grid_pin_0_ , 
    ccff_tail ) ;
input  [0:0] prog_clk ;
input  [0:19] chany_bottom_in ;
input  [0:19] chany_top_in ;
input  [0:0] ccff_head ;
output [0:19] chany_bottom_out ;
output [0:19] chany_top_out ;
output [0:0] right_grid_pin_52_ ;
output [0:0] left_grid_pin_0_ ;
output [0:0] ccff_tail ;

wire [0:3] mux_tree_tapbuf_size10_0_sram ;
wire [0:3] mux_tree_tapbuf_size10_0_sram_inv ;
wire [0:3] mux_tree_tapbuf_size10_1_sram ;
wire [0:3] mux_tree_tapbuf_size10_1_sram_inv ;
wire [0:0] mux_tree_tapbuf_size10_mem_0_ccff_tail ;

mux_tree_tapbuf_size10_0_4 mux_left_ipin_0 (
    .in ( { chany_bottom_in[0] , chany_top_in[0] , chany_bottom_in[2] , 
        chany_top_in[2] , chany_bottom_in[4] , chany_top_in[4] , 
        chany_bottom_in[10] , chany_top_in[10] , chany_bottom_in[16] , 
        chany_top_in[16] } ) ,
    .sram ( mux_tree_tapbuf_size10_0_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size10_0_sram_inv ) , 
    .out ( right_grid_pin_52_ ) , .p0 ( optlc_net_144 ) ) ;
mux_tree_tapbuf_size10_15 mux_right_ipin_0 (
    .in ( { chany_bottom_in[1] , chany_top_in[1] , chany_bottom_in[3] , 
        chany_top_in[3] , chany_bottom_in[5] , chany_top_in[5] , 
        chany_bottom_in[11] , chany_top_in[11] , chany_bottom_in[17] , 
        chany_top_in[17] } ) ,
    .sram ( mux_tree_tapbuf_size10_1_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size10_1_sram_inv ) , 
    .out ( left_grid_pin_0_ ) , .p0 ( optlc_net_145 ) ) ;
mux_tree_tapbuf_size10_mem_0_4 mem_left_ipin_0 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( ccff_head ) , 
    .ccff_tail ( mux_tree_tapbuf_size10_mem_0_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size10_0_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size10_0_sram_inv ) ) ;
mux_tree_tapbuf_size10_mem_15 mem_right_ipin_0 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size10_mem_0_ccff_tail ) , 
    .ccff_tail ( ccff_tail ) , .mem_out ( mux_tree_tapbuf_size10_1_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size10_1_sram_inv ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_1__0 ( .A ( chany_bottom_in[0] ) , 
    .X ( chany_top_out[0] ) ) ;
sky130_fd_sc_hd__conb_1 optlc_144 ( .LO ( SYNOPSYS_UNCONNECTED_1 ) , 
    .HI ( optlc_net_144 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_3__2 ( .A ( chany_bottom_in[2] ) , 
    .X ( ropt_net_173 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_145 ( .LO ( SYNOPSYS_UNCONNECTED_2 ) , 
    .HI ( optlc_net_145 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_724 ( .A ( chany_bottom_in[8] ) , 
    .X ( ropt_net_202 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_758 ( .A ( ropt_net_177 ) , 
    .X ( chany_bottom_out[1] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_759 ( .A ( ropt_net_178 ) , 
    .X ( chany_bottom_out[2] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_8__7 ( .A ( chany_bottom_in[7] ) , 
    .X ( chany_top_out[7] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_725 ( .A ( chany_bottom_in[6] ) , 
    .X ( ropt_net_201 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_726 ( .A ( chany_bottom_in[5] ) , 
    .X ( ropt_net_182 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_727 ( .A ( chany_top_in[18] ) , 
    .X ( chany_bottom_out[18] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_728 ( .A ( chany_top_in[5] ) , 
    .X ( ropt_net_200 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_729 ( .A ( ropt_net_151 ) , 
    .X ( chany_bottom_out[8] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_730 ( .A ( chany_top_in[13] ) , 
    .X ( ropt_net_199 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_731 ( .A ( ropt_net_153 ) , 
    .X ( ropt_net_178 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_732 ( .A ( ropt_net_154 ) , 
    .X ( ropt_net_177 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_733 ( .A ( ropt_net_155 ) , 
    .X ( ropt_net_181 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_734 ( .A ( ropt_net_156 ) , 
    .X ( ropt_net_187 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_735 ( .A ( ropt_net_157 ) , 
    .X ( ropt_net_186 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_736 ( .A ( ropt_net_158 ) , 
    .X ( ropt_net_184 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_21__20 ( .A ( chany_top_in[0] ) , 
    .X ( ropt_net_204 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_737 ( .A ( ropt_net_159 ) , 
    .X ( ropt_net_198 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_738 ( .A ( ropt_net_160 ) , 
    .X ( chany_bottom_out[15] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_739 ( .A ( ropt_net_161 ) , 
    .X ( ropt_net_189 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_25__24 ( .A ( chany_top_in[4] ) , 
    .X ( ropt_net_169 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_740 ( .A ( ropt_net_162 ) , 
    .X ( chany_bottom_out[19] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_741 ( .A ( ropt_net_163 ) , 
    .X ( chany_bottom_out[10] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_742 ( .A ( ropt_net_164 ) , 
    .X ( ropt_net_195 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_743 ( .A ( ropt_net_165 ) , 
    .X ( ropt_net_193 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_744 ( .A ( ropt_net_166 ) , 
    .X ( ropt_net_190 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_745 ( .A ( ropt_net_167 ) , 
    .X ( ropt_net_183 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_746 ( .A ( ropt_net_168 ) , 
    .X ( ropt_net_179 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_747 ( .A ( ropt_net_169 ) , 
    .X ( ropt_net_192 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_748 ( .A ( ropt_net_170 ) , 
    .X ( ropt_net_185 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_749 ( .A ( ropt_net_171 ) , 
    .X ( ropt_net_191 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_750 ( .A ( ropt_net_172 ) , 
    .X ( ropt_net_196 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_751 ( .A ( ropt_net_173 ) , 
    .X ( ropt_net_180 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_752 ( .A ( ropt_net_174 ) , 
    .X ( ropt_net_194 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_754 ( .A ( ropt_net_175 ) , 
    .X ( ropt_net_188 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_755 ( .A ( ropt_net_176 ) , 
    .X ( ropt_net_197 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_760 ( .A ( ropt_net_179 ) , 
    .X ( chany_bottom_out[6] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_761 ( .A ( ropt_net_180 ) , 
    .X ( chany_top_out[2] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_762 ( .A ( ropt_net_181 ) , 
    .X ( chany_top_out[16] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_RR_45 ( .A ( chany_bottom_in[3] ) , 
    .X ( chany_top_out[3] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_763 ( .A ( ropt_net_182 ) , 
    .X ( chany_top_out[5] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_764 ( .A ( ropt_net_183 ) , 
    .X ( chany_top_out[13] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_765 ( .A ( ropt_net_184 ) , 
    .X ( chany_bottom_out[12] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_766 ( .A ( ropt_net_185 ) , 
    .X ( chany_bottom_out[11] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_767 ( .A ( ropt_net_186 ) , 
    .X ( chany_top_out[19] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_51 ( .A ( chany_bottom_in[10] ) , 
    .X ( ropt_net_175 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_769 ( .A ( ropt_net_187 ) , 
    .X ( chany_top_out[15] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_770 ( .A ( ropt_net_188 ) , 
    .X ( chany_top_out[10] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_771 ( .A ( ropt_net_189 ) , 
    .X ( chany_top_out[18] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_772 ( .A ( ropt_net_190 ) , 
    .X ( chany_top_out[4] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_773 ( .A ( ropt_net_191 ) , 
    .X ( chany_bottom_out[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_57 ( .A ( chany_bottom_in[17] ) , 
    .X ( ropt_net_165 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_58 ( .A ( chany_bottom_in[19] ) , 
    .X ( ropt_net_157 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_59 ( .A ( chany_top_in[1] ) , 
    .X ( ropt_net_154 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_60 ( .A ( chany_top_in[2] ) , 
    .X ( ropt_net_153 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_774 ( .A ( ropt_net_192 ) , 
    .X ( chany_bottom_out[4] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_775 ( .A ( ropt_net_193 ) , 
    .X ( chany_top_out[17] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_776 ( .A ( ropt_net_194 ) , 
    .X ( chany_top_out[12] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_64 ( .A ( chany_top_in[7] ) , 
    .X ( ropt_net_164 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_RR_65 ( .A ( chany_top_in[8] ) , 
    .X ( ropt_net_151 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_66 ( .A ( chany_top_in[9] ) , 
    .X ( BUF_net_66 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_777 ( .A ( ropt_net_195 ) , 
    .X ( chany_bottom_out[7] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_68 ( .A ( chany_top_in[11] ) , 
    .X ( ropt_net_170 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_69 ( .A ( chany_top_in[12] ) , 
    .X ( ropt_net_158 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_778 ( .A ( ropt_net_196 ) , 
    .X ( chany_top_out[11] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_779 ( .A ( ropt_net_197 ) , 
    .X ( chany_top_out[14] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_780 ( .A ( ropt_net_198 ) , 
    .X ( chany_top_out[9] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_RR_73 ( .A ( chany_top_in[17] ) , 
    .X ( chany_bottom_out[17] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_783 ( .A ( ropt_net_199 ) , 
    .X ( chany_bottom_out[13] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_787 ( .A ( ropt_net_200 ) , 
    .X ( chany_bottom_out[5] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_789 ( .A ( ropt_net_201 ) , 
    .X ( chany_top_out[6] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_790 ( .A ( ropt_net_202 ) , 
    .X ( chany_top_out[8] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_792 ( .A ( ropt_net_203 ) , 
    .X ( chany_bottom_out[16] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_794 ( .A ( ropt_net_204 ) , 
    .X ( chany_bottom_out[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_95 ( .A ( chany_top_in[3] ) , 
    .X ( ropt_net_171 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_RR_101 ( .A ( chany_top_in[10] ) , 
    .X ( ropt_net_163 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_P_110 ( .A ( chany_bottom_in[16] ) , 
    .X ( ropt_net_155 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_P_111 ( .A ( chany_bottom_in[18] ) , 
    .X ( ropt_net_161 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_P_112 ( .A ( chany_top_in[16] ) , 
    .X ( ropt_net_203 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_P_113 ( .A ( chany_top_in[19] ) , 
    .X ( ropt_net_162 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_P_115 ( .A ( chany_bottom_in[1] ) , 
    .X ( chany_top_out[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_P_117 ( .A ( chany_bottom_in[4] ) , 
    .X ( ropt_net_166 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_P_119 ( .A ( chany_bottom_in[9] ) , 
    .X ( ropt_net_159 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_P_120 ( .A ( chany_bottom_in[11] ) , 
    .X ( ropt_net_172 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_P_121 ( .A ( chany_bottom_in[12] ) , 
    .X ( ropt_net_174 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_P_122 ( .A ( chany_bottom_in[13] ) , 
    .X ( ropt_net_167 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_P_123 ( .A ( chany_bottom_in[14] ) , 
    .X ( ropt_net_176 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_P_124 ( .A ( chany_bottom_in[15] ) , 
    .X ( ropt_net_156 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_P_131 ( .A ( chany_top_in[6] ) , 
    .X ( ropt_net_168 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 BUFT_P_134 ( .A ( BUF_net_66 ) , 
    .X ( chany_bottom_out[9] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_P_139 ( .A ( chany_top_in[14] ) , 
    .X ( chany_bottom_out[14] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_P_140 ( .A ( chany_top_in[15] ) , 
    .X ( ropt_net_160 ) ) ;
endmodule


module mux_tree_tapbuf_size10_mem_14 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_1__40 ( .A ( mem_out[3] ) , 
    .X ( net_net_74 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_115 ( .A ( net_net_74 ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_42 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size10_14 ( in , sram , sram_inv , out , p0 ) ;
input  [0:9] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

const1_42 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[6] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[8] ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[9] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
endmodule


module cbx_1__2_ ( prog_clk , chanx_left_in , chanx_right_in , ccff_head , 
    chanx_left_out , chanx_right_out , top_grid_pin_0_ , ccff_tail ) ;
input  [0:0] prog_clk ;
input  [0:19] chanx_left_in ;
input  [0:19] chanx_right_in ;
input  [0:0] ccff_head ;
output [0:19] chanx_left_out ;
output [0:19] chanx_right_out ;
output [0:0] top_grid_pin_0_ ;
output [0:0] ccff_tail ;

wire [0:3] mux_tree_tapbuf_size10_0_sram ;
wire [0:3] mux_tree_tapbuf_size10_0_sram_inv ;

mux_tree_tapbuf_size10_14 mux_bottom_ipin_0 (
    .in ( { chanx_left_in[0] , chanx_right_in[0] , chanx_left_in[2] , 
        chanx_right_in[2] , chanx_left_in[4] , chanx_right_in[4] , 
        chanx_left_in[10] , chanx_right_in[10] , chanx_left_in[16] , 
        chanx_right_in[16] } ) ,
    .sram ( mux_tree_tapbuf_size10_0_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size10_0_sram_inv ) , 
    .out ( top_grid_pin_0_ ) , .p0 ( optlc_net_143 ) ) ;
mux_tree_tapbuf_size10_mem_14 mem_bottom_ipin_0 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( ccff_head ) ,
    .ccff_tail ( { ropt_net_181 } ) ,
    .mem_out ( mux_tree_tapbuf_size10_0_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size10_0_sram_inv ) ) ;
sky130_fd_sc_hd__conb_1 optlc_143 ( .LO ( SYNOPSYS_UNCONNECTED_1 ) , 
    .HI ( optlc_net_143 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_722 ( .A ( ropt_net_144 ) , 
    .X ( ropt_net_196 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_723 ( .A ( chanx_right_in[4] ) , 
    .X ( ropt_net_207 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_724 ( .A ( chanx_left_in[13] ) , 
    .X ( ropt_net_215 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_725 ( .A ( ropt_net_147 ) , 
    .X ( chanx_left_out[8] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_762 ( .A ( ropt_net_184 ) , 
    .X ( chanx_left_out[9] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_726 ( .A ( ropt_net_148 ) , 
    .X ( ropt_net_192 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_727 ( .A ( ropt_net_149 ) , 
    .X ( ropt_net_191 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_728 ( .A ( chanx_left_in[18] ) , 
    .X ( ropt_net_210 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_729 ( .A ( chanx_right_in[5] ) , 
    .X ( ropt_net_208 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_730 ( .A ( ropt_net_152 ) , 
    .X ( ropt_net_185 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_731 ( .A ( chanx_right_in[18] ) , 
    .X ( ropt_net_213 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_732 ( .A ( chanx_right_in[13] ) , 
    .X ( ropt_net_209 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_733 ( .A ( ropt_net_155 ) , 
    .X ( ropt_net_193 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_734 ( .A ( chanx_left_in[17] ) , 
    .X ( ropt_net_202 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_735 ( .A ( chanx_left_in[16] ) , 
    .X ( ropt_net_201 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_736 ( .A ( chanx_right_in[14] ) , 
    .X ( ropt_net_200 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_737 ( .A ( chanx_left_in[14] ) , 
    .X ( ropt_net_204 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_738 ( .A ( chanx_left_in[6] ) , 
    .X ( ropt_net_214 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_739 ( .A ( chanx_right_in[17] ) , 
    .X ( ropt_net_203 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_740 ( .A ( chanx_left_in[19] ) , 
    .X ( ropt_net_212 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_741 ( .A ( chanx_right_in[15] ) , 
    .X ( ropt_net_206 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_763 ( .A ( ropt_net_185 ) , 
    .X ( chanx_left_out[6] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_742 ( .A ( chanx_left_in[12] ) , 
    .X ( ropt_net_216 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_743 ( .A ( chanx_right_in[16] ) , 
    .X ( ropt_net_205 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_744 ( .A ( chanx_right_in[10] ) , 
    .X ( ropt_net_188 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_745 ( .A ( ropt_net_167 ) , 
    .X ( ropt_net_184 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_746 ( .A ( chanx_left_in[5] ) , 
    .X ( ropt_net_211 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_747 ( .A ( chanx_right_in[0] ) , 
    .X ( ropt_net_187 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_748 ( .A ( ropt_net_170 ) , 
    .X ( chanx_right_out[7] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_749 ( .A ( ropt_net_171 ) , 
    .X ( ropt_net_195 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_750 ( .A ( ropt_net_172 ) , 
    .X ( ropt_net_197 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_751 ( .A ( ropt_net_173 ) , 
    .X ( ropt_net_190 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_752 ( .A ( ropt_net_174 ) , 
    .X ( ropt_net_189 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_753 ( .A ( ropt_net_175 ) , 
    .X ( ropt_net_186 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_754 ( .A ( ropt_net_176 ) , 
    .X ( chanx_right_out[11] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_755 ( .A ( ropt_net_177 ) , 
    .X ( ropt_net_194 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_756 ( .A ( ropt_net_178 ) , 
    .X ( chanx_right_out[15] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_757 ( .A ( ropt_net_179 ) , 
    .X ( ropt_net_198 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_758 ( .A ( ropt_net_180 ) , 
    .X ( chanx_right_out[9] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_764 ( .A ( ropt_net_186 ) , 
    .X ( chanx_left_out[1] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_759 ( .A ( ropt_net_181 ) , 
    .X ( ropt_net_199 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_765 ( .A ( ropt_net_187 ) , 
    .X ( chanx_left_out[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_44 ( .A ( chanx_left_in[8] ) , 
    .X ( BUF_net_44 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_760 ( .A ( ropt_net_182 ) , 
    .X ( chanx_right_out[0] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_761 ( .A ( ropt_net_183 ) , 
    .X ( chanx_right_out[4] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_766 ( .A ( ropt_net_188 ) , 
    .X ( chanx_left_out[10] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_767 ( .A ( ropt_net_189 ) , 
    .X ( chanx_left_out[11] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_768 ( .A ( ropt_net_190 ) , 
    .X ( chanx_left_out[7] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_769 ( .A ( ropt_net_191 ) , 
    .X ( chanx_left_out[3] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_770 ( .A ( ropt_net_192 ) , 
    .X ( chanx_right_out[1] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_771 ( .A ( ropt_net_193 ) , 
    .X ( chanx_left_out[12] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_772 ( .A ( ropt_net_194 ) , 
    .X ( chanx_left_out[19] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_54 ( .A ( chanx_right_in[1] ) , 
    .X ( ropt_net_175 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_773 ( .A ( ropt_net_195 ) , 
    .X ( chanx_right_out[10] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_774 ( .A ( ropt_net_196 ) , 
    .X ( chanx_left_out[2] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_775 ( .A ( ropt_net_197 ) , 
    .X ( chanx_right_out[2] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_776 ( .A ( ropt_net_198 ) , 
    .X ( chanx_right_out[3] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_777 ( .A ( ropt_net_199 ) , 
    .X ( ccff_tail[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_60 ( .A ( chanx_right_in[7] ) , 
    .X ( ropt_net_173 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_778 ( .A ( ropt_net_200 ) , 
    .X ( chanx_left_out[14] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_62 ( .A ( chanx_right_in[9] ) , 
    .X ( ropt_net_167 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_779 ( .A ( ropt_net_201 ) , 
    .X ( chanx_right_out[16] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_64 ( .A ( chanx_right_in[11] ) , 
    .X ( ropt_net_174 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_780 ( .A ( ropt_net_202 ) , 
    .X ( chanx_right_out[17] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_781 ( .A ( ropt_net_203 ) , 
    .X ( chanx_left_out[17] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_782 ( .A ( ropt_net_204 ) , 
    .X ( chanx_right_out[14] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_783 ( .A ( ropt_net_205 ) , 
    .X ( chanx_left_out[16] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_784 ( .A ( ropt_net_206 ) , 
    .X ( chanx_left_out[15] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_785 ( .A ( ropt_net_207 ) , 
    .X ( chanx_left_out[4] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_786 ( .A ( ropt_net_208 ) , 
    .X ( chanx_left_out[5] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_72 ( .A ( chanx_right_in[19] ) , 
    .X ( ropt_net_177 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_787 ( .A ( ropt_net_209 ) , 
    .X ( chanx_left_out[13] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_788 ( .A ( ropt_net_210 ) , 
    .X ( chanx_right_out[18] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_789 ( .A ( ropt_net_211 ) , 
    .X ( chanx_right_out[5] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_790 ( .A ( ropt_net_212 ) , 
    .X ( chanx_right_out[19] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_791 ( .A ( ropt_net_213 ) , 
    .X ( chanx_left_out[18] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_792 ( .A ( ropt_net_214 ) , 
    .X ( chanx_right_out[6] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_793 ( .A ( ropt_net_215 ) , 
    .X ( chanx_right_out[13] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_794 ( .A ( ropt_net_216 ) , 
    .X ( chanx_right_out[12] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_P_102 ( .A ( chanx_left_in[0] ) , 
    .X ( ropt_net_182 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_P_103 ( .A ( chanx_left_in[2] ) , 
    .X ( ropt_net_172 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_P_104 ( .A ( chanx_left_in[3] ) , 
    .X ( ropt_net_179 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_P_105 ( .A ( chanx_left_in[7] ) , 
    .X ( ropt_net_170 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_P_106 ( .A ( chanx_left_in[11] ) , 
    .X ( ropt_net_176 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_P_108 ( .A ( chanx_left_in[15] ) , 
    .X ( ropt_net_178 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_P_110 ( .A ( chanx_right_in[2] ) , 
    .X ( ropt_net_144 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_P_116 ( .A ( chanx_left_in[1] ) , 
    .X ( ropt_net_148 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_P_117 ( .A ( chanx_left_in[4] ) , 
    .X ( ropt_net_183 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 BUFT_P_119 ( .A ( BUF_net_44 ) , 
    .X ( chanx_right_out[8] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_P_120 ( .A ( chanx_left_in[9] ) , 
    .X ( ropt_net_180 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_P_121 ( .A ( chanx_left_in[10] ) , 
    .X ( ropt_net_171 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_P_129 ( .A ( chanx_right_in[3] ) , 
    .X ( ropt_net_149 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_P_132 ( .A ( chanx_right_in[6] ) , 
    .X ( ropt_net_152 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 BUFT_P_133 ( .A ( chanx_right_in[8] ) , 
    .X ( ropt_net_147 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_P_136 ( .A ( chanx_right_in[12] ) , 
    .X ( ropt_net_155 ) ) ;
endmodule


module mux_tree_tapbuf_size8_mem_3_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_16__55 ( .A ( mem_out[3] ) , 
    .X ( net_net_72 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_71 ( .A ( net_net_72 ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size8_mem_2_2 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_15__54 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size8_mem_1_3 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_14__53 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size8_mem_0_3 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_13__52 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size8_mem_8 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_12__51 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size8_mem_6_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_11__50 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size8_mem_5_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_10__49 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size8_mem_4_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_9__48 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_41 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size8_3_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:7] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;

const1_41 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( in[2] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[4] ) , .A1 ( in[3] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[6] ) , .A1 ( in[5] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
endmodule


module const1_14_10 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size8_2_2 ( in , sram , sram_inv , out , p0 ) ;
input  [0:7] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;

const1_14_10 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( in[2] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[4] ) , .A1 ( in[3] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[6] ) , .A1 ( in[5] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
endmodule


module const1_13_10 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size8_1_3 ( in , sram , sram_inv , out , p0 ) ;
input  [0:7] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;

const1_13_10 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( in[2] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[4] ) , .A1 ( in[3] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[6] ) , .A1 ( in[5] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
endmodule


module const1_12_10 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size8_0_3 ( in , sram , sram_inv , out , p0 ) ;
input  [0:7] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;

const1_12_10 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( in[2] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[4] ) , .A1 ( in[3] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[6] ) , .A1 ( in[5] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
endmodule


module const1_11_10 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size8_8 ( in , sram , sram_inv , out , p0 ) ;
input  [0:7] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;

const1_11_10 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( in[2] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[4] ) , .A1 ( in[3] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[6] ) , .A1 ( in[5] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_8 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[3] ) , .X ( out[0] ) ) ;
endmodule


module const1_10_10 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size8_6_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:7] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;

const1_10_10 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( in[2] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[4] ) , .A1 ( in[3] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[6] ) , .A1 ( in[5] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
endmodule


module const1_9_10 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size8_5_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:7] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;

const1_9_10 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( in[2] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[4] ) , .A1 ( in[3] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[6] ) , .A1 ( in[5] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
endmodule


module const1_8_10 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size8_4_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:7] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;

const1_8_10 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( in[2] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[4] ) , .A1 ( in[3] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[6] ) , .A1 ( in[5] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
endmodule


module mux_tree_tapbuf_size10_mem_3_2 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_8__47 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size10_mem_2_2 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_7__46 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size10_mem_13 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_6__45 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size10_mem_6_2 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_5__44 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size10_mem_5_2 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_4__43 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size10_mem_4_2 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_3__42 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size10_mem_1_2 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_2__41 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size10_mem_0_3 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_1__40 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_7_10 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size10_3_2 ( in , sram , sram_inv , out , p0 ) ;
input  [0:9] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

const1_7_10 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[6] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[8] ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[9] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
endmodule


module const1_6_11 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size10_2_2 ( in , sram , sram_inv , out , p0 ) ;
input  [0:9] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

const1_6_11 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[6] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[8] ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[9] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
endmodule


module const1_5_11 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size10_13 ( in , sram , sram_inv , out , p0 ) ;
input  [0:9] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

const1_5_11 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[6] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[8] ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[9] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
endmodule


module const1_4_11 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size10_6_2 ( in , sram , sram_inv , out , p0 ) ;
input  [0:9] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

const1_4_11 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[6] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[8] ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[9] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
endmodule


module const1_3_11 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size10_5_2 ( in , sram , sram_inv , out , p0 ) ;
input  [0:9] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

const1_3_11 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[6] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[8] ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[9] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
endmodule


module const1_2_11 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size10_4_2 ( in , sram , sram_inv , out , p0 ) ;
input  [0:9] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

const1_2_11 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[6] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[8] ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[9] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
endmodule


module const1_1_11 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size10_1_2 ( in , sram , sram_inv , out , p0 ) ;
input  [0:9] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

const1_1_11 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[6] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[8] ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[9] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
endmodule


module const1_0_11 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size10_0_3 ( in , sram , sram_inv , out , p0 ) ;
input  [0:9] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

const1_0_11 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[6] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[8] ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[9] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
endmodule


module cbx_1__1_ ( prog_clk , chanx_left_in , chanx_right_in , ccff_head , 
    chanx_left_out , chanx_right_out , top_grid_pin_16_ , top_grid_pin_17_ , 
    top_grid_pin_18_ , top_grid_pin_19_ , top_grid_pin_20_ , 
    top_grid_pin_21_ , top_grid_pin_22_ , top_grid_pin_23_ , 
    top_grid_pin_24_ , top_grid_pin_25_ , top_grid_pin_26_ , 
    top_grid_pin_27_ , top_grid_pin_28_ , top_grid_pin_29_ , 
    top_grid_pin_30_ , top_grid_pin_31_ , ccff_tail ) ;
input  [0:0] prog_clk ;
input  [0:19] chanx_left_in ;
input  [0:19] chanx_right_in ;
input  [0:0] ccff_head ;
output [0:19] chanx_left_out ;
output [0:19] chanx_right_out ;
output [0:0] top_grid_pin_16_ ;
output [0:0] top_grid_pin_17_ ;
output [0:0] top_grid_pin_18_ ;
output [0:0] top_grid_pin_19_ ;
output [0:0] top_grid_pin_20_ ;
output [0:0] top_grid_pin_21_ ;
output [0:0] top_grid_pin_22_ ;
output [0:0] top_grid_pin_23_ ;
output [0:0] top_grid_pin_24_ ;
output [0:0] top_grid_pin_25_ ;
output [0:0] top_grid_pin_26_ ;
output [0:0] top_grid_pin_27_ ;
output [0:0] top_grid_pin_28_ ;
output [0:0] top_grid_pin_29_ ;
output [0:0] top_grid_pin_30_ ;
output [0:0] top_grid_pin_31_ ;
output [0:0] ccff_tail ;

wire [0:3] mux_tree_tapbuf_size10_0_sram ;
wire [0:3] mux_tree_tapbuf_size10_0_sram_inv ;
wire [0:3] mux_tree_tapbuf_size10_1_sram ;
wire [0:3] mux_tree_tapbuf_size10_1_sram_inv ;
wire [0:3] mux_tree_tapbuf_size10_2_sram ;
wire [0:3] mux_tree_tapbuf_size10_2_sram_inv ;
wire [0:3] mux_tree_tapbuf_size10_3_sram ;
wire [0:3] mux_tree_tapbuf_size10_3_sram_inv ;
wire [0:3] mux_tree_tapbuf_size10_4_sram ;
wire [0:3] mux_tree_tapbuf_size10_4_sram_inv ;
wire [0:3] mux_tree_tapbuf_size10_5_sram ;
wire [0:3] mux_tree_tapbuf_size10_5_sram_inv ;
wire [0:3] mux_tree_tapbuf_size10_6_sram ;
wire [0:3] mux_tree_tapbuf_size10_6_sram_inv ;
wire [0:3] mux_tree_tapbuf_size10_7_sram ;
wire [0:3] mux_tree_tapbuf_size10_7_sram_inv ;
wire [0:0] mux_tree_tapbuf_size10_mem_0_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size10_mem_1_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size10_mem_2_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size10_mem_3_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size10_mem_4_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size10_mem_5_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size10_mem_6_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size10_mem_7_ccff_tail ;
wire [0:3] mux_tree_tapbuf_size8_0_sram ;
wire [0:3] mux_tree_tapbuf_size8_0_sram_inv ;
wire [0:3] mux_tree_tapbuf_size8_1_sram ;
wire [0:3] mux_tree_tapbuf_size8_1_sram_inv ;
wire [0:3] mux_tree_tapbuf_size8_2_sram ;
wire [0:3] mux_tree_tapbuf_size8_2_sram_inv ;
wire [0:3] mux_tree_tapbuf_size8_3_sram ;
wire [0:3] mux_tree_tapbuf_size8_3_sram_inv ;
wire [0:3] mux_tree_tapbuf_size8_4_sram ;
wire [0:3] mux_tree_tapbuf_size8_4_sram_inv ;
wire [0:3] mux_tree_tapbuf_size8_5_sram ;
wire [0:3] mux_tree_tapbuf_size8_5_sram_inv ;
wire [0:3] mux_tree_tapbuf_size8_6_sram ;
wire [0:3] mux_tree_tapbuf_size8_6_sram_inv ;
wire [0:3] mux_tree_tapbuf_size8_7_sram ;
wire [0:3] mux_tree_tapbuf_size8_7_sram_inv ;
wire [0:0] mux_tree_tapbuf_size8_mem_0_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size8_mem_1_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size8_mem_2_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size8_mem_3_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size8_mem_4_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size8_mem_5_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size8_mem_6_ccff_tail ;

mux_tree_tapbuf_size10_0_3 mux_bottom_ipin_0 (
    .in ( { chanx_left_in[0] , chanx_right_in[0] , chanx_left_in[2] , 
        chanx_right_in[2] , chanx_left_in[4] , chanx_right_in[4] , 
        chanx_left_in[10] , chanx_right_in[10] , chanx_left_in[16] , 
        chanx_right_in[16] } ) ,
    .sram ( mux_tree_tapbuf_size10_0_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size10_0_sram_inv ) , 
    .out ( top_grid_pin_16_ ) , .p0 ( optlc_net_94 ) ) ;
mux_tree_tapbuf_size10_1_2 mux_bottom_ipin_1 (
    .in ( { chanx_left_in[1] , chanx_right_in[1] , chanx_left_in[3] , 
        chanx_right_in[3] , chanx_left_in[5] , chanx_right_in[5] , 
        chanx_left_in[11] , chanx_right_in[11] , chanx_left_in[17] , 
        chanx_right_in[17] } ) ,
    .sram ( mux_tree_tapbuf_size10_1_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size10_1_sram_inv ) , 
    .out ( top_grid_pin_17_ ) , .p0 ( optlc_net_95 ) ) ;
mux_tree_tapbuf_size10_4_2 mux_bottom_ipin_4 (
    .in ( { chanx_left_in[0] , chanx_right_in[0] , chanx_left_in[2] , 
        chanx_right_in[2] , chanx_left_in[4] , chanx_right_in[4] , 
        chanx_left_in[8] , chanx_right_in[8] , chanx_left_in[14] , 
        chanx_right_in[14] } ) ,
    .sram ( mux_tree_tapbuf_size10_2_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size10_2_sram_inv ) , 
    .out ( top_grid_pin_20_ ) , .p0 ( optlc_net_94 ) ) ;
mux_tree_tapbuf_size10_5_2 mux_bottom_ipin_5 (
    .in ( { chanx_left_in[1] , chanx_right_in[1] , chanx_left_in[3] , 
        chanx_right_in[3] , chanx_left_in[5] , chanx_right_in[5] , 
        chanx_left_in[9] , chanx_right_in[9] , chanx_left_in[15] , 
        chanx_right_in[15] } ) ,
    .sram ( mux_tree_tapbuf_size10_3_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size10_3_sram_inv ) , 
    .out ( top_grid_pin_21_ ) , .p0 ( optlc_net_94 ) ) ;
mux_tree_tapbuf_size10_6_2 mux_bottom_ipin_8 (
    .in ( { chanx_left_in[0] , chanx_right_in[0] , chanx_left_in[2] , 
        chanx_right_in[2] , chanx_left_in[8] , chanx_right_in[8] , 
        chanx_left_in[12] , chanx_right_in[12] , chanx_left_in[18] , 
        chanx_right_in[18] } ) ,
    .sram ( mux_tree_tapbuf_size10_4_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size10_4_sram_inv ) , 
    .out ( top_grid_pin_24_ ) , .p0 ( optlc_net_94 ) ) ;
mux_tree_tapbuf_size10_13 mux_bottom_ipin_9 (
    .in ( { chanx_left_in[1] , chanx_right_in[1] , chanx_left_in[3] , 
        chanx_right_in[3] , chanx_left_in[9] , chanx_right_in[9] , 
        chanx_left_in[13] , chanx_right_in[13] , chanx_left_in[19] , 
        chanx_right_in[19] } ) ,
    .sram ( mux_tree_tapbuf_size10_5_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size10_5_sram_inv ) , 
    .out ( top_grid_pin_25_ ) , .p0 ( optlc_net_95 ) ) ;
mux_tree_tapbuf_size10_2_2 mux_bottom_ipin_12 (
    .in ( { chanx_left_in[0] , chanx_right_in[0] , chanx_left_in[2] , 
        chanx_right_in[2] , chanx_left_in[6] , chanx_right_in[6] , 
        chanx_left_in[12] , chanx_right_in[12] , chanx_left_in[16] , 
        chanx_right_in[16] } ) ,
    .sram ( mux_tree_tapbuf_size10_6_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size10_6_sram_inv ) , 
    .out ( top_grid_pin_28_ ) , .p0 ( optlc_net_94 ) ) ;
mux_tree_tapbuf_size10_3_2 mux_bottom_ipin_13 (
    .in ( { chanx_left_in[1] , chanx_right_in[1] , chanx_left_in[3] , 
        chanx_right_in[3] , chanx_left_in[7] , chanx_right_in[7] , 
        chanx_left_in[13] , chanx_right_in[13] , chanx_left_in[17] , 
        chanx_right_in[17] } ) ,
    .sram ( mux_tree_tapbuf_size10_7_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size10_7_sram_inv ) , 
    .out ( top_grid_pin_29_ ) , .p0 ( optlc_net_95 ) ) ;
mux_tree_tapbuf_size10_mem_0_3 mem_bottom_ipin_0 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( ccff_head ) , 
    .ccff_tail ( mux_tree_tapbuf_size10_mem_0_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size10_0_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size10_0_sram_inv ) ) ;
mux_tree_tapbuf_size10_mem_1_2 mem_bottom_ipin_1 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size10_mem_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size10_mem_1_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size10_1_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size10_1_sram_inv ) ) ;
mux_tree_tapbuf_size10_mem_4_2 mem_bottom_ipin_4 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size8_mem_1_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size10_mem_2_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size10_2_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size10_2_sram_inv ) ) ;
mux_tree_tapbuf_size10_mem_5_2 mem_bottom_ipin_5 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size10_mem_2_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size10_mem_3_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size10_3_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size10_3_sram_inv ) ) ;
mux_tree_tapbuf_size10_mem_6_2 mem_bottom_ipin_8 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size8_mem_3_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size10_mem_4_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size10_4_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size10_4_sram_inv ) ) ;
mux_tree_tapbuf_size10_mem_13 mem_bottom_ipin_9 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size10_mem_4_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size10_mem_5_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size10_5_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size10_5_sram_inv ) ) ;
mux_tree_tapbuf_size10_mem_2_2 mem_bottom_ipin_12 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size8_mem_5_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size10_mem_6_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size10_6_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size10_6_sram_inv ) ) ;
mux_tree_tapbuf_size10_mem_3_2 mem_bottom_ipin_13 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size10_mem_6_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size10_mem_7_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size10_7_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size10_7_sram_inv ) ) ;
mux_tree_tapbuf_size8_4_1 mux_bottom_ipin_2 (
    .in ( { chanx_left_in[0] , chanx_right_in[0] , chanx_left_in[2] , 
        chanx_right_in[2] , chanx_left_in[6] , chanx_right_in[6] , 
        chanx_left_in[14] , chanx_right_in[14] } ) ,
    .sram ( mux_tree_tapbuf_size8_0_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size8_0_sram_inv ) , 
    .out ( top_grid_pin_18_ ) , .p0 ( optlc_net_94 ) ) ;
mux_tree_tapbuf_size8_5_1 mux_bottom_ipin_3 (
    .in ( { chanx_left_in[1] , chanx_right_in[1] , chanx_left_in[3] , 
        chanx_right_in[3] , chanx_left_in[7] , chanx_right_in[7] , 
        chanx_left_in[15] , chanx_right_in[15] } ) ,
    .sram ( mux_tree_tapbuf_size8_1_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size8_1_sram_inv ) , 
    .out ( top_grid_pin_19_ ) , .p0 ( optlc_net_95 ) ) ;
mux_tree_tapbuf_size8_6_1 mux_bottom_ipin_6 (
    .in ( { chanx_left_in[0] , chanx_right_in[0] , chanx_left_in[2] , 
        chanx_right_in[2] , chanx_left_in[10] , chanx_right_in[10] , 
        chanx_left_in[18] , chanx_right_in[18] } ) ,
    .sram ( mux_tree_tapbuf_size8_2_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size8_2_sram_inv ) , 
    .out ( top_grid_pin_22_ ) , .p0 ( optlc_net_95 ) ) ;
mux_tree_tapbuf_size8_8 mux_bottom_ipin_7 (
    .in ( { chanx_left_in[1] , chanx_right_in[1] , chanx_left_in[3] , 
        chanx_right_in[3] , chanx_left_in[11] , chanx_right_in[11] , 
        chanx_left_in[19] , chanx_right_in[19] } ) ,
    .sram ( mux_tree_tapbuf_size8_3_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size8_3_sram_inv ) , 
    .out ( top_grid_pin_23_ ) , .p0 ( optlc_net_95 ) ) ;
mux_tree_tapbuf_size8_0_3 mux_bottom_ipin_10 (
    .in ( { chanx_left_in[0] , chanx_right_in[0] , chanx_left_in[2] , 
        chanx_right_in[2] , chanx_left_in[6] , chanx_right_in[6] , 
        chanx_left_in[14] , chanx_right_in[14] } ) ,
    .sram ( mux_tree_tapbuf_size8_4_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size8_4_sram_inv ) , 
    .out ( top_grid_pin_26_ ) , .p0 ( optlc_net_94 ) ) ;
mux_tree_tapbuf_size8_1_3 mux_bottom_ipin_11 (
    .in ( { chanx_left_in[1] , chanx_right_in[1] , chanx_left_in[3] , 
        chanx_right_in[3] , chanx_left_in[7] , chanx_right_in[7] , 
        chanx_left_in[15] , chanx_right_in[15] } ) ,
    .sram ( mux_tree_tapbuf_size8_5_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size8_5_sram_inv ) , 
    .out ( top_grid_pin_27_ ) , .p0 ( optlc_net_94 ) ) ;
mux_tree_tapbuf_size8_2_2 mux_bottom_ipin_14 (
    .in ( { chanx_left_in[0] , chanx_right_in[0] , chanx_left_in[2] , 
        chanx_right_in[2] , chanx_left_in[10] , chanx_right_in[10] , 
        chanx_left_in[18] , chanx_right_in[18] } ) ,
    .sram ( mux_tree_tapbuf_size8_6_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size8_6_sram_inv ) , 
    .out ( top_grid_pin_30_ ) , .p0 ( optlc_net_95 ) ) ;
mux_tree_tapbuf_size8_3_1 mux_bottom_ipin_15 (
    .in ( { chanx_left_in[1] , chanx_right_in[1] , chanx_left_in[3] , 
        chanx_right_in[3] , chanx_left_in[11] , chanx_right_in[11] , 
        chanx_left_in[19] , chanx_right_in[19] } ) ,
    .sram ( mux_tree_tapbuf_size8_7_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size8_7_sram_inv ) , 
    .out ( top_grid_pin_31_ ) , .p0 ( optlc_net_95 ) ) ;
mux_tree_tapbuf_size8_mem_4_1 mem_bottom_ipin_2 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size10_mem_1_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size8_mem_0_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size8_0_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size8_0_sram_inv ) ) ;
mux_tree_tapbuf_size8_mem_5_1 mem_bottom_ipin_3 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size8_mem_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size8_mem_1_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size8_1_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size8_1_sram_inv ) ) ;
mux_tree_tapbuf_size8_mem_6_1 mem_bottom_ipin_6 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size10_mem_3_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size8_mem_2_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size8_2_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size8_2_sram_inv ) ) ;
mux_tree_tapbuf_size8_mem_8 mem_bottom_ipin_7 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size8_mem_2_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size8_mem_3_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size8_3_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size8_3_sram_inv ) ) ;
mux_tree_tapbuf_size8_mem_0_3 mem_bottom_ipin_10 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size10_mem_5_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size8_mem_4_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size8_4_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size8_4_sram_inv ) ) ;
mux_tree_tapbuf_size8_mem_1_3 mem_bottom_ipin_11 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size8_mem_4_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size8_mem_5_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size8_5_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size8_5_sram_inv ) ) ;
mux_tree_tapbuf_size8_mem_2_2 mem_bottom_ipin_14 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size10_mem_7_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size8_mem_6_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size8_6_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size8_6_sram_inv ) ) ;
mux_tree_tapbuf_size8_mem_3_1 mem_bottom_ipin_15 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size8_mem_6_ccff_tail ) ,
    .ccff_tail ( { ropt_net_97 } ) ,
    .mem_out ( mux_tree_tapbuf_size8_7_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size8_7_sram_inv ) ) ;
sky130_fd_sc_hd__conb_1 optlc_92 ( .LO ( SYNOPSYS_UNCONNECTED_1 ) , 
    .HI ( optlc_net_94 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_2__1 ( .A ( chanx_left_in[1] ) , 
    .X ( chanx_right_out[1] ) ) ;
sky130_fd_sc_hd__conb_1 optlc_94 ( .LO ( SYNOPSYS_UNCONNECTED_2 ) , 
    .HI ( optlc_net_95 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_4__3 ( .A ( chanx_left_in[3] ) , 
    .X ( chanx_right_out[3] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_684 ( .A ( ropt_net_105 ) , 
    .X ( chanx_right_out[8] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_6__5 ( .A ( chanx_left_in[5] ) , 
    .X ( chanx_right_out[5] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_7__6 ( .A ( chanx_left_in[6] ) , 
    .X ( chanx_right_out[6] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_8__7 ( .A ( chanx_left_in[7] ) , 
    .X ( chanx_right_out[7] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_673 ( .A ( chanx_left_in[15] ) , 
    .X ( chanx_right_out[15] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_685 ( .A ( ropt_net_106 ) , 
    .X ( chanx_right_out[12] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_11__10 ( .A ( chanx_left_in[10] ) , 
    .X ( chanx_right_out[10] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_12__11 ( .A ( chanx_left_in[11] ) , 
    .X ( chanx_right_out[11] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_686 ( .A ( ropt_net_107 ) , 
    .X ( chanx_left_out[13] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_14__13 ( .A ( chanx_left_in[13] ) , 
    .X ( chanx_right_out[13] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_675 ( .A ( ropt_net_97 ) , 
    .X ( ropt_net_108 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_687 ( .A ( ropt_net_108 ) , 
    .X ( ccff_tail[0] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_17__16 ( .A ( chanx_left_in[16] ) , 
    .X ( chanx_right_out[16] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_676 ( .A ( ropt_net_98 ) , 
    .X ( chanx_right_out[4] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_678 ( .A ( chanx_right_in[4] ) , 
    .X ( chanx_left_out[4] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_679 ( .A ( chanx_left_in[12] ) , 
    .X ( ropt_net_106 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_21__20 ( .A ( chanx_right_in[0] ) , 
    .X ( chanx_left_out[0] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_22__21 ( .A ( chanx_right_in[1] ) , 
    .X ( chanx_left_out[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd1_1 FTB_23__22 ( .A ( chanx_right_in[2] ) , 
    .X ( chanx_left_out[2] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_680 ( .A ( chanx_right_in[16] ) , 
    .X ( chanx_left_out[16] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_26__25 ( .A ( chanx_right_in[5] ) , 
    .X ( aps_rename_2_ ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_681 ( .A ( ropt_net_102 ) , 
    .X ( chanx_left_out[12] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_28__27 ( .A ( chanx_right_in[7] ) , 
    .X ( chanx_left_out[7] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_682 ( .A ( ropt_net_103 ) , 
    .X ( chanx_left_out[18] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_30__29 ( .A ( chanx_right_in[9] ) , 
    .X ( chanx_left_out[9] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_31__30 ( .A ( chanx_right_in[10] ) , 
    .X ( ropt_net_104 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_32__31 ( .A ( chanx_right_in[11] ) , 
    .X ( aps_rename_3_ ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_683 ( .A ( ropt_net_104 ) , 
    .X ( chanx_left_out[10] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_34__33 ( .A ( chanx_right_in[13] ) , 
    .X ( ropt_net_107 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_35__34 ( .A ( chanx_right_in[14] ) , 
    .X ( chanx_left_out[14] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_36__35 ( .A ( chanx_right_in[15] ) , 
    .X ( chanx_left_out[15] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_38__37 ( .A ( chanx_right_in[17] ) , 
    .X ( chanx_left_out[17] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_39__38 ( .A ( chanx_right_in[18] ) , 
    .X ( ropt_net_103 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_40__39 ( .A ( chanx_right_in[19] ) , 
    .X ( chanx_left_out[19] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 BUFT_RR_59 ( .A ( chanx_left_in[4] ) , 
    .X ( ropt_net_98 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_RR_60 ( .A ( chanx_left_in[8] ) , 
    .X ( ropt_net_105 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_61 ( .A ( chanx_left_in[9] ) , 
    .X ( BUF_net_61 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_RR_64 ( .A ( chanx_left_in[19] ) , 
    .X ( chanx_right_out[19] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_RR_67 ( .A ( chanx_right_in[8] ) , 
    .X ( chanx_left_out[8] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 BUFT_RR_76 ( .A ( BUF_net_61 ) , 
    .X ( chanx_right_out[9] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_RR_78 ( .A ( chanx_left_in[14] ) , 
    .X ( chanx_right_out[14] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 BUFT_RR_79 ( .A ( aps_rename_3_ ) , 
    .X ( chanx_left_out[11] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_RR_80 ( .A ( chanx_right_in[12] ) , 
    .X ( ropt_net_102 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_P_82 ( .A ( chanx_left_in[0] ) , 
    .X ( chanx_right_out[0] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_P_83 ( .A ( chanx_left_in[2] ) , 
    .X ( chanx_right_out[2] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_P_84 ( .A ( chanx_left_in[17] ) , 
    .X ( chanx_right_out[17] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_P_85 ( .A ( chanx_left_in[18] ) , 
    .X ( chanx_right_out[18] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_P_86 ( .A ( chanx_right_in[3] ) , 
    .X ( chanx_left_out[3] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_P_87 ( .A ( chanx_right_in[6] ) , 
    .X ( chanx_left_out[6] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 BUFT_P_89 ( .A ( aps_rename_2_ ) , 
    .X ( chanx_left_out[5] ) ) ;
endmodule


module mux_tree_tapbuf_size8_mem_3 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_17__56 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size8_mem_2_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_16__55 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size8_mem_1_2 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_15__54 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size8_mem_0_2 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_14__53 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size8_mem_7 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_13__52 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size8_mem_6 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_12__51 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size8_mem_5 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_11__50 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size8_mem_4 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_10__49 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_40 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size8_3 ( in , sram , sram_inv , out , p0 ) ;
input  [0:7] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;

const1_40 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( in[2] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[4] ) , .A1 ( in[3] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[6] ) , .A1 ( in[5] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
endmodule


module const1_15_9 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size8_2_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:7] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;

const1_15_9 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( in[2] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[4] ) , .A1 ( in[3] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[6] ) , .A1 ( in[5] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
endmodule


module const1_14_9 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size8_1_2 ( in , sram , sram_inv , out , p0 ) ;
input  [0:7] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;

const1_14_9 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( in[2] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[4] ) , .A1 ( in[3] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[6] ) , .A1 ( in[5] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
endmodule


module const1_13_9 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size8_0_2 ( in , sram , sram_inv , out , p0 ) ;
input  [0:7] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;

const1_13_9 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( in[2] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[4] ) , .A1 ( in[3] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[6] ) , .A1 ( in[5] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
endmodule


module const1_12_9 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size8_7 ( in , sram , sram_inv , out , p0 ) ;
input  [0:7] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;

const1_12_9 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( in[2] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[4] ) , .A1 ( in[3] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[6] ) , .A1 ( in[5] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_4 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[3] ) , .X ( out[0] ) ) ;
endmodule


module const1_11_9 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size8_6 ( in , sram , sram_inv , out , p0 ) ;
input  [0:7] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;

const1_11_9 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( in[2] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[4] ) , .A1 ( in[3] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[6] ) , .A1 ( in[5] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
endmodule


module const1_10_9 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size8_5 ( in , sram , sram_inv , out , p0 ) ;
input  [0:7] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;

const1_10_9 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( in[2] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[4] ) , .A1 ( in[3] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[6] ) , .A1 ( in[5] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_4 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[3] ) , .X ( out[0] ) ) ;
endmodule


module const1_9_9 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size8_4 ( in , sram , sram_inv , out , p0 ) ;
input  [0:7] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;

const1_9_9 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( in[2] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[4] ) , .A1 ( in[3] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[6] ) , .A1 ( in[5] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
endmodule


module mux_tree_tapbuf_size10_mem_12 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd1_1 FTB_9__48 ( .A ( mem_out[3] ) , 
    .X ( net_net_69 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_P_86 ( .A ( net_net_69 ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size10_mem_3_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_8__47 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size10_mem_2_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_7__46 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size10_mem_7_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_6__45 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size10_mem_6_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_5__44 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size10_mem_5_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_4__43 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size10_mem_4_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_3__42 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size10_mem_1_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_2__41 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size10_mem_0_2 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_1__40 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_8_9 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size10_12 ( in , sram , sram_inv , out , p0 ) ;
input  [0:9] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

const1_8_9 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[6] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[8] ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[9] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
endmodule


module const1_7_9 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size10_3_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:9] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

const1_7_9 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[6] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[8] ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[9] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
endmodule


module const1_6_10 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size10_2_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:9] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

const1_6_10 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[6] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[8] ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[9] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
endmodule


module const1_5_10 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size10_7_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:9] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

const1_5_10 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[6] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[8] ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[9] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
endmodule


module const1_4_10 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size10_6_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:9] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

const1_4_10 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[6] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[8] ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[9] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
endmodule


module const1_3_10 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size10_5_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:9] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

const1_3_10 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[6] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[8] ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[9] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
endmodule


module const1_2_10 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size10_4_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:9] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

const1_2_10 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[6] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[8] ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[9] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
endmodule


module const1_1_10 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size10_1_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:9] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

const1_1_10 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[6] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[8] ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[9] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
endmodule


module const1_0_10 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size10_0_2 ( in , sram , sram_inv , out , p0 ) ;
input  [0:9] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

const1_0_10 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[6] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[8] ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[9] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
endmodule


module cbx_1__0_ ( prog_clk , chanx_left_in , chanx_right_in , ccff_head , 
    chanx_left_out , chanx_right_out , top_grid_pin_16_ , top_grid_pin_17_ , 
    top_grid_pin_18_ , top_grid_pin_19_ , top_grid_pin_20_ , 
    top_grid_pin_21_ , top_grid_pin_22_ , top_grid_pin_23_ , 
    top_grid_pin_24_ , top_grid_pin_25_ , top_grid_pin_26_ , 
    top_grid_pin_27_ , top_grid_pin_28_ , top_grid_pin_29_ , 
    top_grid_pin_30_ , top_grid_pin_31_ , bottom_grid_pin_0_ , ccff_tail ) ;
input  [0:0] prog_clk ;
input  [0:19] chanx_left_in ;
input  [0:19] chanx_right_in ;
input  [0:0] ccff_head ;
output [0:19] chanx_left_out ;
output [0:19] chanx_right_out ;
output [0:0] top_grid_pin_16_ ;
output [0:0] top_grid_pin_17_ ;
output [0:0] top_grid_pin_18_ ;
output [0:0] top_grid_pin_19_ ;
output [0:0] top_grid_pin_20_ ;
output [0:0] top_grid_pin_21_ ;
output [0:0] top_grid_pin_22_ ;
output [0:0] top_grid_pin_23_ ;
output [0:0] top_grid_pin_24_ ;
output [0:0] top_grid_pin_25_ ;
output [0:0] top_grid_pin_26_ ;
output [0:0] top_grid_pin_27_ ;
output [0:0] top_grid_pin_28_ ;
output [0:0] top_grid_pin_29_ ;
output [0:0] top_grid_pin_30_ ;
output [0:0] top_grid_pin_31_ ;
output [0:0] bottom_grid_pin_0_ ;
output [0:0] ccff_tail ;

wire [0:3] mux_tree_tapbuf_size10_0_sram ;
wire [0:3] mux_tree_tapbuf_size10_0_sram_inv ;
wire [0:3] mux_tree_tapbuf_size10_1_sram ;
wire [0:3] mux_tree_tapbuf_size10_1_sram_inv ;
wire [0:3] mux_tree_tapbuf_size10_2_sram ;
wire [0:3] mux_tree_tapbuf_size10_2_sram_inv ;
wire [0:3] mux_tree_tapbuf_size10_3_sram ;
wire [0:3] mux_tree_tapbuf_size10_3_sram_inv ;
wire [0:3] mux_tree_tapbuf_size10_4_sram ;
wire [0:3] mux_tree_tapbuf_size10_4_sram_inv ;
wire [0:3] mux_tree_tapbuf_size10_5_sram ;
wire [0:3] mux_tree_tapbuf_size10_5_sram_inv ;
wire [0:3] mux_tree_tapbuf_size10_6_sram ;
wire [0:3] mux_tree_tapbuf_size10_6_sram_inv ;
wire [0:3] mux_tree_tapbuf_size10_7_sram ;
wire [0:3] mux_tree_tapbuf_size10_7_sram_inv ;
wire [0:3] mux_tree_tapbuf_size10_8_sram ;
wire [0:3] mux_tree_tapbuf_size10_8_sram_inv ;
wire [0:0] mux_tree_tapbuf_size10_mem_0_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size10_mem_1_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size10_mem_2_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size10_mem_3_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size10_mem_4_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size10_mem_5_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size10_mem_6_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size10_mem_7_ccff_tail ;
wire [0:3] mux_tree_tapbuf_size8_0_sram ;
wire [0:3] mux_tree_tapbuf_size8_0_sram_inv ;
wire [0:3] mux_tree_tapbuf_size8_1_sram ;
wire [0:3] mux_tree_tapbuf_size8_1_sram_inv ;
wire [0:3] mux_tree_tapbuf_size8_2_sram ;
wire [0:3] mux_tree_tapbuf_size8_2_sram_inv ;
wire [0:3] mux_tree_tapbuf_size8_3_sram ;
wire [0:3] mux_tree_tapbuf_size8_3_sram_inv ;
wire [0:3] mux_tree_tapbuf_size8_4_sram ;
wire [0:3] mux_tree_tapbuf_size8_4_sram_inv ;
wire [0:3] mux_tree_tapbuf_size8_5_sram ;
wire [0:3] mux_tree_tapbuf_size8_5_sram_inv ;
wire [0:3] mux_tree_tapbuf_size8_6_sram ;
wire [0:3] mux_tree_tapbuf_size8_6_sram_inv ;
wire [0:3] mux_tree_tapbuf_size8_7_sram ;
wire [0:3] mux_tree_tapbuf_size8_7_sram_inv ;
wire [0:0] mux_tree_tapbuf_size8_mem_0_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size8_mem_1_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size8_mem_2_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size8_mem_3_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size8_mem_4_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size8_mem_5_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size8_mem_6_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size8_mem_7_ccff_tail ;

mux_tree_tapbuf_size10_0_2 mux_bottom_ipin_0 (
    .in ( { chanx_left_in[0] , chanx_right_in[0] , chanx_left_in[2] , 
        chanx_right_in[2] , chanx_left_in[4] , chanx_right_in[4] , 
        chanx_left_in[10] , chanx_right_in[10] , chanx_left_in[16] , 
        chanx_right_in[16] } ) ,
    .sram ( mux_tree_tapbuf_size10_0_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size10_0_sram_inv ) , 
    .out ( top_grid_pin_16_ ) , .p0 ( optlc_net_90 ) ) ;
mux_tree_tapbuf_size10_1_1 mux_bottom_ipin_1 (
    .in ( { chanx_left_in[1] , chanx_right_in[1] , chanx_left_in[3] , 
        chanx_right_in[3] , chanx_left_in[5] , chanx_right_in[5] , 
        chanx_left_in[11] , chanx_right_in[11] , chanx_left_in[17] , 
        chanx_right_in[17] } ) ,
    .sram ( mux_tree_tapbuf_size10_1_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size10_1_sram_inv ) , 
    .out ( top_grid_pin_17_ ) , .p0 ( optlc_net_91 ) ) ;
mux_tree_tapbuf_size10_4_1 mux_bottom_ipin_4 (
    .in ( { chanx_left_in[0] , chanx_right_in[0] , chanx_left_in[2] , 
        chanx_right_in[2] , chanx_left_in[4] , chanx_right_in[4] , 
        chanx_left_in[8] , chanx_right_in[8] , chanx_left_in[14] , 
        chanx_right_in[14] } ) ,
    .sram ( mux_tree_tapbuf_size10_2_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size10_2_sram_inv ) , 
    .out ( top_grid_pin_20_ ) , .p0 ( optlc_net_91 ) ) ;
mux_tree_tapbuf_size10_5_1 mux_bottom_ipin_5 (
    .in ( { chanx_left_in[1] , chanx_right_in[1] , chanx_left_in[3] , 
        chanx_right_in[3] , chanx_left_in[5] , chanx_right_in[5] , 
        chanx_left_in[9] , chanx_right_in[9] , chanx_left_in[15] , 
        chanx_right_in[15] } ) ,
    .sram ( mux_tree_tapbuf_size10_3_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size10_3_sram_inv ) , 
    .out ( top_grid_pin_21_ ) , .p0 ( optlc_net_91 ) ) ;
mux_tree_tapbuf_size10_6_1 mux_bottom_ipin_8 (
    .in ( { chanx_left_in[0] , chanx_right_in[0] , chanx_left_in[2] , 
        chanx_right_in[2] , chanx_left_in[8] , chanx_right_in[8] , 
        chanx_left_in[12] , chanx_right_in[12] , chanx_left_in[18] , 
        chanx_right_in[18] } ) ,
    .sram ( mux_tree_tapbuf_size10_4_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size10_4_sram_inv ) , 
    .out ( top_grid_pin_24_ ) , .p0 ( optlc_net_91 ) ) ;
mux_tree_tapbuf_size10_7_1 mux_bottom_ipin_9 (
    .in ( { chanx_left_in[1] , chanx_right_in[1] , chanx_left_in[3] , 
        chanx_right_in[3] , chanx_left_in[9] , chanx_right_in[9] , 
        chanx_left_in[13] , chanx_right_in[13] , chanx_left_in[19] , 
        chanx_right_in[19] } ) ,
    .sram ( mux_tree_tapbuf_size10_5_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size10_5_sram_inv ) , 
    .out ( top_grid_pin_25_ ) , .p0 ( optlc_net_91 ) ) ;
mux_tree_tapbuf_size10_2_1 mux_bottom_ipin_12 (
    .in ( { chanx_left_in[0] , chanx_right_in[0] , chanx_left_in[2] , 
        chanx_right_in[2] , chanx_left_in[6] , chanx_right_in[6] , 
        chanx_left_in[12] , chanx_right_in[12] , chanx_left_in[16] , 
        chanx_right_in[16] } ) ,
    .sram ( mux_tree_tapbuf_size10_6_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size10_6_sram_inv ) , 
    .out ( top_grid_pin_28_ ) , .p0 ( optlc_net_90 ) ) ;
mux_tree_tapbuf_size10_3_1 mux_bottom_ipin_13 (
    .in ( { chanx_left_in[1] , chanx_right_in[1] , chanx_left_in[3] , 
        chanx_right_in[3] , chanx_left_in[7] , chanx_right_in[7] , 
        chanx_left_in[13] , chanx_right_in[13] , chanx_left_in[17] , 
        chanx_right_in[17] } ) ,
    .sram ( mux_tree_tapbuf_size10_7_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size10_7_sram_inv ) , 
    .out ( top_grid_pin_29_ ) , .p0 ( optlc_net_90 ) ) ;
mux_tree_tapbuf_size10_12 mux_top_ipin_0 (
    .in ( { chanx_left_in[0] , chanx_right_in[0] , chanx_left_in[2] , 
        chanx_right_in[2] , chanx_left_in[4] , chanx_right_in[4] , 
        chanx_left_in[10] , chanx_right_in[10] , chanx_left_in[16] , 
        chanx_right_in[16] } ) ,
    .sram ( mux_tree_tapbuf_size10_8_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size10_8_sram_inv ) , 
    .out ( bottom_grid_pin_0_ ) , .p0 ( optlc_net_90 ) ) ;
mux_tree_tapbuf_size10_mem_0_2 mem_bottom_ipin_0 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( ccff_head ) , 
    .ccff_tail ( mux_tree_tapbuf_size10_mem_0_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size10_0_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size10_0_sram_inv ) ) ;
mux_tree_tapbuf_size10_mem_1_1 mem_bottom_ipin_1 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size10_mem_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size10_mem_1_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size10_1_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size10_1_sram_inv ) ) ;
mux_tree_tapbuf_size10_mem_4_1 mem_bottom_ipin_4 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size8_mem_1_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size10_mem_2_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size10_2_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size10_2_sram_inv ) ) ;
mux_tree_tapbuf_size10_mem_5_1 mem_bottom_ipin_5 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size10_mem_2_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size10_mem_3_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size10_3_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size10_3_sram_inv ) ) ;
mux_tree_tapbuf_size10_mem_6_1 mem_bottom_ipin_8 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size8_mem_3_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size10_mem_4_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size10_4_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size10_4_sram_inv ) ) ;
mux_tree_tapbuf_size10_mem_7_1 mem_bottom_ipin_9 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size10_mem_4_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size10_mem_5_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size10_5_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size10_5_sram_inv ) ) ;
mux_tree_tapbuf_size10_mem_2_1 mem_bottom_ipin_12 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size8_mem_5_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size10_mem_6_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size10_6_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size10_6_sram_inv ) ) ;
mux_tree_tapbuf_size10_mem_3_1 mem_bottom_ipin_13 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size10_mem_6_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size10_mem_7_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size10_7_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size10_7_sram_inv ) ) ;
mux_tree_tapbuf_size10_mem_12 mem_top_ipin_0 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size8_mem_7_ccff_tail ) , 
    .ccff_tail ( ccff_tail ) , .mem_out ( mux_tree_tapbuf_size10_8_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size10_8_sram_inv ) ) ;
mux_tree_tapbuf_size8_4 mux_bottom_ipin_2 (
    .in ( { chanx_left_in[0] , chanx_right_in[0] , chanx_left_in[2] , 
        chanx_right_in[2] , chanx_left_in[6] , chanx_right_in[6] , 
        chanx_left_in[14] , chanx_right_in[14] } ) ,
    .sram ( mux_tree_tapbuf_size8_0_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size8_0_sram_inv ) , 
    .out ( top_grid_pin_18_ ) , .p0 ( optlc_net_90 ) ) ;
mux_tree_tapbuf_size8_5 mux_bottom_ipin_3 (
    .in ( { chanx_left_in[1] , chanx_right_in[1] , chanx_left_in[3] , 
        chanx_right_in[3] , chanx_left_in[7] , chanx_right_in[7] , 
        chanx_left_in[15] , chanx_right_in[15] } ) ,
    .sram ( mux_tree_tapbuf_size8_1_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size8_1_sram_inv ) , 
    .out ( top_grid_pin_19_ ) , .p0 ( optlc_net_91 ) ) ;
mux_tree_tapbuf_size8_6 mux_bottom_ipin_6 (
    .in ( { chanx_left_in[0] , chanx_right_in[0] , chanx_left_in[2] , 
        chanx_right_in[2] , chanx_left_in[10] , chanx_right_in[10] , 
        chanx_left_in[18] , chanx_right_in[18] } ) ,
    .sram ( mux_tree_tapbuf_size8_2_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size8_2_sram_inv ) , 
    .out ( top_grid_pin_22_ ) , .p0 ( optlc_net_90 ) ) ;
mux_tree_tapbuf_size8_7 mux_bottom_ipin_7 (
    .in ( { chanx_left_in[1] , chanx_right_in[1] , chanx_left_in[3] , 
        chanx_right_in[3] , chanx_left_in[11] , chanx_right_in[11] , 
        chanx_left_in[19] , chanx_right_in[19] } ) ,
    .sram ( mux_tree_tapbuf_size8_3_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size8_3_sram_inv ) , 
    .out ( top_grid_pin_23_ ) , .p0 ( optlc_net_91 ) ) ;
mux_tree_tapbuf_size8_0_2 mux_bottom_ipin_10 (
    .in ( { chanx_left_in[0] , chanx_right_in[0] , chanx_left_in[2] , 
        chanx_right_in[2] , chanx_left_in[6] , chanx_right_in[6] , 
        chanx_left_in[14] , chanx_right_in[14] } ) ,
    .sram ( mux_tree_tapbuf_size8_4_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size8_4_sram_inv ) , 
    .out ( top_grid_pin_26_ ) , .p0 ( optlc_net_91 ) ) ;
mux_tree_tapbuf_size8_1_2 mux_bottom_ipin_11 (
    .in ( { chanx_left_in[1] , chanx_right_in[1] , chanx_left_in[3] , 
        chanx_right_in[3] , chanx_left_in[7] , chanx_right_in[7] , 
        chanx_left_in[15] , chanx_right_in[15] } ) ,
    .sram ( mux_tree_tapbuf_size8_5_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size8_5_sram_inv ) , 
    .out ( top_grid_pin_27_ ) , .p0 ( optlc_net_91 ) ) ;
mux_tree_tapbuf_size8_2_1 mux_bottom_ipin_14 (
    .in ( { chanx_left_in[0] , chanx_right_in[0] , chanx_left_in[2] , 
        chanx_right_in[2] , chanx_left_in[10] , chanx_right_in[10] , 
        chanx_left_in[18] , chanx_right_in[18] } ) ,
    .sram ( mux_tree_tapbuf_size8_6_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size8_6_sram_inv ) , 
    .out ( top_grid_pin_30_ ) , .p0 ( optlc_net_90 ) ) ;
mux_tree_tapbuf_size8_3 mux_bottom_ipin_15 (
    .in ( { chanx_left_in[1] , chanx_right_in[1] , chanx_left_in[3] , 
        chanx_right_in[3] , chanx_left_in[11] , chanx_right_in[11] , 
        chanx_left_in[19] , chanx_right_in[19] } ) ,
    .sram ( mux_tree_tapbuf_size8_7_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size8_7_sram_inv ) , 
    .out ( top_grid_pin_31_ ) , .p0 ( optlc_net_90 ) ) ;
mux_tree_tapbuf_size8_mem_4 mem_bottom_ipin_2 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size10_mem_1_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size8_mem_0_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size8_0_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size8_0_sram_inv ) ) ;
mux_tree_tapbuf_size8_mem_5 mem_bottom_ipin_3 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size8_mem_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size8_mem_1_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size8_1_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size8_1_sram_inv ) ) ;
mux_tree_tapbuf_size8_mem_6 mem_bottom_ipin_6 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size10_mem_3_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size8_mem_2_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size8_2_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size8_2_sram_inv ) ) ;
mux_tree_tapbuf_size8_mem_7 mem_bottom_ipin_7 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size8_mem_2_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size8_mem_3_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size8_3_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size8_3_sram_inv ) ) ;
mux_tree_tapbuf_size8_mem_0_2 mem_bottom_ipin_10 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size10_mem_5_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size8_mem_4_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size8_4_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size8_4_sram_inv ) ) ;
mux_tree_tapbuf_size8_mem_1_2 mem_bottom_ipin_11 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size8_mem_4_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size8_mem_5_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size8_5_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size8_5_sram_inv ) ) ;
mux_tree_tapbuf_size8_mem_2_1 mem_bottom_ipin_14 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size10_mem_7_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size8_mem_6_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size8_6_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size8_6_sram_inv ) ) ;
mux_tree_tapbuf_size8_mem_3 mem_bottom_ipin_15 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size8_mem_6_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size8_mem_7_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size8_7_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size8_7_sram_inv ) ) ;
sky130_fd_sc_hd__dlygate4sd1_1 FTB_1__0 ( .A ( chanx_left_in[0] ) , 
    .X ( chanx_right_out[0] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_2__1 ( .A ( chanx_left_in[1] ) , 
    .X ( chanx_right_out[1] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_4__3 ( .A ( chanx_left_in[3] ) , 
    .X ( chanx_right_out[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd1_1 FTB_5__4 ( .A ( chanx_left_in[4] ) , 
    .X ( chanx_right_out[4] ) ) ;
sky130_fd_sc_hd__conb_1 optlc_89 ( .LO ( SYNOPSYS_UNCONNECTED_1 ) , 
    .HI ( optlc_net_90 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_8__7 ( .A ( chanx_left_in[7] ) , 
    .X ( chanx_right_out[7] ) ) ;
sky130_fd_sc_hd__conb_1 optlc_91 ( .LO ( SYNOPSYS_UNCONNECTED_2 ) , 
    .HI ( optlc_net_91 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_670 ( .A ( ropt_net_92 ) , 
    .X ( chanx_left_out[4] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_672 ( .A ( chanx_left_in[2] ) , 
    .X ( chanx_right_out[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd1_1 FTB_12__11 ( .A ( chanx_left_in[11] ) , 
    .X ( chanx_right_out[11] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_13__12 ( .A ( chanx_left_in[12] ) , 
    .X ( chanx_right_out[12] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_673 ( .A ( chanx_left_in[6] ) , 
    .X ( chanx_right_out[6] ) ) ;
sky130_fd_sc_hd__dlygate4sd1_1 FTB_15__14 ( .A ( chanx_left_in[14] ) , 
    .X ( chanx_right_out[14] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_16__15 ( .A ( chanx_left_in[15] ) , 
    .X ( chanx_right_out[15] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_679 ( .A ( chanx_right_in[1] ) , 
    .X ( chanx_left_out[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_18__17 ( .A ( chanx_left_in[17] ) , 
    .X ( aps_rename_2_ ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_20__19 ( .A ( chanx_left_in[19] ) , 
    .X ( chanx_right_out[19] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_23__22 ( .A ( chanx_right_in[2] ) , 
    .X ( chanx_left_out[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd1_1 FTB_24__23 ( .A ( chanx_right_in[3] ) , 
    .X ( chanx_left_out[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd1_1 FTB_25__24 ( .A ( chanx_right_in[4] ) , 
    .X ( ropt_net_92 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_26__25 ( .A ( chanx_right_in[5] ) , 
    .X ( chanx_left_out[5] ) ) ;
sky130_fd_sc_hd__dlygate4sd1_1 FTB_27__26 ( .A ( chanx_right_in[6] ) , 
    .X ( chanx_left_out[6] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_28__27 ( .A ( chanx_right_in[7] ) , 
    .X ( chanx_left_out[7] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_29__28 ( .A ( chanx_right_in[8] ) , 
    .X ( chanx_left_out[8] ) ) ;
sky130_fd_sc_hd__dlygate4sd1_1 FTB_30__29 ( .A ( chanx_right_in[9] ) , 
    .X ( chanx_left_out[9] ) ) ;
sky130_fd_sc_hd__dlygate4sd1_1 FTB_33__32 ( .A ( chanx_right_in[12] ) , 
    .X ( chanx_left_out[12] ) ) ;
sky130_fd_sc_hd__dlygate4sd1_1 FTB_34__33 ( .A ( chanx_right_in[13] ) , 
    .X ( chanx_left_out[13] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_35__34 ( .A ( chanx_right_in[14] ) , 
    .X ( chanx_left_out[14] ) ) ;
sky130_fd_sc_hd__dlygate4sd1_1 FTB_36__35 ( .A ( chanx_right_in[15] ) , 
    .X ( chanx_left_out[15] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_37__36 ( .A ( chanx_right_in[16] ) , 
    .X ( aps_rename_1_ ) ) ;
sky130_fd_sc_hd__dlygate4sd1_1 FTB_40__39 ( .A ( chanx_right_in[19] ) , 
    .X ( chanx_left_out[19] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_RR_60 ( .A ( chanx_left_in[5] ) , 
    .X ( chanx_right_out[5] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_RR_61 ( .A ( chanx_left_in[8] ) , 
    .X ( chanx_right_out[8] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_RR_62 ( .A ( chanx_left_in[9] ) , 
    .X ( chanx_right_out[9] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_RR_68 ( .A ( chanx_right_in[18] ) , 
    .X ( chanx_left_out[18] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_RR_70 ( .A ( chanx_left_in[16] ) , 
    .X ( chanx_right_out[16] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_RR_71 ( .A ( chanx_left_in[18] ) , 
    .X ( chanx_right_out[18] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 BUFT_RR_73 ( .A ( aps_rename_1_ ) , 
    .X ( chanx_left_out[16] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_P_76 ( .A ( chanx_right_in[0] ) , 
    .X ( chanx_left_out[0] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_P_77 ( .A ( chanx_right_in[10] ) , 
    .X ( chanx_left_out[10] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_P_78 ( .A ( chanx_right_in[11] ) , 
    .X ( chanx_left_out[11] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_P_81 ( .A ( chanx_left_in[10] ) , 
    .X ( chanx_right_out[10] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_P_82 ( .A ( chanx_left_in[13] ) , 
    .X ( chanx_right_out[13] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 BUFT_P_83 ( .A ( aps_rename_2_ ) , 
    .X ( chanx_right_out[17] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_P_85 ( .A ( chanx_right_in[17] ) , 
    .X ( chanx_left_out[17] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_15_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd1_1 FTB_24__39 ( .A ( mem_out[1] ) , 
    .X ( net_net_59 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_86 ( .A ( net_net_59 ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_22 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_23__38 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_16_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_22__37 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_14_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_21__36 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_13_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_20__35 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_12_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_19__34 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_11_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_18__33 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_10_2 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_17__32 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_9_2 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_16__31 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_8_2 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_15__30 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_7_2 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_14__29 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_6_3 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_13__28 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_5_4 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_12__27 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_4_4 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_11__26 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_3_5 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_10__25 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_2_5 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_9__24 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_1_5 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_8__23 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_0_5 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_7__22 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_39 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_15_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_39 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
endmodule


module const1_22_7 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_22 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_22_7 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
endmodule


module const1_21_7 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_16_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_21_7 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
endmodule


module const1_20_7 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_14_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_20_7 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
endmodule


module const1_19_7 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_13_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_19_7 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
endmodule


module const1_18_7 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_12_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;

const1_18_7 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_8 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , .X ( out[0] ) ) ;
endmodule


module const1_17_7 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_11_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_17_7 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
endmodule


module const1_16_8 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_10_2 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_16_8 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
endmodule


module const1_15_8 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_9_2 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_15_8 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_42 ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
endmodule


module const1_14_8 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_8_2 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_14_8 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
endmodule


module const1_13_8 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_7_2 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_13_8 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
endmodule


module const1_12_8 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_6_3 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_12_8 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
endmodule


module const1_11_8 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_5_4 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_11_8 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
endmodule


module const1_10_8 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_4_4 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_10_8 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
endmodule


module const1_9_8 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_3_5 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_9_8 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
endmodule


module const1_8_8 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_2_5 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_8_8 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
endmodule


module const1_7_8 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_1_5 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_7_8 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
endmodule


module const1_6_9 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_0_5 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_6_9 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
endmodule


module mux_tree_tapbuf_size3_mem_0_6 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_6__21 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size3_mem_11 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_5__20 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_5_9 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size3_0_6 ( in , sram , sram_inv , out , p0 ) ;
input  [0:2] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;

const1_5_9 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( p0 ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_41 ( 
    .A ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .X ( BUF_net_41 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_P_88 ( .A ( BUF_net_41 ) , 
    .X ( out[0] ) ) ;
endmodule


module const1_4_9 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size3_11 ( in , sram , sram_inv , out , p0 ) ;
input  [0:2] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;

const1_4_9 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( p0 ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
endmodule


module mux_tree_tapbuf_size5_mem_8 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_4__19 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size5_mem_0_4 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_3__18 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_3_9 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size5_8 ( in , sram , sram_inv , out , p0 ) ;
input  [0:4] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;

const1_3_9 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , .A1 ( in[4] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
endmodule


module const1_2_9 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size5_0_4 ( in , sram , sram_inv , out , p0 ) ;
input  [0:4] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;

const1_2_9 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , .A1 ( in[4] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_P_87 ( 
    .A ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .X ( out[0] ) ) ;
endmodule


module mux_tree_tapbuf_size6_mem_10 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_2__17 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size6_mem_0_6 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_1__16 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_1_9 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size6_10 ( in , sram , sram_inv , out , p0 ) ;
input  [0:5] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;

const1_1_9 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
endmodule


module const1_0_9 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size6_0_6 ( in , sram , sram_inv , out , p0 ) ;
input  [0:5] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;

const1_0_9 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
endmodule


module sb_2__2_ ( prog_clk , chany_bottom_in , bottom_right_grid_pin_1_ , 
    bottom_left_grid_pin_34_ , bottom_left_grid_pin_35_ , 
    bottom_left_grid_pin_36_ , bottom_left_grid_pin_37_ , 
    bottom_left_grid_pin_38_ , bottom_left_grid_pin_39_ , 
    bottom_left_grid_pin_40_ , bottom_left_grid_pin_41_ , chanx_left_in , 
    left_top_grid_pin_1_ , ccff_head , chany_bottom_out , chanx_left_out , 
    ccff_tail ) ;
input  [0:0] prog_clk ;
input  [0:19] chany_bottom_in ;
input  [0:0] bottom_right_grid_pin_1_ ;
input  [0:0] bottom_left_grid_pin_34_ ;
input  [0:0] bottom_left_grid_pin_35_ ;
input  [0:0] bottom_left_grid_pin_36_ ;
input  [0:0] bottom_left_grid_pin_37_ ;
input  [0:0] bottom_left_grid_pin_38_ ;
input  [0:0] bottom_left_grid_pin_39_ ;
input  [0:0] bottom_left_grid_pin_40_ ;
input  [0:0] bottom_left_grid_pin_41_ ;
input  [0:19] chanx_left_in ;
input  [0:0] left_top_grid_pin_1_ ;
input  [0:0] ccff_head ;
output [0:19] chany_bottom_out ;
output [0:19] chanx_left_out ;
output [0:0] ccff_tail ;

wire [0:1] mux_tree_tapbuf_size2_0_sram ;
wire [0:1] mux_tree_tapbuf_size2_0_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_10_sram ;
wire [0:1] mux_tree_tapbuf_size2_10_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_11_sram ;
wire [0:1] mux_tree_tapbuf_size2_11_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_12_sram ;
wire [0:1] mux_tree_tapbuf_size2_12_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_13_sram ;
wire [0:1] mux_tree_tapbuf_size2_13_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_14_sram ;
wire [0:1] mux_tree_tapbuf_size2_14_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_15_sram ;
wire [0:1] mux_tree_tapbuf_size2_15_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_16_sram ;
wire [0:1] mux_tree_tapbuf_size2_16_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_17_sram ;
wire [0:1] mux_tree_tapbuf_size2_17_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_1_sram ;
wire [0:1] mux_tree_tapbuf_size2_1_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_2_sram ;
wire [0:1] mux_tree_tapbuf_size2_2_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_3_sram ;
wire [0:1] mux_tree_tapbuf_size2_3_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_4_sram ;
wire [0:1] mux_tree_tapbuf_size2_4_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_5_sram ;
wire [0:1] mux_tree_tapbuf_size2_5_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_6_sram ;
wire [0:1] mux_tree_tapbuf_size2_6_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_7_sram ;
wire [0:1] mux_tree_tapbuf_size2_7_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_8_sram ;
wire [0:1] mux_tree_tapbuf_size2_8_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_9_sram ;
wire [0:1] mux_tree_tapbuf_size2_9_sram_inv ;
wire [0:0] mux_tree_tapbuf_size2_mem_0_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_10_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_11_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_12_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_13_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_14_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_15_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_16_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_1_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_2_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_3_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_4_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_5_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_6_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_7_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_8_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_9_ccff_tail ;
wire [0:1] mux_tree_tapbuf_size3_0_sram ;
wire [0:1] mux_tree_tapbuf_size3_0_sram_inv ;
wire [0:1] mux_tree_tapbuf_size3_1_sram ;
wire [0:1] mux_tree_tapbuf_size3_1_sram_inv ;
wire [0:0] mux_tree_tapbuf_size3_mem_0_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size3_mem_1_ccff_tail ;
wire [0:2] mux_tree_tapbuf_size5_0_sram ;
wire [0:2] mux_tree_tapbuf_size5_0_sram_inv ;
wire [0:2] mux_tree_tapbuf_size5_1_sram ;
wire [0:2] mux_tree_tapbuf_size5_1_sram_inv ;
wire [0:0] mux_tree_tapbuf_size5_mem_0_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size5_mem_1_ccff_tail ;
wire [0:2] mux_tree_tapbuf_size6_0_sram ;
wire [0:2] mux_tree_tapbuf_size6_0_sram_inv ;
wire [0:2] mux_tree_tapbuf_size6_1_sram ;
wire [0:2] mux_tree_tapbuf_size6_1_sram_inv ;
wire [0:0] mux_tree_tapbuf_size6_mem_0_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size6_mem_1_ccff_tail ;

mux_tree_tapbuf_size6_0_6 mux_bottom_track_1 (
    .in ( { bottom_right_grid_pin_1_[0] , bottom_left_grid_pin_35_[0] , 
        bottom_left_grid_pin_37_[0] , bottom_left_grid_pin_39_[0] , 
        bottom_left_grid_pin_41_[0] , chanx_left_in[1] } ) ,
    .sram ( mux_tree_tapbuf_size6_0_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size6_0_sram_inv ) , 
    .out ( chany_bottom_out[0] ) , .p0 ( optlc_net_114 ) ) ;
mux_tree_tapbuf_size6_10 mux_bottom_track_5 (
    .in ( { bottom_right_grid_pin_1_[0] , bottom_left_grid_pin_35_[0] , 
        bottom_left_grid_pin_37_[0] , bottom_left_grid_pin_39_[0] , 
        bottom_left_grid_pin_41_[0] , chanx_left_in[3] } ) ,
    .sram ( mux_tree_tapbuf_size6_1_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size6_1_sram_inv ) , 
    .out ( chany_bottom_out[2] ) , .p0 ( optlc_net_114 ) ) ;
mux_tree_tapbuf_size6_mem_0_6 mem_bottom_track_1 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( ccff_head ) , 
    .ccff_tail ( mux_tree_tapbuf_size6_mem_0_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size6_0_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size6_0_sram_inv ) ) ;
mux_tree_tapbuf_size6_mem_10 mem_bottom_track_5 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size5_mem_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size6_mem_1_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size6_1_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size6_1_sram_inv ) ) ;
mux_tree_tapbuf_size5_0_4 mux_bottom_track_3 (
    .in ( { bottom_left_grid_pin_34_[0] , bottom_left_grid_pin_36_[0] , 
        bottom_left_grid_pin_38_[0] , bottom_left_grid_pin_40_[0] , 
        chanx_left_in[2] } ) ,
    .sram ( mux_tree_tapbuf_size5_0_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size5_0_sram_inv ) ,
    .out ( { ropt_net_123 } ) ,
    .p0 ( optlc_net_114 ) ) ;
mux_tree_tapbuf_size5_8 mux_bottom_track_7 (
    .in ( { bottom_left_grid_pin_34_[0] , bottom_left_grid_pin_36_[0] , 
        bottom_left_grid_pin_38_[0] , bottom_left_grid_pin_40_[0] , 
        chanx_left_in[4] } ) ,
    .sram ( mux_tree_tapbuf_size5_1_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size5_1_sram_inv ) , 
    .out ( chany_bottom_out[3] ) , .p0 ( optlc_net_114 ) ) ;
mux_tree_tapbuf_size5_mem_0_4 mem_bottom_track_3 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size6_mem_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size5_mem_0_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size5_0_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size5_0_sram_inv ) ) ;
mux_tree_tapbuf_size5_mem_8 mem_bottom_track_7 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size6_mem_1_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size5_mem_1_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size5_1_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size5_1_sram_inv ) ) ;
mux_tree_tapbuf_size3_11 mux_bottom_track_9 (
    .in ( { bottom_right_grid_pin_1_[0] , bottom_left_grid_pin_41_[0] , 
        chanx_left_in[5] } ) ,
    .sram ( mux_tree_tapbuf_size3_0_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size3_0_sram_inv ) , 
    .out ( chany_bottom_out[4] ) , .p0 ( optlc_net_114 ) ) ;
mux_tree_tapbuf_size3_0_6 mux_bottom_track_25 (
    .in ( { bottom_right_grid_pin_1_[0] , bottom_left_grid_pin_41_[0] , 
        chanx_left_in[13] } ) ,
    .sram ( mux_tree_tapbuf_size3_1_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size3_1_sram_inv ) ,
    .out ( { ropt_net_130 } ) ,
    .p0 ( optlc_net_115 ) ) ;
mux_tree_tapbuf_size3_mem_11 mem_bottom_track_9 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size5_mem_1_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size3_mem_0_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size3_0_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size3_0_sram_inv ) ) ;
mux_tree_tapbuf_size3_mem_0_6 mem_bottom_track_25 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_6_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size3_mem_1_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size3_1_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size3_1_sram_inv ) ) ;
mux_tree_tapbuf_size2_0_5 mux_bottom_track_11 (
    .in ( { bottom_left_grid_pin_34_[0] , chanx_left_in[6] } ) ,
    .sram ( mux_tree_tapbuf_size2_0_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_0_sram_inv ) , 
    .out ( chany_bottom_out[5] ) , .p0 ( optlc_net_114 ) ) ;
mux_tree_tapbuf_size2_1_5 mux_bottom_track_13 (
    .in ( { bottom_left_grid_pin_35_[0] , chanx_left_in[7] } ) ,
    .sram ( mux_tree_tapbuf_size2_1_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_1_sram_inv ) , 
    .out ( chany_bottom_out[6] ) , .p0 ( optlc_net_115 ) ) ;
mux_tree_tapbuf_size2_2_5 mux_bottom_track_15 (
    .in ( { bottom_left_grid_pin_36_[0] , chanx_left_in[8] } ) ,
    .sram ( mux_tree_tapbuf_size2_2_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_2_sram_inv ) , 
    .out ( chany_bottom_out[7] ) , .p0 ( optlc_net_115 ) ) ;
mux_tree_tapbuf_size2_3_5 mux_bottom_track_17 (
    .in ( { bottom_left_grid_pin_37_[0] , chanx_left_in[9] } ) ,
    .sram ( mux_tree_tapbuf_size2_3_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_3_sram_inv ) , 
    .out ( chany_bottom_out[8] ) , .p0 ( optlc_net_112 ) ) ;
mux_tree_tapbuf_size2_4_4 mux_bottom_track_19 (
    .in ( { bottom_left_grid_pin_38_[0] , chanx_left_in[10] } ) ,
    .sram ( mux_tree_tapbuf_size2_4_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_4_sram_inv ) , 
    .out ( chany_bottom_out[9] ) , .p0 ( optlc_net_114 ) ) ;
mux_tree_tapbuf_size2_5_4 mux_bottom_track_21 (
    .in ( { bottom_left_grid_pin_39_[0] , chanx_left_in[11] } ) ,
    .sram ( mux_tree_tapbuf_size2_5_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_5_sram_inv ) , 
    .out ( chany_bottom_out[10] ) , .p0 ( optlc_net_115 ) ) ;
mux_tree_tapbuf_size2_6_3 mux_bottom_track_23 (
    .in ( { bottom_left_grid_pin_40_[0] , chanx_left_in[12] } ) ,
    .sram ( mux_tree_tapbuf_size2_6_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_6_sram_inv ) , 
    .out ( chany_bottom_out[11] ) , .p0 ( optlc_net_113 ) ) ;
mux_tree_tapbuf_size2_7_2 mux_bottom_track_27 (
    .in ( { bottom_left_grid_pin_34_[0] , chanx_left_in[14] } ) ,
    .sram ( mux_tree_tapbuf_size2_7_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_7_sram_inv ) , 
    .out ( chany_bottom_out[13] ) , .p0 ( optlc_net_114 ) ) ;
mux_tree_tapbuf_size2_8_2 mux_bottom_track_29 (
    .in ( { bottom_left_grid_pin_35_[0] , chanx_left_in[15] } ) ,
    .sram ( mux_tree_tapbuf_size2_8_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_8_sram_inv ) , 
    .out ( chany_bottom_out[14] ) , .p0 ( optlc_net_115 ) ) ;
mux_tree_tapbuf_size2_9_2 mux_bottom_track_31 (
    .in ( { bottom_left_grid_pin_36_[0] , chanx_left_in[16] } ) ,
    .sram ( mux_tree_tapbuf_size2_9_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_9_sram_inv ) ,
    .out ( { ropt_net_120 } ) ,
    .p0 ( optlc_net_115 ) ) ;
mux_tree_tapbuf_size2_10_2 mux_bottom_track_33 (
    .in ( { bottom_left_grid_pin_37_[0] , chanx_left_in[17] } ) ,
    .sram ( mux_tree_tapbuf_size2_10_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_10_sram_inv ) , 
    .out ( chany_bottom_out[16] ) , .p0 ( optlc_net_112 ) ) ;
mux_tree_tapbuf_size2_11_1 mux_bottom_track_35 (
    .in ( { bottom_left_grid_pin_38_[0] , chanx_left_in[18] } ) ,
    .sram ( mux_tree_tapbuf_size2_11_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_11_sram_inv ) , 
    .out ( chany_bottom_out[17] ) , .p0 ( optlc_net_112 ) ) ;
mux_tree_tapbuf_size2_12_1 mux_bottom_track_37 (
    .in ( { bottom_left_grid_pin_39_[0] , chanx_left_in[19] } ) ,
    .sram ( mux_tree_tapbuf_size2_12_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_12_sram_inv ) , 
    .out ( chany_bottom_out[18] ) , .p0 ( optlc_net_115 ) ) ;
mux_tree_tapbuf_size2_13_1 mux_bottom_track_39 (
    .in ( { bottom_left_grid_pin_40_[0] , chanx_left_in[0] } ) ,
    .sram ( mux_tree_tapbuf_size2_13_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_13_sram_inv ) , 
    .out ( chany_bottom_out[19] ) , .p0 ( optlc_net_114 ) ) ;
mux_tree_tapbuf_size2_14_1 mux_left_track_1 (
    .in ( { chany_bottom_in[19] , left_top_grid_pin_1_[0] } ) ,
    .sram ( mux_tree_tapbuf_size2_14_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_14_sram_inv ) , 
    .out ( chanx_left_out[0] ) , .p0 ( optlc_net_113 ) ) ;
mux_tree_tapbuf_size2_16_1 mux_left_track_5 (
    .in ( { chany_bottom_in[1] , left_top_grid_pin_1_[0] } ) ,
    .sram ( mux_tree_tapbuf_size2_15_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_15_sram_inv ) , 
    .out ( chanx_left_out[2] ) , .p0 ( optlc_net_113 ) ) ;
mux_tree_tapbuf_size2_22 mux_left_track_9 (
    .in ( { chany_bottom_in[3] , left_top_grid_pin_1_[0] } ) ,
    .sram ( mux_tree_tapbuf_size2_16_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_16_sram_inv ) , 
    .out ( chanx_left_out[4] ) , .p0 ( optlc_net_113 ) ) ;
mux_tree_tapbuf_size2_15_1 mux_left_track_25 (
    .in ( { chany_bottom_in[11] , left_top_grid_pin_1_[0] } ) ,
    .sram ( mux_tree_tapbuf_size2_17_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_17_sram_inv ) , 
    .out ( chanx_left_out[12] ) , .p0 ( optlc_net_113 ) ) ;
mux_tree_tapbuf_size2_mem_0_5 mem_bottom_track_11 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size3_mem_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_0_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_0_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_0_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem_1_5 mem_bottom_track_13 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_1_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_1_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_1_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem_2_5 mem_bottom_track_15 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_1_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_2_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_2_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_2_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem_3_5 mem_bottom_track_17 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_2_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_3_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_3_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_3_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem_4_4 mem_bottom_track_19 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_3_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_4_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_4_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_4_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem_5_4 mem_bottom_track_21 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_4_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_5_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_5_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_5_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem_6_3 mem_bottom_track_23 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_5_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_6_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_6_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_6_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem_7_2 mem_bottom_track_27 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size3_mem_1_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_7_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_7_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_7_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem_8_2 mem_bottom_track_29 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_7_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_8_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_8_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_8_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem_9_2 mem_bottom_track_31 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_8_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_9_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_9_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_9_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem_10_2 mem_bottom_track_33 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_9_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_10_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_10_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_10_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem_11_1 mem_bottom_track_35 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_10_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_11_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_11_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_11_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem_12_1 mem_bottom_track_37 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_11_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_12_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_12_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_12_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem_13_1 mem_bottom_track_39 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_12_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_13_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_13_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_13_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem_14_1 mem_left_track_1 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_13_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_14_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_14_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_14_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem_16_1 mem_left_track_5 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_14_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_15_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_15_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_15_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem_22 mem_left_track_9 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_15_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_16_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_16_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_16_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem_15_1 mem_left_track_25 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_16_ccff_tail ) ,
    .ccff_tail ( { ropt_net_128 } ) ,
    .mem_out ( mux_tree_tapbuf_size2_17_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_17_sram_inv ) ) ;
sky130_fd_sc_hd__conb_1 optlc_107 ( .LO ( SYNOPSYS_UNCONNECTED_1 ) , 
    .HI ( optlc_net_112 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_109 ( .LO ( SYNOPSYS_UNCONNECTED_2 ) , 
    .HI ( optlc_net_113 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_111 ( .LO ( SYNOPSYS_UNCONNECTED_3 ) , 
    .HI ( optlc_net_114 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_113 ( .LO ( SYNOPSYS_UNCONNECTED_4 ) , 
    .HI ( optlc_net_115 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_703 ( .A ( chany_bottom_in[2] ) , 
    .X ( chanx_left_out[3] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_704 ( .A ( chany_bottom_in[7] ) , 
    .X ( ropt_net_138 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_705 ( 
    .A ( chany_bottom_in[16] ) , .X ( chanx_left_out[17] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_706 ( .A ( ropt_net_120 ) , 
    .X ( ropt_net_137 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_707 ( 
    .A ( chany_bottom_in[17] ) , .X ( chanx_left_out[18] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_708 ( .A ( chany_bottom_in[8] ) , 
    .X ( chanx_left_out[9] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_709 ( .A ( ropt_net_123 ) , 
    .X ( ropt_net_141 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_710 ( 
    .A ( chany_bottom_in[15] ) , .X ( ropt_net_135 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_711 ( .A ( chany_bottom_in[0] ) , 
    .X ( chanx_left_out[1] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_712 ( 
    .A ( chany_bottom_in[12] ) , .X ( ropt_net_134 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_719 ( .A ( ropt_net_133 ) , 
    .X ( chanx_left_out[6] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_713 ( 
    .A ( chany_bottom_in[18] ) , .X ( chanx_left_out[19] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_714 ( .A ( ropt_net_128 ) , 
    .X ( ropt_net_140 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_715 ( .A ( ropt_net_129 ) , 
    .X ( ropt_net_136 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_46 ( .A ( chany_bottom_in[4] ) , 
    .X ( BUF_net_46 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_47 ( .A ( chany_bottom_in[5] ) , 
    .X ( ropt_net_131 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_716 ( .A ( ropt_net_130 ) , 
    .X ( chany_bottom_out[12] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_720 ( .A ( ropt_net_134 ) , 
    .X ( chanx_left_out[13] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_721 ( .A ( ropt_net_135 ) , 
    .X ( chanx_left_out[16] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_51 ( .A ( chany_bottom_in[9] ) , 
    .X ( BUF_net_51 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_52 ( .A ( chany_bottom_in[10] ) , 
    .X ( BUF_net_52 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_722 ( .A ( ropt_net_136 ) , 
    .X ( chanx_left_out[7] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_54 ( .A ( chany_bottom_in[13] ) , 
    .X ( BUF_net_54 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_55 ( .A ( chany_bottom_in[14] ) , 
    .X ( BUF_net_55 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_718 ( .A ( ropt_net_131 ) , 
    .X ( ropt_net_133 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_723 ( .A ( ropt_net_137 ) , 
    .X ( chany_bottom_out[15] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_724 ( .A ( ropt_net_138 ) , 
    .X ( chanx_left_out[8] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_725 ( .A ( ropt_net_139 ) , 
    .X ( chanx_left_out[5] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_726 ( .A ( ropt_net_140 ) , 
    .X ( ccff_tail[0] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_727 ( .A ( ropt_net_141 ) , 
    .X ( chany_bottom_out[1] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 BUFT_P_93 ( .A ( BUF_net_46 ) , 
    .X ( ropt_net_139 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_P_95 ( .A ( chany_bottom_in[6] ) , 
    .X ( ropt_net_129 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 BUFT_P_98 ( .A ( BUF_net_51 ) , 
    .X ( chanx_left_out[10] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 BUFT_P_99 ( .A ( BUF_net_52 ) , 
    .X ( chanx_left_out[11] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 BUFT_P_101 ( .A ( BUF_net_54 ) , 
    .X ( chanx_left_out[14] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 BUFT_P_102 ( .A ( BUF_net_55 ) , 
    .X ( chanx_left_out[15] ) ) ;
endmodule


module mux_tree_tapbuf_size3_mem_10 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_27__59 ( .A ( mem_out[1] ) , 
    .X ( net_net_80 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_79 ( .A ( net_net_80 ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size3_mem_3_3 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_26__58 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size3_mem_2_4 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_25__57 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size3_mem_1_4 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_24__56 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size3_mem_0_5 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_23__55 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_38 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size3_10 ( in , sram , sram_inv , out , p0 ) ;
input  [0:2] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;

const1_38 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( p0 ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
endmodule


module const1_25_6 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size3_3_3 ( in , sram , sram_inv , out , p0 ) ;
input  [0:2] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;

const1_25_6 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( p0 ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
endmodule


module const1_24_6 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size3_2_4 ( in , sram , sram_inv , out , p0 ) ;
input  [0:2] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;

const1_24_6 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( p0 ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
endmodule


module const1_23_6 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size3_1_4 ( in , sram , sram_inv , out , p0 ) ;
input  [0:2] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;

const1_23_6 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( p0 ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
endmodule


module const1_22_6 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size3_0_5 ( in , sram , sram_inv , out , p0 ) ;
input  [0:2] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;

const1_22_6 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( p0 ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
endmodule


module mux_tree_tapbuf_size4_mem_2_2 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_22__54 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size4_mem_1_2 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_21__53 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size4_mem_0_3 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_20__52 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size4_mem_8 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_19__51 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_21_6 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size4_2_2 ( in , sram , sram_inv , out , p0 ) ;
input  [0:3] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;

const1_21_6 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( in[2] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , .A1 ( in[3] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
endmodule


module const1_20_6 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size4_1_2 ( in , sram , sram_inv , out , p0 ) ;
input  [0:3] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;

const1_20_6 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( in[2] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , .A1 ( in[3] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
endmodule


module const1_19_6 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size4_0_3 ( in , sram , sram_inv , out , p0 ) ;
input  [0:3] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;

const1_19_6 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( in[2] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , .A1 ( in[3] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_105 ( 
    .A ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .X ( out[0] ) ) ;
endmodule


module const1_18_6 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size4_8 ( in , sram , sram_inv , out , p0 ) ;
input  [0:3] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;

const1_18_6 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( in[2] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , .A1 ( in[3] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
endmodule


module mux_tree_tapbuf_size9_mem_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_18__50 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_17_6 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size9_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:8] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;

const1_17_6 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[7] ) , .A1 ( in[6] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[8] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 BUFT_P_104 ( 
    .A ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , .X ( out[0] ) ) ;
endmodule


module mux_tree_tapbuf_size6_mem_1_3 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_17__49 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size6_mem_0_5 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_16__48 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size6_mem_9 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_15__47 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_16_7 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size6_1_3 ( in , sram , sram_inv , out , p0 ) ;
input  [0:5] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;

const1_16_7 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
endmodule


module const1_15_7 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size6_0_5 ( in , sram , sram_inv , out , p0 ) ;
input  [0:5] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;

const1_15_7 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
endmodule


module const1_14_7 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size6_9 ( in , sram , sram_inv , out , p0 ) ;
input  [0:5] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;

const1_14_7 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
endmodule


module mux_tree_tapbuf_size7_mem_4_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_14__46 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size7_mem_3_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_13__45 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size7_mem_2_3 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_12__44 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size7_mem_1_4 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_11__43 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size7_mem_0_4 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_10__42 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size7_mem_8 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_9__41 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size7_mem_5_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_8__40 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_13_7 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size7_4_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:6] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;

const1_13_7 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_3_ ( .A0 ( p0 ) , .A1 ( in[6] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
endmodule


module const1_12_7 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size7_3_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:6] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;

const1_12_7 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_3_ ( .A0 ( p0 ) , .A1 ( in[6] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
endmodule


module const1_11_7 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size7_2_3 ( in , sram , sram_inv , out , p0 ) ;
input  [0:6] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;

const1_11_7 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_3_ ( .A0 ( p0 ) , .A1 ( in[6] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
endmodule


module const1_10_7 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size7_1_4 ( in , sram , sram_inv , out , p0 ) ;
input  [0:6] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;

const1_10_7 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_3_ ( .A0 ( p0 ) , .A1 ( in[6] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
endmodule


module const1_9_7 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size7_0_4 ( in , sram , sram_inv , out , p0 ) ;
input  [0:6] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;

const1_9_7 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_3_ ( .A0 ( p0 ) , .A1 ( in[6] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
endmodule


module const1_8_7 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size7_8 ( in , sram , sram_inv , out , p0 ) ;
input  [0:6] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;

const1_8_7 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_3_ ( .A0 ( p0 ) , .A1 ( in[6] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
endmodule


module const1_7_7 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size7_5_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:6] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;

const1_7_7 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_3_ ( .A0 ( p0 ) , .A1 ( in[6] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
endmodule


module mux_tree_tapbuf_size14_mem_0_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_7__39 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size14_mem_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_6__38 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_6_8 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size14_0_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:13] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_10_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_11_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_12_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_13_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

const1_6_8 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_13_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_3_ ( .A0 ( in[7] ) , .A1 ( in[6] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_4_ ( .A0 ( in[9] ) , .A1 ( in[8] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_5_ ( .A0 ( in[11] ) , .A1 ( in[10] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_6_ ( .A0 ( in[13] ) , .A1 ( in[12] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_10_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_11_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_10_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_12_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_12_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_11_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_13_X[0] ) ) ;
endmodule


module const1_5_8 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size14_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:13] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_10_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_11_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_12_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_13_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

const1_5_8 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_13_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_3_ ( .A0 ( in[7] ) , .A1 ( in[6] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_4_ ( .A0 ( in[9] ) , .A1 ( in[8] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_5_ ( .A0 ( in[11] ) , .A1 ( in[10] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_6_ ( .A0 ( in[13] ) , .A1 ( in[12] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_10_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_11_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_10_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_12_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_12_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_11_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_13_X[0] ) ) ;
endmodule


module mux_tree_tapbuf_size8_mem_0_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_5__37 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size8_mem_3 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_4__36 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size8_mem_1_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_3__35 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_4_8 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size8_0_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:7] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;

const1_4_8 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( in[2] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[4] ) , .A1 ( in[3] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[6] ) , .A1 ( in[5] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
endmodule


module const1_3_8 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size8_3 ( in , sram , sram_inv , out , p0 ) ;
input  [0:7] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;

const1_3_8 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( in[2] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[4] ) , .A1 ( in[3] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[6] ) , .A1 ( in[5] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
endmodule


module const1_2_8 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size8_1_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:7] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;

const1_2_8 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( in[2] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[4] ) , .A1 ( in[3] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[6] ) , .A1 ( in[5] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
endmodule


module mux_tree_tapbuf_size10_mem_0_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_2__34 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size10_mem_11 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_1__33 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_1_8 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size10_0_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:9] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

const1_1_8 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[6] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[8] ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[9] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
endmodule


module const1_0_8 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size10_11 ( in , sram , sram_inv , out , p0 ) ;
input  [0:9] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

const1_0_8 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[6] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[8] ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[9] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
endmodule


module sb_2__1_ ( prog_clk , chany_top_in , top_left_grid_pin_34_ , 
    top_left_grid_pin_35_ , top_left_grid_pin_36_ , top_left_grid_pin_37_ , 
    top_left_grid_pin_38_ , top_left_grid_pin_39_ , top_left_grid_pin_40_ , 
    top_left_grid_pin_41_ , top_right_grid_pin_1_ , chany_bottom_in , 
    bottom_right_grid_pin_1_ , bottom_left_grid_pin_34_ , 
    bottom_left_grid_pin_35_ , bottom_left_grid_pin_36_ , 
    bottom_left_grid_pin_37_ , bottom_left_grid_pin_38_ , 
    bottom_left_grid_pin_39_ , bottom_left_grid_pin_40_ , 
    bottom_left_grid_pin_41_ , chanx_left_in , left_top_grid_pin_42_ , 
    left_top_grid_pin_43_ , left_top_grid_pin_44_ , left_top_grid_pin_45_ , 
    left_top_grid_pin_46_ , left_top_grid_pin_47_ , left_top_grid_pin_48_ , 
    left_top_grid_pin_49_ , ccff_head , chany_top_out , chany_bottom_out , 
    chanx_left_out , ccff_tail ) ;
input  [0:0] prog_clk ;
input  [0:19] chany_top_in ;
input  [0:0] top_left_grid_pin_34_ ;
input  [0:0] top_left_grid_pin_35_ ;
input  [0:0] top_left_grid_pin_36_ ;
input  [0:0] top_left_grid_pin_37_ ;
input  [0:0] top_left_grid_pin_38_ ;
input  [0:0] top_left_grid_pin_39_ ;
input  [0:0] top_left_grid_pin_40_ ;
input  [0:0] top_left_grid_pin_41_ ;
input  [0:0] top_right_grid_pin_1_ ;
input  [0:19] chany_bottom_in ;
input  [0:0] bottom_right_grid_pin_1_ ;
input  [0:0] bottom_left_grid_pin_34_ ;
input  [0:0] bottom_left_grid_pin_35_ ;
input  [0:0] bottom_left_grid_pin_36_ ;
input  [0:0] bottom_left_grid_pin_37_ ;
input  [0:0] bottom_left_grid_pin_38_ ;
input  [0:0] bottom_left_grid_pin_39_ ;
input  [0:0] bottom_left_grid_pin_40_ ;
input  [0:0] bottom_left_grid_pin_41_ ;
input  [0:19] chanx_left_in ;
input  [0:0] left_top_grid_pin_42_ ;
input  [0:0] left_top_grid_pin_43_ ;
input  [0:0] left_top_grid_pin_44_ ;
input  [0:0] left_top_grid_pin_45_ ;
input  [0:0] left_top_grid_pin_46_ ;
input  [0:0] left_top_grid_pin_47_ ;
input  [0:0] left_top_grid_pin_48_ ;
input  [0:0] left_top_grid_pin_49_ ;
input  [0:0] ccff_head ;
output [0:19] chany_top_out ;
output [0:19] chany_bottom_out ;
output [0:19] chanx_left_out ;
output [0:0] ccff_tail ;

wire [0:3] mux_tree_tapbuf_size10_0_sram ;
wire [0:3] mux_tree_tapbuf_size10_0_sram_inv ;
wire [0:3] mux_tree_tapbuf_size10_1_sram ;
wire [0:3] mux_tree_tapbuf_size10_1_sram_inv ;
wire [0:0] mux_tree_tapbuf_size10_mem_0_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size10_mem_1_ccff_tail ;
wire [0:3] mux_tree_tapbuf_size14_0_sram ;
wire [0:3] mux_tree_tapbuf_size14_0_sram_inv ;
wire [0:3] mux_tree_tapbuf_size14_1_sram ;
wire [0:3] mux_tree_tapbuf_size14_1_sram_inv ;
wire [0:0] mux_tree_tapbuf_size14_mem_0_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size14_mem_1_ccff_tail ;
wire [0:1] mux_tree_tapbuf_size3_0_sram ;
wire [0:1] mux_tree_tapbuf_size3_0_sram_inv ;
wire [0:1] mux_tree_tapbuf_size3_1_sram ;
wire [0:1] mux_tree_tapbuf_size3_1_sram_inv ;
wire [0:1] mux_tree_tapbuf_size3_2_sram ;
wire [0:1] mux_tree_tapbuf_size3_2_sram_inv ;
wire [0:1] mux_tree_tapbuf_size3_3_sram ;
wire [0:1] mux_tree_tapbuf_size3_3_sram_inv ;
wire [0:1] mux_tree_tapbuf_size3_4_sram ;
wire [0:1] mux_tree_tapbuf_size3_4_sram_inv ;
wire [0:0] mux_tree_tapbuf_size3_mem_0_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size3_mem_1_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size3_mem_2_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size3_mem_3_ccff_tail ;
wire [0:2] mux_tree_tapbuf_size4_0_sram ;
wire [0:2] mux_tree_tapbuf_size4_0_sram_inv ;
wire [0:2] mux_tree_tapbuf_size4_1_sram ;
wire [0:2] mux_tree_tapbuf_size4_1_sram_inv ;
wire [0:2] mux_tree_tapbuf_size4_2_sram ;
wire [0:2] mux_tree_tapbuf_size4_2_sram_inv ;
wire [0:2] mux_tree_tapbuf_size4_3_sram ;
wire [0:2] mux_tree_tapbuf_size4_3_sram_inv ;
wire [0:0] mux_tree_tapbuf_size4_mem_0_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size4_mem_1_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size4_mem_2_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size4_mem_3_ccff_tail ;
wire [0:2] mux_tree_tapbuf_size6_0_sram ;
wire [0:2] mux_tree_tapbuf_size6_0_sram_inv ;
wire [0:2] mux_tree_tapbuf_size6_1_sram ;
wire [0:2] mux_tree_tapbuf_size6_1_sram_inv ;
wire [0:2] mux_tree_tapbuf_size6_2_sram ;
wire [0:2] mux_tree_tapbuf_size6_2_sram_inv ;
wire [0:0] mux_tree_tapbuf_size6_mem_0_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size6_mem_1_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size6_mem_2_ccff_tail ;
wire [0:2] mux_tree_tapbuf_size7_0_sram ;
wire [0:2] mux_tree_tapbuf_size7_0_sram_inv ;
wire [0:2] mux_tree_tapbuf_size7_1_sram ;
wire [0:2] mux_tree_tapbuf_size7_1_sram_inv ;
wire [0:2] mux_tree_tapbuf_size7_2_sram ;
wire [0:2] mux_tree_tapbuf_size7_2_sram_inv ;
wire [0:2] mux_tree_tapbuf_size7_3_sram ;
wire [0:2] mux_tree_tapbuf_size7_3_sram_inv ;
wire [0:2] mux_tree_tapbuf_size7_4_sram ;
wire [0:2] mux_tree_tapbuf_size7_4_sram_inv ;
wire [0:2] mux_tree_tapbuf_size7_5_sram ;
wire [0:2] mux_tree_tapbuf_size7_5_sram_inv ;
wire [0:2] mux_tree_tapbuf_size7_6_sram ;
wire [0:2] mux_tree_tapbuf_size7_6_sram_inv ;
wire [0:0] mux_tree_tapbuf_size7_mem_0_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size7_mem_1_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size7_mem_2_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size7_mem_3_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size7_mem_4_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size7_mem_5_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size7_mem_6_ccff_tail ;
wire [0:3] mux_tree_tapbuf_size8_0_sram ;
wire [0:3] mux_tree_tapbuf_size8_0_sram_inv ;
wire [0:3] mux_tree_tapbuf_size8_1_sram ;
wire [0:3] mux_tree_tapbuf_size8_1_sram_inv ;
wire [0:3] mux_tree_tapbuf_size8_2_sram ;
wire [0:3] mux_tree_tapbuf_size8_2_sram_inv ;
wire [0:0] mux_tree_tapbuf_size8_mem_0_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size8_mem_1_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size8_mem_2_ccff_tail ;
wire [0:3] mux_tree_tapbuf_size9_0_sram ;
wire [0:3] mux_tree_tapbuf_size9_0_sram_inv ;
wire [0:0] mux_tree_tapbuf_size9_mem_0_ccff_tail ;

mux_tree_tapbuf_size10_11 mux_top_track_0 (
    .in ( { top_left_grid_pin_34_[0] , top_left_grid_pin_36_[0] , 
        top_left_grid_pin_38_[0] , top_left_grid_pin_40_[0] , 
        top_right_grid_pin_1_[0] , chany_bottom_in[2] , chany_bottom_in[12] , 
        chanx_left_in[0] , chanx_left_in[7] , chanx_left_in[14] } ) ,
    .sram ( mux_tree_tapbuf_size10_0_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size10_0_sram_inv ) , 
    .out ( chany_top_out[0] ) , .p0 ( optlc_net_123 ) ) ;
mux_tree_tapbuf_size10_0_1 mux_bottom_track_1 (
    .in ( { chany_top_in[2] , chany_top_in[12] , bottom_right_grid_pin_1_[0] , 
        bottom_left_grid_pin_35_[0] , bottom_left_grid_pin_37_[0] , 
        bottom_left_grid_pin_39_[0] , bottom_left_grid_pin_41_[0] , 
        chanx_left_in[1] , chanx_left_in[8] , chanx_left_in[15] } ) ,
    .sram ( mux_tree_tapbuf_size10_1_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size10_1_sram_inv ) , 
    .out ( chany_bottom_out[0] ) , .p0 ( optlc_net_124 ) ) ;
mux_tree_tapbuf_size10_mem_11 mem_top_track_0 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( ccff_head ) , 
    .ccff_tail ( mux_tree_tapbuf_size10_mem_0_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size10_0_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size10_0_sram_inv ) ) ;
mux_tree_tapbuf_size10_mem_0_1 mem_bottom_track_1 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size6_mem_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size10_mem_1_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size10_1_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size10_1_sram_inv ) ) ;
mux_tree_tapbuf_size8_1_1 mux_top_track_2 (
    .in ( { top_left_grid_pin_35_[0] , top_left_grid_pin_37_[0] , 
        top_left_grid_pin_39_[0] , top_left_grid_pin_41_[0] , 
        chany_bottom_in[4] , chany_bottom_in[13] , chanx_left_in[6] , 
        chanx_left_in[13] } ) ,
    .sram ( mux_tree_tapbuf_size8_0_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size8_0_sram_inv ) , 
    .out ( chany_top_out[1] ) , .p0 ( optlc_net_123 ) ) ;
mux_tree_tapbuf_size8_3 mux_top_track_8 (
    .in ( { top_left_grid_pin_34_[0] , top_left_grid_pin_38_[0] , 
        top_right_grid_pin_1_[0] , chany_bottom_in[6] , chany_bottom_in[16] , 
        chanx_left_in[4] , chanx_left_in[11] , chanx_left_in[18] } ) ,
    .sram ( mux_tree_tapbuf_size8_1_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size8_1_sram_inv ) , 
    .out ( chany_top_out[4] ) , .p0 ( optlc_net_125 ) ) ;
mux_tree_tapbuf_size8_0_1 mux_bottom_track_9 (
    .in ( { chany_top_in[6] , chany_top_in[16] , bottom_right_grid_pin_1_[0] , 
        bottom_left_grid_pin_37_[0] , bottom_left_grid_pin_41_[0] , 
        chanx_left_in[4] , chanx_left_in[11] , chanx_left_in[18] } ) ,
    .sram ( mux_tree_tapbuf_size8_2_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size8_2_sram_inv ) , 
    .out ( chany_bottom_out[4] ) , .p0 ( optlc_net_122 ) ) ;
mux_tree_tapbuf_size8_mem_1_1 mem_top_track_2 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size10_mem_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size8_mem_0_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size8_0_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size8_0_sram_inv ) ) ;
mux_tree_tapbuf_size8_mem_3 mem_top_track_8 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size14_mem_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size8_mem_1_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size8_1_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size8_1_sram_inv ) ) ;
mux_tree_tapbuf_size8_mem_0_1 mem_bottom_track_9 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size14_mem_1_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size8_mem_2_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size8_2_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size8_2_sram_inv ) ) ;
mux_tree_tapbuf_size14_1 mux_top_track_4 (
    .in ( { top_left_grid_pin_34_[0] , top_left_grid_pin_35_[0] , 
        top_left_grid_pin_36_[0] , top_left_grid_pin_37_[0] , 
        top_left_grid_pin_38_[0] , top_left_grid_pin_39_[0] , 
        top_left_grid_pin_40_[0] , top_left_grid_pin_41_[0] , 
        top_right_grid_pin_1_[0] , chany_bottom_in[5] , chany_bottom_in[14] , 
        chanx_left_in[5] , chanx_left_in[12] , chanx_left_in[19] } ) ,
    .sram ( mux_tree_tapbuf_size14_0_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size14_0_sram_inv ) , 
    .out ( chany_top_out[2] ) , .p0 ( optlc_net_125 ) ) ;
mux_tree_tapbuf_size14_0_1 mux_bottom_track_5 (
    .in ( { chany_top_in[5] , chany_top_in[14] , bottom_right_grid_pin_1_[0] , 
        bottom_left_grid_pin_34_[0] , bottom_left_grid_pin_35_[0] , 
        bottom_left_grid_pin_36_[0] , bottom_left_grid_pin_37_[0] , 
        bottom_left_grid_pin_38_[0] , bottom_left_grid_pin_39_[0] , 
        bottom_left_grid_pin_40_[0] , bottom_left_grid_pin_41_[0] , 
        chanx_left_in[3] , chanx_left_in[10] , chanx_left_in[17] } ) ,
    .sram ( mux_tree_tapbuf_size14_1_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size14_1_sram_inv ) , 
    .out ( chany_bottom_out[2] ) , .p0 ( optlc_net_122 ) ) ;
mux_tree_tapbuf_size14_mem_1 mem_top_track_4 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size8_mem_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size14_mem_0_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size14_0_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size14_0_sram_inv ) ) ;
mux_tree_tapbuf_size14_mem_0_1 mem_bottom_track_5 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size9_mem_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size14_mem_1_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size14_1_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size14_1_sram_inv ) ) ;
mux_tree_tapbuf_size7_5_1 mux_top_track_16 (
    .in ( { top_left_grid_pin_35_[0] , top_left_grid_pin_39_[0] , 
        chany_bottom_in[8] , chany_bottom_in[17] , chanx_left_in[3] , 
        chanx_left_in[10] , chanx_left_in[17] } ) ,
    .sram ( mux_tree_tapbuf_size7_0_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size7_0_sram_inv ) , 
    .out ( chany_top_out[8] ) , .p0 ( optlc_net_123 ) ) ;
mux_tree_tapbuf_size7_8 mux_top_track_24 (
    .in ( { top_left_grid_pin_36_[0] , top_left_grid_pin_40_[0] , 
        chany_bottom_in[9] , chany_bottom_in[18] , chanx_left_in[2] , 
        chanx_left_in[9] , chanx_left_in[16] } ) ,
    .sram ( mux_tree_tapbuf_size7_1_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size7_1_sram_inv ) , 
    .out ( chany_top_out[12] ) , .p0 ( optlc_net_123 ) ) ;
mux_tree_tapbuf_size7_0_4 mux_bottom_track_17 (
    .in ( { chany_top_in[8] , chany_top_in[17] , bottom_left_grid_pin_34_[0] , 
        bottom_left_grid_pin_38_[0] , chanx_left_in[5] , chanx_left_in[12] , 
        chanx_left_in[19] } ) ,
    .sram ( mux_tree_tapbuf_size7_2_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size7_2_sram_inv ) , 
    .out ( chany_bottom_out[8] ) , .p0 ( optlc_net_122 ) ) ;
mux_tree_tapbuf_size7_1_4 mux_left_track_1 (
    .in ( { chany_top_in[0] , chany_top_in[2] , chany_bottom_in[2] , 
        left_top_grid_pin_42_[0] , left_top_grid_pin_44_[0] , 
        left_top_grid_pin_46_[0] , left_top_grid_pin_48_[0] } ) ,
    .sram ( mux_tree_tapbuf_size7_3_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size7_3_sram_inv ) , 
    .out ( chanx_left_out[0] ) , .p0 ( optlc_net_125 ) ) ;
mux_tree_tapbuf_size7_2_3 mux_left_track_3 (
    .in ( { chany_top_in[4] , chany_bottom_in[0] , chany_bottom_in[4] , 
        left_top_grid_pin_43_[0] , left_top_grid_pin_45_[0] , 
        left_top_grid_pin_47_[0] , left_top_grid_pin_49_[0] } ) ,
    .sram ( mux_tree_tapbuf_size7_4_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size7_4_sram_inv ) , 
    .out ( chanx_left_out[1] ) , .p0 ( optlc_net_125 ) ) ;
mux_tree_tapbuf_size7_3_1 mux_left_track_5 (
    .in ( { chany_top_in[5] , chany_bottom_in[1] , chany_bottom_in[5] , 
        left_top_grid_pin_42_[0] , left_top_grid_pin_44_[0] , 
        left_top_grid_pin_46_[0] , left_top_grid_pin_48_[0] } ) ,
    .sram ( mux_tree_tapbuf_size7_5_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size7_5_sram_inv ) , 
    .out ( chanx_left_out[2] ) , .p0 ( optlc_net_125 ) ) ;
mux_tree_tapbuf_size7_4_1 mux_left_track_7 (
    .in ( { chany_top_in[6] , chany_bottom_in[3] , chany_bottom_in[6] , 
        left_top_grid_pin_43_[0] , left_top_grid_pin_45_[0] , 
        left_top_grid_pin_47_[0] , left_top_grid_pin_49_[0] } ) ,
    .sram ( mux_tree_tapbuf_size7_6_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size7_6_sram_inv ) , 
    .out ( chanx_left_out[3] ) , .p0 ( optlc_net_125 ) ) ;
mux_tree_tapbuf_size7_mem_5_1 mem_top_track_16 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size8_mem_1_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size7_mem_0_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size7_0_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size7_0_sram_inv ) ) ;
mux_tree_tapbuf_size7_mem_8 mem_top_track_24 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size7_mem_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size7_mem_1_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size7_1_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size7_1_sram_inv ) ) ;
mux_tree_tapbuf_size7_mem_0_4 mem_bottom_track_17 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size8_mem_2_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size7_mem_2_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size7_2_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size7_2_sram_inv ) ) ;
mux_tree_tapbuf_size7_mem_1_4 mem_left_track_1 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size6_mem_2_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size7_mem_3_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size7_3_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size7_3_sram_inv ) ) ;
mux_tree_tapbuf_size7_mem_2_3 mem_left_track_3 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size7_mem_3_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size7_mem_4_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size7_4_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size7_4_sram_inv ) ) ;
mux_tree_tapbuf_size7_mem_3_1 mem_left_track_5 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size7_mem_4_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size7_mem_5_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size7_5_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size7_5_sram_inv ) ) ;
mux_tree_tapbuf_size7_mem_4_1 mem_left_track_7 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size7_mem_5_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size7_mem_6_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size7_6_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size7_6_sram_inv ) ) ;
mux_tree_tapbuf_size6_9 mux_top_track_32 (
    .in ( { top_left_grid_pin_37_[0] , top_left_grid_pin_41_[0] , 
        chany_bottom_in[10] , chanx_left_in[1] , chanx_left_in[8] , 
        chanx_left_in[15] } ) ,
    .sram ( mux_tree_tapbuf_size6_0_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size6_0_sram_inv ) , 
    .out ( chany_top_out[16] ) , .p0 ( optlc_net_123 ) ) ;
mux_tree_tapbuf_size6_0_5 mux_bottom_track_25 (
    .in ( { chany_top_in[9] , chany_top_in[18] , bottom_left_grid_pin_35_[0] , 
        bottom_left_grid_pin_39_[0] , chanx_left_in[6] , chanx_left_in[13] } ) ,
    .sram ( mux_tree_tapbuf_size6_1_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size6_1_sram_inv ) , 
    .out ( chany_bottom_out[12] ) , .p0 ( optlc_net_122 ) ) ;
mux_tree_tapbuf_size6_1_3 mux_bottom_track_33 (
    .in ( { chany_top_in[10] , bottom_left_grid_pin_36_[0] , 
        bottom_left_grid_pin_40_[0] , chanx_left_in[0] , chanx_left_in[7] , 
        chanx_left_in[14] } ) ,
    .sram ( mux_tree_tapbuf_size6_2_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size6_2_sram_inv ) , 
    .out ( chany_bottom_out[16] ) , .p0 ( optlc_net_123 ) ) ;
mux_tree_tapbuf_size6_mem_9 mem_top_track_32 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size7_mem_1_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size6_mem_0_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size6_0_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size6_0_sram_inv ) ) ;
mux_tree_tapbuf_size6_mem_0_5 mem_bottom_track_25 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size7_mem_2_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size6_mem_1_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size6_1_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size6_1_sram_inv ) ) ;
mux_tree_tapbuf_size6_mem_1_3 mem_bottom_track_33 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size6_mem_1_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size6_mem_2_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size6_2_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size6_2_sram_inv ) ) ;
mux_tree_tapbuf_size9_1 mux_bottom_track_3 (
    .in ( { chany_top_in[4] , chany_top_in[13] , bottom_left_grid_pin_34_[0] , 
        bottom_left_grid_pin_36_[0] , bottom_left_grid_pin_38_[0] , 
        bottom_left_grid_pin_40_[0] , chanx_left_in[2] , chanx_left_in[9] , 
        chanx_left_in[16] } ) ,
    .sram ( mux_tree_tapbuf_size9_0_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size9_0_sram_inv ) ,
    .out ( { ropt_net_130 } ) ,
    .p0 ( optlc_net_124 ) ) ;
mux_tree_tapbuf_size9_mem_1 mem_bottom_track_3 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size10_mem_1_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size9_mem_0_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size9_0_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size9_0_sram_inv ) ) ;
mux_tree_tapbuf_size4_8 mux_left_track_9 (
    .in ( { chany_top_in[8] , chany_bottom_in[7] , chany_bottom_in[8] , 
        left_top_grid_pin_42_[0] } ) ,
    .sram ( mux_tree_tapbuf_size4_0_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size4_0_sram_inv ) , 
    .out ( chanx_left_out[4] ) , .p0 ( optlc_net_125 ) ) ;
mux_tree_tapbuf_size4_0_3 mux_left_track_11 (
    .in ( { chany_top_in[9] , chany_bottom_in[9] , chany_bottom_in[11] , 
        left_top_grid_pin_43_[0] } ) ,
    .sram ( mux_tree_tapbuf_size4_1_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size4_1_sram_inv ) ,
    .out ( { ropt_net_129 } ) ,
    .p0 ( optlc_net_122 ) ) ;
mux_tree_tapbuf_size4_1_2 mux_left_track_13 (
    .in ( { chany_top_in[10] , chany_bottom_in[10] , chany_bottom_in[15] , 
        left_top_grid_pin_44_[0] } ) ,
    .sram ( mux_tree_tapbuf_size4_2_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size4_2_sram_inv ) , 
    .out ( chanx_left_out[6] ) , .p0 ( optlc_net_122 ) ) ;
mux_tree_tapbuf_size4_2_2 mux_left_track_15 (
    .in ( { chany_top_in[12] , chany_bottom_in[12] , chany_bottom_in[19] , 
        left_top_grid_pin_45_[0] } ) ,
    .sram ( mux_tree_tapbuf_size4_3_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size4_3_sram_inv ) , 
    .out ( chanx_left_out[7] ) , .p0 ( optlc_net_123 ) ) ;
mux_tree_tapbuf_size4_mem_8 mem_left_track_9 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size7_mem_6_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size4_mem_0_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size4_0_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size4_0_sram_inv ) ) ;
mux_tree_tapbuf_size4_mem_0_3 mem_left_track_11 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size4_mem_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size4_mem_1_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size4_1_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size4_1_sram_inv ) ) ;
mux_tree_tapbuf_size4_mem_1_2 mem_left_track_13 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size4_mem_1_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size4_mem_2_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size4_2_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size4_2_sram_inv ) ) ;
mux_tree_tapbuf_size4_mem_2_2 mem_left_track_15 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size4_mem_2_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size4_mem_3_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size4_3_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size4_3_sram_inv ) ) ;
mux_tree_tapbuf_size3_0_5 mux_left_track_17 (
    .in ( { chany_top_in[13] , chany_bottom_in[13] , 
        left_top_grid_pin_46_[0] } ) ,
    .sram ( mux_tree_tapbuf_size3_0_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size3_0_sram_inv ) , 
    .out ( chanx_left_out[8] ) , .p0 ( optlc_net_125 ) ) ;
mux_tree_tapbuf_size3_1_4 mux_left_track_19 (
    .in ( { chany_top_in[14] , chany_bottom_in[14] , 
        left_top_grid_pin_47_[0] } ) ,
    .sram ( mux_tree_tapbuf_size3_1_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size3_1_sram_inv ) , 
    .out ( chanx_left_out[9] ) , .p0 ( optlc_net_125 ) ) ;
mux_tree_tapbuf_size3_2_4 mux_left_track_21 (
    .in ( { chany_top_in[16] , chany_bottom_in[16] , 
        left_top_grid_pin_48_[0] } ) ,
    .sram ( mux_tree_tapbuf_size3_2_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size3_2_sram_inv ) , 
    .out ( chanx_left_out[10] ) , .p0 ( optlc_net_125 ) ) ;
mux_tree_tapbuf_size3_3_3 mux_left_track_23 (
    .in ( { chany_top_in[17] , chany_bottom_in[17] , 
        left_top_grid_pin_49_[0] } ) ,
    .sram ( mux_tree_tapbuf_size3_3_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size3_3_sram_inv ) , 
    .out ( chanx_left_out[11] ) , .p0 ( optlc_net_123 ) ) ;
mux_tree_tapbuf_size3_10 mux_left_track_25 (
    .in ( { chany_top_in[18] , chany_bottom_in[18] , 
        left_top_grid_pin_42_[0] } ) ,
    .sram ( mux_tree_tapbuf_size3_4_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size3_4_sram_inv ) , 
    .out ( chanx_left_out[12] ) , .p0 ( optlc_net_123 ) ) ;
mux_tree_tapbuf_size3_mem_0_5 mem_left_track_17 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size4_mem_3_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size3_mem_0_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size3_0_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size3_0_sram_inv ) ) ;
mux_tree_tapbuf_size3_mem_1_4 mem_left_track_19 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size3_mem_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size3_mem_1_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size3_1_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size3_1_sram_inv ) ) ;
mux_tree_tapbuf_size3_mem_2_4 mem_left_track_21 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size3_mem_1_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size3_mem_2_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size3_2_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size3_2_sram_inv ) ) ;
mux_tree_tapbuf_size3_mem_3_3 mem_left_track_23 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size3_mem_2_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size3_mem_3_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size3_3_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size3_3_sram_inv ) ) ;
mux_tree_tapbuf_size3_mem_10 mem_left_track_25 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size3_mem_3_ccff_tail ) ,
    .ccff_tail ( { ropt_net_127 } ) ,
    .mem_out ( mux_tree_tapbuf_size3_4_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size3_4_sram_inv ) ) ;
sky130_fd_sc_hd__conb_1 optlc_111 ( .LO ( SYNOPSYS_UNCONNECTED_1 ) , 
    .HI ( optlc_net_122 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_113 ( .LO ( SYNOPSYS_UNCONNECTED_2 ) , 
    .HI ( optlc_net_123 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_758 ( .A ( ropt_net_154 ) , 
    .X ( chany_bottom_out[3] ) ) ;
sky130_fd_sc_hd__conb_1 optlc_115 ( .LO ( SYNOPSYS_UNCONNECTED_3 ) , 
    .HI ( optlc_net_124 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_5__4 ( .A ( chany_top_in[5] ) , 
    .X ( ropt_net_146 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_117 ( .LO ( SYNOPSYS_UNCONNECTED_4 ) , 
    .HI ( optlc_net_125 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_760 ( .A ( ropt_net_155 ) , 
    .X ( chany_top_out[15] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_761 ( .A ( ropt_net_156 ) , 
    .X ( chany_top_out[19] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_719 ( .A ( ropt_net_126 ) , 
    .X ( ropt_net_164 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_720 ( .A ( ropt_net_127 ) , 
    .X ( ropt_net_170 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_721 ( .A ( chany_top_in[1] ) , 
    .X ( chanx_left_out[19] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_12__11 ( .A ( chany_top_in[12] ) , 
    .X ( ropt_net_150 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_722 ( .A ( ropt_net_129 ) , 
    .X ( ropt_net_169 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_14__13 ( .A ( chany_top_in[14] ) , 
    .X ( chany_bottom_out[15] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_15__14 ( .A ( chany_top_in[15] ) , 
    .X ( ropt_net_167 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_16__15 ( .A ( chany_top_in[16] ) , 
    .X ( chany_bottom_out[17] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_723 ( .A ( ropt_net_130 ) , 
    .X ( chany_bottom_out[1] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_18__17 ( .A ( chany_top_in[18] ) , 
    .X ( ropt_net_138 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_765 ( .A ( ropt_net_157 ) , 
    .X ( chany_top_out[3] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_724 ( .A ( chany_top_in[4] ) , 
    .X ( chany_bottom_out[5] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_21__20 ( .A ( chany_bottom_in[4] ) , 
    .X ( ropt_net_141 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_725 ( .A ( chany_top_in[13] ) , 
    .X ( ropt_net_160 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_726 ( 
    .A ( chany_bottom_in[13] ) , .X ( chany_top_out[14] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_24__23 ( .A ( chany_bottom_in[8] ) , 
    .X ( ropt_net_148 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_727 ( .A ( chany_top_in[8] ) , 
    .X ( chany_bottom_out[9] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_728 ( .A ( chany_top_in[3] ) , 
    .X ( ropt_net_159 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_27__26 ( .A ( chany_bottom_in[12] ) , 
    .X ( ropt_net_149 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_729 ( .A ( ropt_net_136 ) , 
    .X ( ropt_net_158 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_730 ( 
    .A ( chany_bottom_in[16] ) , .X ( chany_top_out[17] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_731 ( .A ( ropt_net_138 ) , 
    .X ( chany_bottom_out[19] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_732 ( .A ( chany_top_in[19] ) , 
    .X ( ropt_net_171 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_32__31 ( .A ( chany_bottom_in[18] ) , 
    .X ( ropt_net_147 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_33__32 ( .A ( left_top_grid_pin_43_[0] ) , 
    .X ( chanx_left_out[13] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_766 ( .A ( ropt_net_158 ) , 
    .X ( chany_bottom_out[10] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_767 ( .A ( ropt_net_159 ) , 
    .X ( chanx_left_out[18] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_67 ( .A ( chany_top_in[7] ) , 
    .X ( ropt_net_126 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_68 ( .A ( chany_top_in[9] ) , 
    .X ( ropt_net_136 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_734 ( .A ( ropt_net_140 ) , 
    .X ( ropt_net_155 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_70 ( .A ( chany_bottom_in[2] ) , 
    .X ( ropt_net_145 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_RR_71 ( .A ( chany_bottom_in[5] ) , 
    .X ( ropt_net_143 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_RR_72 ( .A ( chany_bottom_in[6] ) , 
    .X ( chany_top_out[7] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_73 ( .A ( chany_bottom_in[9] ) , 
    .X ( ropt_net_142 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_RR_74 ( .A ( chany_bottom_in[10] ) , 
    .X ( chany_top_out[11] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_768 ( .A ( ropt_net_160 ) , 
    .X ( chany_bottom_out[14] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_76 ( .A ( chany_bottom_in[14] ) , 
    .X ( ropt_net_140 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_770 ( .A ( ropt_net_161 ) , 
    .X ( chanx_left_out[16] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_RR_78 ( .A ( chany_bottom_in[17] ) , 
    .X ( chany_top_out[18] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_735 ( .A ( ropt_net_141 ) , 
    .X ( chany_top_out[5] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_736 ( .A ( ropt_net_142 ) , 
    .X ( ropt_net_162 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_737 ( .A ( ropt_net_143 ) , 
    .X ( chany_top_out[6] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_738 ( .A ( ropt_net_144 ) , 
    .X ( ropt_net_161 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_P_97 ( .A ( chany_top_in[2] ) , 
    .X ( ropt_net_153 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_P_98 ( .A ( chany_top_in[6] ) , 
    .X ( chany_bottom_out[7] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_P_99 ( .A ( chany_top_in[10] ) , 
    .X ( ropt_net_151 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_P_100 ( .A ( chany_top_in[11] ) , 
    .X ( ropt_net_144 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_772 ( .A ( ropt_net_162 ) , 
    .X ( chany_top_out[10] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_P_102 ( .A ( chany_top_in[17] ) , 
    .X ( ropt_net_152 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_739 ( .A ( ropt_net_145 ) , 
    .X ( ropt_net_157 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_775 ( .A ( ropt_net_163 ) , 
    .X ( chany_top_out[13] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_741 ( .A ( ropt_net_146 ) , 
    .X ( ropt_net_168 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_743 ( .A ( ropt_net_147 ) , 
    .X ( ropt_net_156 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_745 ( .A ( ropt_net_148 ) , 
    .X ( chany_top_out[9] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_746 ( .A ( ropt_net_149 ) , 
    .X ( ropt_net_163 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_750 ( .A ( ropt_net_150 ) , 
    .X ( chany_bottom_out[13] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_753 ( .A ( ropt_net_151 ) , 
    .X ( ropt_net_165 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_754 ( .A ( ropt_net_152 ) , 
    .X ( ropt_net_166 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_755 ( .A ( ropt_net_153 ) , 
    .X ( ropt_net_154 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_776 ( .A ( ropt_net_164 ) , 
    .X ( chanx_left_out[17] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_778 ( .A ( ropt_net_165 ) , 
    .X ( chany_bottom_out[11] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_779 ( .A ( ropt_net_166 ) , 
    .X ( chany_bottom_out[18] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_781 ( .A ( ropt_net_167 ) , 
    .X ( chanx_left_out[15] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_782 ( .A ( ropt_net_168 ) , 
    .X ( chany_bottom_out[6] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_783 ( .A ( ropt_net_169 ) , 
    .X ( chanx_left_out[5] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_784 ( .A ( ropt_net_170 ) , 
    .X ( ccff_tail[0] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_786 ( .A ( ropt_net_171 ) , 
    .X ( chanx_left_out[14] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_7_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_34__39 ( .A ( mem_out[1] ) , 
    .X ( net_net_49 ) ) ;
sky130_fd_sc_hd__dlygate4sd1_1 BUFT_RR_49 ( .A ( net_net_49 ) , 
    .X ( net_net_48 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_69 ( .A ( net_net_48 ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_6_2 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_33__38 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_5_3 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_32__37 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_4_3 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_31__36 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_3_4 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_30__35 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_2_4 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_29__34 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_1_4 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_28__33 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_0_4 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_27__32 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_21 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_26__31 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_20 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_25__30 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_19 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_24__29 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_18 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_23__28 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_17 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_22__27 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_16 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_21__26 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_15 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_20__25 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_14 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_19__24 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_13 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_18__23 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_12 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_17__22 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_11 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_16__21 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_10_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_15__20 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_9_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_14__19 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_8_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_13__18 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_37 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_7_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_37 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
endmodule


module const1_32_1 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_6_2 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_32_1 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
endmodule


module const1_31_2 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_5_3 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_31_2 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
endmodule


module const1_30_3 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_4_3 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_30_3 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
endmodule


module const1_29_3 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_3_4 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_29_3 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
endmodule


module const1_28_3 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_2_4 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_28_3 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
endmodule


module const1_27_3 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_1_4 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_27_3 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
endmodule


module const1_26_5 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_0_4 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_26_5 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
endmodule


module const1_25_5 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_21 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_25_5 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
endmodule


module const1_24_5 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_20 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_24_5 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
endmodule


module const1_23_5 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_19 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_23_5 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
endmodule


module const1_22_5 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_18 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_22_5 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
endmodule


module const1_21_5 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_17 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_21_5 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
endmodule


module const1_20_5 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_16 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_20_5 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
endmodule


module const1_19_5 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_15 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_19_5 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
endmodule


module const1_18_5 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_14 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_18_5 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
endmodule


module const1_17_5 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_13 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_17_5 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
endmodule


module const1_16_6 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_12 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_16_6 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
endmodule


module const1_15_6 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_11 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_15_6 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
endmodule


module const1_14_6 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_10_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_14_6 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
endmodule


module const1_13_6 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_9_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_13_6 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
endmodule


module const1_12_6 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_8_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_12_6 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
endmodule


module mux_tree_tapbuf_size3_mem_0_4 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_12__17 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size3_mem_1_3 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_11__16 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size3_mem_2_3 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_10__15 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size3_mem_9 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_9__14 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_11_6 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size3_0_4 ( in , sram , sram_inv , out , p0 ) ;
input  [0:2] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;

const1_11_6 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( p0 ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
endmodule


module const1_10_6 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size3_1_3 ( in , sram , sram_inv , out , p0 ) ;
input  [0:2] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;

const1_10_6 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( p0 ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
endmodule


module const1_9_6 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size3_2_3 ( in , sram , sram_inv , out , p0 ) ;
input  [0:2] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;

const1_9_6 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( p0 ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
endmodule


module const1_8_6 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size3_9 ( in , sram , sram_inv , out , p0 ) ;
input  [0:2] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;

const1_8_6 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( p0 ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_41 ( 
    .A ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .X ( BUF_net_41 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_P_65 ( .A ( BUF_net_41 ) , 
    .X ( out[0] ) ) ;
endmodule


module mux_tree_tapbuf_size5_mem_1_2 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_8__13 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size5_mem_0_3 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_7__12 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size5_mem_7 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_6__11 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size5_mem_2_2 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_5__10 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_7_6 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size5_1_2 ( in , sram , sram_inv , out , p0 ) ;
input  [0:4] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;

const1_7_6 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , .A1 ( in[4] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
endmodule


module const1_6_7 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size5_0_3 ( in , sram , sram_inv , out , p0 ) ;
input  [0:4] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;

const1_6_7 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , .A1 ( in[4] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
endmodule


module const1_5_7 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size5_7 ( in , sram , sram_inv , out , p0 ) ;
input  [0:4] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;

const1_5_7 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , .A1 ( in[4] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
endmodule


module const1_4_7 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size5_2_2 ( in , sram , sram_inv , out , p0 ) ;
input  [0:4] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;

const1_4_7 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , .A1 ( in[4] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
endmodule


module mux_tree_tapbuf_size6_mem_1_2 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_4__9 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size6_mem_0_4 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_3__8 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size6_mem_8 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_2__7 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size6_mem_2_2 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_1__6 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_3_7 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size6_1_2 ( in , sram , sram_inv , out , p0 ) ;
input  [0:5] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;

const1_3_7 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
endmodule


module const1_2_7 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size6_0_4 ( in , sram , sram_inv , out , p0 ) ;
input  [0:5] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;

const1_2_7 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
endmodule


module const1_1_7 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size6_8 ( in , sram , sram_inv , out , p0 ) ;
input  [0:5] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;

const1_1_7 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
endmodule


module const1_0_7 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size6_2_2 ( in , sram , sram_inv , out , p0 ) ;
input  [0:5] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;

const1_0_7 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_8 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , .X ( out[0] ) ) ;
endmodule


module sb_2__0_ ( prog_clk , chany_top_in , top_left_grid_pin_34_ , 
    top_left_grid_pin_35_ , top_left_grid_pin_36_ , top_left_grid_pin_37_ , 
    top_left_grid_pin_38_ , top_left_grid_pin_39_ , top_left_grid_pin_40_ , 
    top_left_grid_pin_41_ , top_right_grid_pin_1_ , chanx_left_in , 
    left_top_grid_pin_42_ , left_top_grid_pin_43_ , left_top_grid_pin_44_ , 
    left_top_grid_pin_45_ , left_top_grid_pin_46_ , left_top_grid_pin_47_ , 
    left_top_grid_pin_48_ , left_top_grid_pin_49_ , left_bottom_grid_pin_1_ , 
    ccff_head , chany_top_out , chanx_left_out , ccff_tail ) ;
input  [0:0] prog_clk ;
input  [0:19] chany_top_in ;
input  [0:0] top_left_grid_pin_34_ ;
input  [0:0] top_left_grid_pin_35_ ;
input  [0:0] top_left_grid_pin_36_ ;
input  [0:0] top_left_grid_pin_37_ ;
input  [0:0] top_left_grid_pin_38_ ;
input  [0:0] top_left_grid_pin_39_ ;
input  [0:0] top_left_grid_pin_40_ ;
input  [0:0] top_left_grid_pin_41_ ;
input  [0:0] top_right_grid_pin_1_ ;
input  [0:19] chanx_left_in ;
input  [0:0] left_top_grid_pin_42_ ;
input  [0:0] left_top_grid_pin_43_ ;
input  [0:0] left_top_grid_pin_44_ ;
input  [0:0] left_top_grid_pin_45_ ;
input  [0:0] left_top_grid_pin_46_ ;
input  [0:0] left_top_grid_pin_47_ ;
input  [0:0] left_top_grid_pin_48_ ;
input  [0:0] left_top_grid_pin_49_ ;
input  [0:0] left_bottom_grid_pin_1_ ;
input  [0:0] ccff_head ;
output [0:19] chany_top_out ;
output [0:19] chanx_left_out ;
output [0:0] ccff_tail ;

wire [0:1] mux_tree_tapbuf_size2_0_sram ;
wire [0:1] mux_tree_tapbuf_size2_0_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_10_sram ;
wire [0:1] mux_tree_tapbuf_size2_10_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_11_sram ;
wire [0:1] mux_tree_tapbuf_size2_11_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_12_sram ;
wire [0:1] mux_tree_tapbuf_size2_12_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_13_sram ;
wire [0:1] mux_tree_tapbuf_size2_13_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_14_sram ;
wire [0:1] mux_tree_tapbuf_size2_14_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_15_sram ;
wire [0:1] mux_tree_tapbuf_size2_15_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_16_sram ;
wire [0:1] mux_tree_tapbuf_size2_16_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_17_sram ;
wire [0:1] mux_tree_tapbuf_size2_17_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_18_sram ;
wire [0:1] mux_tree_tapbuf_size2_18_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_19_sram ;
wire [0:1] mux_tree_tapbuf_size2_19_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_1_sram ;
wire [0:1] mux_tree_tapbuf_size2_1_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_20_sram ;
wire [0:1] mux_tree_tapbuf_size2_20_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_21_sram ;
wire [0:1] mux_tree_tapbuf_size2_21_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_2_sram ;
wire [0:1] mux_tree_tapbuf_size2_2_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_3_sram ;
wire [0:1] mux_tree_tapbuf_size2_3_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_4_sram ;
wire [0:1] mux_tree_tapbuf_size2_4_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_5_sram ;
wire [0:1] mux_tree_tapbuf_size2_5_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_6_sram ;
wire [0:1] mux_tree_tapbuf_size2_6_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_7_sram ;
wire [0:1] mux_tree_tapbuf_size2_7_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_8_sram ;
wire [0:1] mux_tree_tapbuf_size2_8_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_9_sram ;
wire [0:1] mux_tree_tapbuf_size2_9_sram_inv ;
wire [0:0] mux_tree_tapbuf_size2_mem_0_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_10_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_11_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_12_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_13_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_14_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_15_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_16_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_17_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_18_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_19_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_1_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_20_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_2_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_3_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_4_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_5_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_6_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_7_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_8_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_9_ccff_tail ;
wire [0:1] mux_tree_tapbuf_size3_0_sram ;
wire [0:1] mux_tree_tapbuf_size3_0_sram_inv ;
wire [0:1] mux_tree_tapbuf_size3_1_sram ;
wire [0:1] mux_tree_tapbuf_size3_1_sram_inv ;
wire [0:1] mux_tree_tapbuf_size3_2_sram ;
wire [0:1] mux_tree_tapbuf_size3_2_sram_inv ;
wire [0:1] mux_tree_tapbuf_size3_3_sram ;
wire [0:1] mux_tree_tapbuf_size3_3_sram_inv ;
wire [0:0] mux_tree_tapbuf_size3_mem_0_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size3_mem_1_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size3_mem_2_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size3_mem_3_ccff_tail ;
wire [0:2] mux_tree_tapbuf_size5_0_sram ;
wire [0:2] mux_tree_tapbuf_size5_0_sram_inv ;
wire [0:2] mux_tree_tapbuf_size5_1_sram ;
wire [0:2] mux_tree_tapbuf_size5_1_sram_inv ;
wire [0:2] mux_tree_tapbuf_size5_2_sram ;
wire [0:2] mux_tree_tapbuf_size5_2_sram_inv ;
wire [0:2] mux_tree_tapbuf_size5_3_sram ;
wire [0:2] mux_tree_tapbuf_size5_3_sram_inv ;
wire [0:0] mux_tree_tapbuf_size5_mem_0_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size5_mem_1_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size5_mem_2_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size5_mem_3_ccff_tail ;
wire [0:2] mux_tree_tapbuf_size6_0_sram ;
wire [0:2] mux_tree_tapbuf_size6_0_sram_inv ;
wire [0:2] mux_tree_tapbuf_size6_1_sram ;
wire [0:2] mux_tree_tapbuf_size6_1_sram_inv ;
wire [0:2] mux_tree_tapbuf_size6_2_sram ;
wire [0:2] mux_tree_tapbuf_size6_2_sram_inv ;
wire [0:2] mux_tree_tapbuf_size6_3_sram ;
wire [0:2] mux_tree_tapbuf_size6_3_sram_inv ;
wire [0:0] mux_tree_tapbuf_size6_mem_0_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size6_mem_1_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size6_mem_2_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size6_mem_3_ccff_tail ;

mux_tree_tapbuf_size6_2_2 mux_top_track_0 (
    .in ( { top_left_grid_pin_34_[0] , top_left_grid_pin_36_[0] , 
        top_left_grid_pin_38_[0] , top_left_grid_pin_40_[0] , 
        top_right_grid_pin_1_[0] , chanx_left_in[0] } ) ,
    .sram ( mux_tree_tapbuf_size6_0_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size6_0_sram_inv ) , 
    .out ( chany_top_out[0] ) , .p0 ( optlc_net_81 ) ) ;
mux_tree_tapbuf_size6_8 mux_top_track_4 (
    .in ( { top_left_grid_pin_34_[0] , top_left_grid_pin_36_[0] , 
        top_left_grid_pin_38_[0] , top_left_grid_pin_40_[0] , 
        top_right_grid_pin_1_[0] , chanx_left_in[18] } ) ,
    .sram ( mux_tree_tapbuf_size6_1_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size6_1_sram_inv ) , 
    .out ( chany_top_out[2] ) , .p0 ( optlc_net_81 ) ) ;
mux_tree_tapbuf_size6_0_4 mux_left_track_1 (
    .in ( { chany_top_in[0] , left_top_grid_pin_42_[0] , 
        left_top_grid_pin_44_[0] , left_top_grid_pin_46_[0] , 
        left_top_grid_pin_48_[0] , left_bottom_grid_pin_1_[0] } ) ,
    .sram ( mux_tree_tapbuf_size6_2_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size6_2_sram_inv ) , 
    .out ( chanx_left_out[0] ) , .p0 ( optlc_net_78 ) ) ;
mux_tree_tapbuf_size6_1_2 mux_left_track_5 (
    .in ( { chany_top_in[18] , left_top_grid_pin_42_[0] , 
        left_top_grid_pin_44_[0] , left_top_grid_pin_46_[0] , 
        left_top_grid_pin_48_[0] , left_bottom_grid_pin_1_[0] } ) ,
    .sram ( mux_tree_tapbuf_size6_3_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size6_3_sram_inv ) , 
    .out ( chanx_left_out[2] ) , .p0 ( optlc_net_78 ) ) ;
mux_tree_tapbuf_size6_mem_2_2 mem_top_track_0 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( ccff_head ) , 
    .ccff_tail ( mux_tree_tapbuf_size6_mem_0_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size6_0_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size6_0_sram_inv ) ) ;
mux_tree_tapbuf_size6_mem_8 mem_top_track_4 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size5_mem_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size6_mem_1_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size6_1_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size6_1_sram_inv ) ) ;
mux_tree_tapbuf_size6_mem_0_4 mem_left_track_1 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_13_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size6_mem_2_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size6_2_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size6_2_sram_inv ) ) ;
mux_tree_tapbuf_size6_mem_1_2 mem_left_track_5 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size5_mem_2_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size6_mem_3_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size6_3_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size6_3_sram_inv ) ) ;
mux_tree_tapbuf_size5_2_2 mux_top_track_2 (
    .in ( { top_left_grid_pin_35_[0] , top_left_grid_pin_37_[0] , 
        top_left_grid_pin_39_[0] , top_left_grid_pin_41_[0] , 
        chanx_left_in[19] } ) ,
    .sram ( mux_tree_tapbuf_size5_0_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size5_0_sram_inv ) , 
    .out ( chany_top_out[1] ) , .p0 ( optlc_net_80 ) ) ;
mux_tree_tapbuf_size5_7 mux_top_track_6 (
    .in ( { top_left_grid_pin_35_[0] , top_left_grid_pin_37_[0] , 
        top_left_grid_pin_39_[0] , top_left_grid_pin_41_[0] , 
        chanx_left_in[17] } ) ,
    .sram ( mux_tree_tapbuf_size5_1_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size5_1_sram_inv ) , 
    .out ( chany_top_out[3] ) , .p0 ( optlc_net_81 ) ) ;
mux_tree_tapbuf_size5_0_3 mux_left_track_3 (
    .in ( { chany_top_in[19] , left_top_grid_pin_43_[0] , 
        left_top_grid_pin_45_[0] , left_top_grid_pin_47_[0] , 
        left_top_grid_pin_49_[0] } ) ,
    .sram ( mux_tree_tapbuf_size5_2_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size5_2_sram_inv ) , 
    .out ( chanx_left_out[1] ) , .p0 ( optlc_net_80 ) ) ;
mux_tree_tapbuf_size5_1_2 mux_left_track_7 (
    .in ( { chany_top_in[17] , left_top_grid_pin_43_[0] , 
        left_top_grid_pin_45_[0] , left_top_grid_pin_47_[0] , 
        left_top_grid_pin_49_[0] } ) ,
    .sram ( mux_tree_tapbuf_size5_3_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size5_3_sram_inv ) , 
    .out ( chanx_left_out[3] ) , .p0 ( optlc_net_80 ) ) ;
mux_tree_tapbuf_size5_mem_2_2 mem_top_track_2 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size6_mem_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size5_mem_0_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size5_0_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size5_0_sram_inv ) ) ;
mux_tree_tapbuf_size5_mem_7 mem_top_track_6 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size6_mem_1_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size5_mem_1_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size5_1_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size5_1_sram_inv ) ) ;
mux_tree_tapbuf_size5_mem_0_3 mem_left_track_3 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size6_mem_2_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size5_mem_2_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size5_2_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size5_2_sram_inv ) ) ;
mux_tree_tapbuf_size5_mem_1_2 mem_left_track_7 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size6_mem_3_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size5_mem_3_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size5_3_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size5_3_sram_inv ) ) ;
mux_tree_tapbuf_size3_9 mux_top_track_8 (
    .in ( { top_left_grid_pin_34_[0] , top_right_grid_pin_1_[0] , 
        chanx_left_in[16] } ) ,
    .sram ( mux_tree_tapbuf_size3_0_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size3_0_sram_inv ) ,
    .out ( { ropt_net_89 } ) ,
    .p0 ( optlc_net_81 ) ) ;
mux_tree_tapbuf_size3_2_3 mux_top_track_24 (
    .in ( { top_left_grid_pin_34_[0] , top_right_grid_pin_1_[0] , 
        chanx_left_in[8] } ) ,
    .sram ( mux_tree_tapbuf_size3_1_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size3_1_sram_inv ) , 
    .out ( chany_top_out[12] ) , .p0 ( optlc_net_79 ) ) ;
mux_tree_tapbuf_size3_1_3 mux_left_track_9 (
    .in ( { chany_top_in[16] , left_top_grid_pin_42_[0] , 
        left_bottom_grid_pin_1_[0] } ) ,
    .sram ( mux_tree_tapbuf_size3_2_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size3_2_sram_inv ) , 
    .out ( chanx_left_out[4] ) , .p0 ( optlc_net_78 ) ) ;
mux_tree_tapbuf_size3_0_4 mux_left_track_25 (
    .in ( { chany_top_in[8] , left_top_grid_pin_42_[0] , 
        left_bottom_grid_pin_1_[0] } ) ,
    .sram ( mux_tree_tapbuf_size3_3_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size3_3_sram_inv ) , 
    .out ( chanx_left_out[12] ) , .p0 ( optlc_net_81 ) ) ;
mux_tree_tapbuf_size3_mem_9 mem_top_track_8 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size5_mem_1_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size3_mem_0_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size3_0_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size3_0_sram_inv ) ) ;
mux_tree_tapbuf_size3_mem_2_3 mem_top_track_24 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_6_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size3_mem_1_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size3_1_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size3_1_sram_inv ) ) ;
mux_tree_tapbuf_size3_mem_1_3 mem_left_track_9 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size5_mem_3_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size3_mem_2_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size3_2_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size3_2_sram_inv ) ) ;
mux_tree_tapbuf_size3_mem_0_4 mem_left_track_25 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_20_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size3_mem_3_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size3_3_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size3_3_sram_inv ) ) ;
mux_tree_tapbuf_size2_8_1 mux_top_track_10 (
    .in ( { top_left_grid_pin_35_[0] , chanx_left_in[15] } ) ,
    .sram ( mux_tree_tapbuf_size2_0_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_0_sram_inv ) , 
    .out ( chany_top_out[5] ) , .p0 ( optlc_net_81 ) ) ;
mux_tree_tapbuf_size2_9_1 mux_top_track_12 (
    .in ( { top_left_grid_pin_36_[0] , chanx_left_in[14] } ) ,
    .sram ( mux_tree_tapbuf_size2_1_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_1_sram_inv ) , 
    .out ( chany_top_out[6] ) , .p0 ( optlc_net_81 ) ) ;
mux_tree_tapbuf_size2_10_1 mux_top_track_14 (
    .in ( { top_left_grid_pin_37_[0] , chanx_left_in[13] } ) ,
    .sram ( mux_tree_tapbuf_size2_2_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_2_sram_inv ) , 
    .out ( chany_top_out[7] ) , .p0 ( optlc_net_79 ) ) ;
mux_tree_tapbuf_size2_11 mux_top_track_16 (
    .in ( { top_left_grid_pin_38_[0] , chanx_left_in[12] } ) ,
    .sram ( mux_tree_tapbuf_size2_3_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_3_sram_inv ) , 
    .out ( chany_top_out[8] ) , .p0 ( optlc_net_79 ) ) ;
mux_tree_tapbuf_size2_12 mux_top_track_18 (
    .in ( { top_left_grid_pin_39_[0] , chanx_left_in[11] } ) ,
    .sram ( mux_tree_tapbuf_size2_4_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_4_sram_inv ) , 
    .out ( chany_top_out[9] ) , .p0 ( optlc_net_79 ) ) ;
mux_tree_tapbuf_size2_13 mux_top_track_20 (
    .in ( { top_left_grid_pin_40_[0] , chanx_left_in[10] } ) ,
    .sram ( mux_tree_tapbuf_size2_5_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_5_sram_inv ) , 
    .out ( chany_top_out[10] ) , .p0 ( optlc_net_79 ) ) ;
mux_tree_tapbuf_size2_14 mux_top_track_22 (
    .in ( { top_left_grid_pin_41_[0] , chanx_left_in[9] } ) ,
    .sram ( mux_tree_tapbuf_size2_6_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_6_sram_inv ) , 
    .out ( chany_top_out[11] ) , .p0 ( optlc_net_79 ) ) ;
mux_tree_tapbuf_size2_15 mux_top_track_26 (
    .in ( { top_left_grid_pin_35_[0] , chanx_left_in[7] } ) ,
    .sram ( mux_tree_tapbuf_size2_7_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_7_sram_inv ) , 
    .out ( chany_top_out[13] ) , .p0 ( optlc_net_80 ) ) ;
mux_tree_tapbuf_size2_16 mux_top_track_28 (
    .in ( { top_left_grid_pin_36_[0] , chanx_left_in[6] } ) ,
    .sram ( mux_tree_tapbuf_size2_8_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_8_sram_inv ) , 
    .out ( chany_top_out[14] ) , .p0 ( optlc_net_79 ) ) ;
mux_tree_tapbuf_size2_17 mux_top_track_30 (
    .in ( { top_left_grid_pin_37_[0] , chanx_left_in[5] } ) ,
    .sram ( mux_tree_tapbuf_size2_9_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_9_sram_inv ) , 
    .out ( chany_top_out[15] ) , .p0 ( optlc_net_79 ) ) ;
mux_tree_tapbuf_size2_18 mux_top_track_32 (
    .in ( { top_left_grid_pin_38_[0] , chanx_left_in[4] } ) ,
    .sram ( mux_tree_tapbuf_size2_10_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_10_sram_inv ) , 
    .out ( chany_top_out[16] ) , .p0 ( optlc_net_79 ) ) ;
mux_tree_tapbuf_size2_19 mux_top_track_34 (
    .in ( { top_left_grid_pin_39_[0] , chanx_left_in[3] } ) ,
    .sram ( mux_tree_tapbuf_size2_11_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_11_sram_inv ) , 
    .out ( chany_top_out[17] ) , .p0 ( optlc_net_79 ) ) ;
mux_tree_tapbuf_size2_20 mux_top_track_36 (
    .in ( { top_left_grid_pin_40_[0] , chanx_left_in[2] } ) ,
    .sram ( mux_tree_tapbuf_size2_12_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_12_sram_inv ) , 
    .out ( chany_top_out[18] ) , .p0 ( optlc_net_79 ) ) ;
mux_tree_tapbuf_size2_21 mux_top_track_38 (
    .in ( { top_left_grid_pin_41_[0] , chanx_left_in[1] } ) ,
    .sram ( mux_tree_tapbuf_size2_13_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_13_sram_inv ) , 
    .out ( chany_top_out[19] ) , .p0 ( optlc_net_79 ) ) ;
mux_tree_tapbuf_size2_0_4 mux_left_track_11 (
    .in ( { chany_top_in[15] , left_top_grid_pin_43_[0] } ) ,
    .sram ( mux_tree_tapbuf_size2_14_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_14_sram_inv ) , 
    .out ( chanx_left_out[5] ) , .p0 ( optlc_net_80 ) ) ;
mux_tree_tapbuf_size2_1_4 mux_left_track_13 (
    .in ( { chany_top_in[14] , left_top_grid_pin_44_[0] } ) ,
    .sram ( mux_tree_tapbuf_size2_15_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_15_sram_inv ) , 
    .out ( chanx_left_out[6] ) , .p0 ( optlc_net_80 ) ) ;
mux_tree_tapbuf_size2_2_4 mux_left_track_15 (
    .in ( { chany_top_in[13] , left_top_grid_pin_45_[0] } ) ,
    .sram ( mux_tree_tapbuf_size2_16_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_16_sram_inv ) , 
    .out ( chanx_left_out[7] ) , .p0 ( optlc_net_80 ) ) ;
mux_tree_tapbuf_size2_3_4 mux_left_track_17 (
    .in ( { chany_top_in[12] , left_top_grid_pin_46_[0] } ) ,
    .sram ( mux_tree_tapbuf_size2_17_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_17_sram_inv ) , 
    .out ( chanx_left_out[8] ) , .p0 ( optlc_net_80 ) ) ;
mux_tree_tapbuf_size2_4_3 mux_left_track_19 (
    .in ( { chany_top_in[11] , left_top_grid_pin_47_[0] } ) ,
    .sram ( mux_tree_tapbuf_size2_18_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_18_sram_inv ) , 
    .out ( chanx_left_out[9] ) , .p0 ( optlc_net_80 ) ) ;
mux_tree_tapbuf_size2_5_3 mux_left_track_21 (
    .in ( { chany_top_in[10] , left_top_grid_pin_48_[0] } ) ,
    .sram ( mux_tree_tapbuf_size2_19_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_19_sram_inv ) , 
    .out ( chanx_left_out[10] ) , .p0 ( optlc_net_78 ) ) ;
mux_tree_tapbuf_size2_6_2 mux_left_track_23 (
    .in ( { chany_top_in[9] , left_top_grid_pin_49_[0] } ) ,
    .sram ( mux_tree_tapbuf_size2_20_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_20_sram_inv ) , 
    .out ( chanx_left_out[11] ) , .p0 ( optlc_net_80 ) ) ;
mux_tree_tapbuf_size2_7_1 mux_left_track_27 (
    .in ( { chany_top_in[7] , left_top_grid_pin_43_[0] } ) ,
    .sram ( mux_tree_tapbuf_size2_21_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_21_sram_inv ) , 
    .out ( chanx_left_out[13] ) , .p0 ( optlc_net_80 ) ) ;
mux_tree_tapbuf_size2_mem_8_1 mem_top_track_10 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size3_mem_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_0_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_0_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_0_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem_9_1 mem_top_track_12 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_1_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_1_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_1_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem_10_1 mem_top_track_14 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_1_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_2_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_2_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_2_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem_11 mem_top_track_16 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_2_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_3_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_3_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_3_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem_12 mem_top_track_18 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_3_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_4_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_4_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_4_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem_13 mem_top_track_20 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_4_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_5_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_5_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_5_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem_14 mem_top_track_22 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_5_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_6_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_6_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_6_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem_15 mem_top_track_26 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size3_mem_1_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_7_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_7_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_7_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem_16 mem_top_track_28 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_7_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_8_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_8_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_8_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem_17 mem_top_track_30 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_8_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_9_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_9_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_9_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem_18 mem_top_track_32 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_9_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_10_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_10_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_10_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem_19 mem_top_track_34 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_10_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_11_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_11_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_11_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem_20 mem_top_track_36 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_11_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_12_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_12_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_12_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem_21 mem_top_track_38 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_12_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_13_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_13_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_13_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem_0_4 mem_left_track_11 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size3_mem_2_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_14_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_14_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_14_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem_1_4 mem_left_track_13 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_14_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_15_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_15_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_15_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem_2_4 mem_left_track_15 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_15_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_16_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_16_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_16_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem_3_4 mem_left_track_17 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_16_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_17_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_17_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_17_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem_4_3 mem_left_track_19 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_17_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_18_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_18_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_18_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem_5_3 mem_left_track_21 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_18_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_19_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_19_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_19_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem_6_2 mem_left_track_23 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_19_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_20_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_20_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_20_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem_7_1 mem_left_track_27 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size3_mem_3_ccff_tail ) ,
    .ccff_tail ( { ropt_net_88 } ) ,
    .mem_out ( mux_tree_tapbuf_size2_21_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_21_sram_inv ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_676 ( .A ( ropt_net_91 ) , 
    .X ( chanx_left_out[14] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_677 ( .A ( ropt_net_92 ) , 
    .X ( ccff_tail[0] ) ) ;
sky130_fd_sc_hd__conb_1 optlc_72 ( .LO ( SYNOPSYS_UNCONNECTED_1 ) , 
    .HI ( optlc_net_78 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_74 ( .LO ( SYNOPSYS_UNCONNECTED_2 ) , 
    .HI ( optlc_net_79 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_76 ( .LO ( SYNOPSYS_UNCONNECTED_3 ) , 
    .HI ( optlc_net_80 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_6__5 ( .A ( chany_top_in[6] ) , 
    .X ( ropt_net_90 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_678 ( .A ( ropt_net_93 ) , 
    .X ( chanx_left_out[15] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_679 ( .A ( ropt_net_94 ) , 
    .X ( chanx_left_out[18] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_680 ( .A ( ropt_net_95 ) , 
    .X ( chanx_left_out[17] ) ) ;
sky130_fd_sc_hd__conb_1 optlc_78 ( .LO ( SYNOPSYS_UNCONNECTED_4 ) , 
    .HI ( optlc_net_81 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_668 ( .A ( chany_top_in[5] ) , 
    .X ( ropt_net_93 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_669 ( .A ( ropt_net_84 ) , 
    .X ( chanx_left_out[16] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 BUFT_P_63 ( .A ( chany_top_in[1] ) , 
    .X ( ropt_net_85 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_670 ( .A ( ropt_net_85 ) , 
    .X ( chanx_left_out[19] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 BUFT_P_67 ( .A ( chany_top_in[4] ) , 
    .X ( ropt_net_84 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_671 ( .A ( chany_top_in[3] ) , 
    .X ( ropt_net_95 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_672 ( .A ( chany_top_in[2] ) , 
    .X ( ropt_net_94 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_673 ( .A ( ropt_net_88 ) , 
    .X ( ropt_net_92 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_674 ( .A ( ropt_net_89 ) , 
    .X ( chany_top_out[4] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_675 ( .A ( ropt_net_90 ) , 
    .X ( ropt_net_91 ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_14 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_34__59 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_5_2 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_33__58 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_4_2 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_32__57 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_3_3 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_31__56 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_2_3 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_30__55 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_1_3 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_29__54 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_0_3 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_28__53 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_36 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_14 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_36 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
endmodule


module const1_32 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_5_2 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_32 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
endmodule


module const1_31_1 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_4_2 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_31_1 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
endmodule


module const1_30_2 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_3_3 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_30_2 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
endmodule


module const1_29_2 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_2_3 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_29_2 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
endmodule


module const1_28_2 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_1_3 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;

const1_28_2 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_8 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , .X ( out[0] ) ) ;
endmodule


module const1_27_2 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_0_3 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_27_2 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_73 ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
endmodule


module mux_tree_tapbuf_size4_mem_7 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_27__52 ( .A ( mem_out[2] ) , 
    .X ( net_net_95 ) ) ;
sky130_fd_sc_hd__dlygate4sd1_1 BUFT_RR_95 ( .A ( net_net_95 ) , 
    .X ( net_net_94 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_RR_130 ( .A ( net_net_94 ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size4_mem_1_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_26__51 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size4_mem_0_2 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_25__50 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size4_mem_2_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_24__49 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_26_4 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size4_7 ( in , sram , sram_inv , out , p0 ) ;
input  [0:3] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;

const1_26_4 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( in[2] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , .A1 ( in[3] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
endmodule


module const1_25_4 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size4_1_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:3] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;

const1_25_4 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( in[2] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , .A1 ( in[3] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
endmodule


module const1_24_4 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size4_0_2 ( in , sram , sram_inv , out , p0 ) ;
input  [0:3] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;

const1_24_4 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( in[2] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , .A1 ( in[3] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_P_137 ( 
    .A ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .X ( out[0] ) ) ;
endmodule


module const1_23_4 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size4_2_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:3] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;

const1_23_4 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( in[2] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , .A1 ( in[3] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
endmodule


module mux_tree_tapbuf_size7_mem_7 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_23__48 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size7_mem_2_2 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_22__47 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size7_mem_1_3 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_21__46 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size7_mem_0_3 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_20__45 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_22_4 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size7_7 ( in , sram , sram_inv , out , p0 ) ;
input  [0:6] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;

const1_22_4 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_3_ ( .A0 ( p0 ) , .A1 ( in[6] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_69 ( 
    .A ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , .X ( BUF_net_69 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 BUFT_P_136 ( .A ( BUF_net_69 ) , 
    .X ( out[0] ) ) ;
endmodule


module const1_21_4 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size7_2_2 ( in , sram , sram_inv , out , p0 ) ;
input  [0:6] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;

const1_21_4 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_3_ ( .A0 ( p0 ) , .A1 ( in[6] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_68 ( 
    .A ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , .X ( BUF_net_68 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 BUFT_P_135 ( .A ( BUF_net_68 ) , 
    .X ( out[0] ) ) ;
endmodule


module const1_20_4 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size7_1_3 ( in , sram , sram_inv , out , p0 ) ;
input  [0:6] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;

const1_20_4 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_3_ ( .A0 ( p0 ) , .A1 ( in[6] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_8 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .S ( sram[2] ) , .X ( out[0] ) ) ;
endmodule


module const1_19_4 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size7_0_3 ( in , sram , sram_inv , out , p0 ) ;
input  [0:6] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;

const1_19_4 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_3_ ( .A0 ( p0 ) , .A1 ( in[6] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_P_133 ( 
    .A ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , .X ( out[0] ) ) ;
endmodule


module mux_tree_tapbuf_size3_mem_5_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_19__44 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size3_mem_4_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_18__43 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size3_mem_3_2 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_17__42 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size3_mem_2_2 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_16__41 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size3_mem_1_2 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_15__40 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size3_mem_0_3 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_14__39 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size3_mem_8 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_13__38 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_18_4 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size3_5_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:2] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;

const1_18_4 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( p0 ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
endmodule


module const1_17_4 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size3_4_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:2] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;

const1_17_4 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( p0 ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
endmodule


module const1_16_5 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size3_3_2 ( in , sram , sram_inv , out , p0 ) ;
input  [0:2] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;

const1_16_5 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( p0 ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
endmodule


module const1_15_5 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size3_2_2 ( in , sram , sram_inv , out , p0 ) ;
input  [0:2] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;

const1_15_5 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( p0 ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
endmodule


module const1_14_5 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size3_1_2 ( in , sram , sram_inv , out , p0 ) ;
input  [0:2] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;

const1_14_5 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( p0 ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
endmodule


module const1_13_5 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size3_0_3 ( in , sram , sram_inv , out , p0 ) ;
input  [0:2] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;

const1_13_5 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( p0 ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
endmodule


module const1_12_5 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size3_8 ( in , sram , sram_inv , out , p0 ) ;
input  [0:2] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;

const1_12_5 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( p0 ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
endmodule


module mux_tree_tapbuf_size5_mem_2_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_12__37 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size5_mem_1_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_11__36 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size5_mem_3_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_10__35 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size5_mem_0_2 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_9__34 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size5_mem_6 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_8__33 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size5_mem_4 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_7__32 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size5_mem_5 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_6__31 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_11_5 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size5_2_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:4] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;

const1_11_5 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , .A1 ( in[4] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
endmodule


module const1_10_5 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size5_1_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:4] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;

const1_10_5 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , .A1 ( in[4] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
endmodule


module const1_9_5 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size5_3_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:4] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;

const1_9_5 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , .A1 ( in[4] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
endmodule


module const1_8_5 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size5_0_2 ( in , sram , sram_inv , out , p0 ) ;
input  [0:4] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;

const1_8_5 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , .A1 ( in[4] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
endmodule


module const1_7_5 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size5_6 ( in , sram , sram_inv , out , p0 ) ;
input  [0:4] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;

const1_7_5 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , .A1 ( in[4] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
endmodule


module const1_6_6 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size5_4 ( in , sram , sram_inv , out , p0 ) ;
input  [0:4] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;

const1_6_6 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , .A1 ( in[4] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
endmodule


module const1_5_6 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size5_5 ( in , sram , sram_inv , out , p0 ) ;
input  [0:4] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;

const1_5_6 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , .A1 ( in[4] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_62 ( 
    .A ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .X ( out[0] ) ) ;
endmodule


module mux_tree_tapbuf_size6_mem_1_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_5__30 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size6_mem_0_3 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_4__29 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size6_mem_7 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_3__28 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size6_mem_3_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_2__27 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size6_mem_2_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_1__26 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_4_6 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size6_1_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:5] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;

const1_4_6 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
endmodule


module const1_3_6 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size6_0_3 ( in , sram , sram_inv , out , p0 ) ;
input  [0:5] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;

const1_3_6 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
endmodule


module const1_2_6 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size6_7 ( in , sram , sram_inv , out , p0 ) ;
input  [0:5] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;

const1_2_6 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_8 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , .X ( out[0] ) ) ;
endmodule


module const1_1_6 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size6_3_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:5] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;

const1_1_6 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_8 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , .X ( out[0] ) ) ;
endmodule


module const1_0_6 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size6_2_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:5] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;

const1_0_6 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
endmodule


module sb_1__2_ ( prog_clk , chanx_right_in , right_top_grid_pin_1_ , 
    chany_bottom_in , bottom_left_grid_pin_34_ , bottom_left_grid_pin_35_ , 
    bottom_left_grid_pin_36_ , bottom_left_grid_pin_37_ , 
    bottom_left_grid_pin_38_ , bottom_left_grid_pin_39_ , 
    bottom_left_grid_pin_40_ , bottom_left_grid_pin_41_ , chanx_left_in , 
    left_top_grid_pin_1_ , ccff_head , chanx_right_out , chany_bottom_out , 
    chanx_left_out , ccff_tail ) ;
input  [0:0] prog_clk ;
input  [0:19] chanx_right_in ;
input  [0:0] right_top_grid_pin_1_ ;
input  [0:19] chany_bottom_in ;
input  [0:0] bottom_left_grid_pin_34_ ;
input  [0:0] bottom_left_grid_pin_35_ ;
input  [0:0] bottom_left_grid_pin_36_ ;
input  [0:0] bottom_left_grid_pin_37_ ;
input  [0:0] bottom_left_grid_pin_38_ ;
input  [0:0] bottom_left_grid_pin_39_ ;
input  [0:0] bottom_left_grid_pin_40_ ;
input  [0:0] bottom_left_grid_pin_41_ ;
input  [0:19] chanx_left_in ;
input  [0:0] left_top_grid_pin_1_ ;
input  [0:0] ccff_head ;
output [0:19] chanx_right_out ;
output [0:19] chany_bottom_out ;
output [0:19] chanx_left_out ;
output [0:0] ccff_tail ;

wire [0:1] mux_tree_tapbuf_size2_0_sram ;
wire [0:1] mux_tree_tapbuf_size2_0_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_1_sram ;
wire [0:1] mux_tree_tapbuf_size2_1_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_2_sram ;
wire [0:1] mux_tree_tapbuf_size2_2_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_3_sram ;
wire [0:1] mux_tree_tapbuf_size2_3_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_4_sram ;
wire [0:1] mux_tree_tapbuf_size2_4_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_5_sram ;
wire [0:1] mux_tree_tapbuf_size2_5_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_6_sram ;
wire [0:1] mux_tree_tapbuf_size2_6_sram_inv ;
wire [0:0] mux_tree_tapbuf_size2_mem_0_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_1_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_2_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_3_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_4_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_5_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_6_ccff_tail ;
wire [0:1] mux_tree_tapbuf_size3_0_sram ;
wire [0:1] mux_tree_tapbuf_size3_0_sram_inv ;
wire [0:1] mux_tree_tapbuf_size3_1_sram ;
wire [0:1] mux_tree_tapbuf_size3_1_sram_inv ;
wire [0:1] mux_tree_tapbuf_size3_2_sram ;
wire [0:1] mux_tree_tapbuf_size3_2_sram_inv ;
wire [0:1] mux_tree_tapbuf_size3_3_sram ;
wire [0:1] mux_tree_tapbuf_size3_3_sram_inv ;
wire [0:1] mux_tree_tapbuf_size3_4_sram ;
wire [0:1] mux_tree_tapbuf_size3_4_sram_inv ;
wire [0:1] mux_tree_tapbuf_size3_5_sram ;
wire [0:1] mux_tree_tapbuf_size3_5_sram_inv ;
wire [0:1] mux_tree_tapbuf_size3_6_sram ;
wire [0:1] mux_tree_tapbuf_size3_6_sram_inv ;
wire [0:0] mux_tree_tapbuf_size3_mem_0_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size3_mem_1_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size3_mem_2_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size3_mem_3_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size3_mem_4_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size3_mem_5_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size3_mem_6_ccff_tail ;
wire [0:2] mux_tree_tapbuf_size4_0_sram ;
wire [0:2] mux_tree_tapbuf_size4_0_sram_inv ;
wire [0:2] mux_tree_tapbuf_size4_1_sram ;
wire [0:2] mux_tree_tapbuf_size4_1_sram_inv ;
wire [0:2] mux_tree_tapbuf_size4_2_sram ;
wire [0:2] mux_tree_tapbuf_size4_2_sram_inv ;
wire [0:2] mux_tree_tapbuf_size4_3_sram ;
wire [0:2] mux_tree_tapbuf_size4_3_sram_inv ;
wire [0:0] mux_tree_tapbuf_size4_mem_0_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size4_mem_1_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size4_mem_2_ccff_tail ;
wire [0:2] mux_tree_tapbuf_size5_0_sram ;
wire [0:2] mux_tree_tapbuf_size5_0_sram_inv ;
wire [0:2] mux_tree_tapbuf_size5_1_sram ;
wire [0:2] mux_tree_tapbuf_size5_1_sram_inv ;
wire [0:2] mux_tree_tapbuf_size5_2_sram ;
wire [0:2] mux_tree_tapbuf_size5_2_sram_inv ;
wire [0:2] mux_tree_tapbuf_size5_3_sram ;
wire [0:2] mux_tree_tapbuf_size5_3_sram_inv ;
wire [0:2] mux_tree_tapbuf_size5_4_sram ;
wire [0:2] mux_tree_tapbuf_size5_4_sram_inv ;
wire [0:2] mux_tree_tapbuf_size5_5_sram ;
wire [0:2] mux_tree_tapbuf_size5_5_sram_inv ;
wire [0:2] mux_tree_tapbuf_size5_6_sram ;
wire [0:2] mux_tree_tapbuf_size5_6_sram_inv ;
wire [0:0] mux_tree_tapbuf_size5_mem_0_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size5_mem_1_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size5_mem_2_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size5_mem_3_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size5_mem_4_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size5_mem_5_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size5_mem_6_ccff_tail ;
wire [0:2] mux_tree_tapbuf_size6_0_sram ;
wire [0:2] mux_tree_tapbuf_size6_0_sram_inv ;
wire [0:2] mux_tree_tapbuf_size6_1_sram ;
wire [0:2] mux_tree_tapbuf_size6_1_sram_inv ;
wire [0:2] mux_tree_tapbuf_size6_2_sram ;
wire [0:2] mux_tree_tapbuf_size6_2_sram_inv ;
wire [0:2] mux_tree_tapbuf_size6_3_sram ;
wire [0:2] mux_tree_tapbuf_size6_3_sram_inv ;
wire [0:2] mux_tree_tapbuf_size6_4_sram ;
wire [0:2] mux_tree_tapbuf_size6_4_sram_inv ;
wire [0:0] mux_tree_tapbuf_size6_mem_0_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size6_mem_1_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size6_mem_2_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size6_mem_3_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size6_mem_4_ccff_tail ;
wire [0:2] mux_tree_tapbuf_size7_0_sram ;
wire [0:2] mux_tree_tapbuf_size7_0_sram_inv ;
wire [0:2] mux_tree_tapbuf_size7_1_sram ;
wire [0:2] mux_tree_tapbuf_size7_1_sram_inv ;
wire [0:2] mux_tree_tapbuf_size7_2_sram ;
wire [0:2] mux_tree_tapbuf_size7_2_sram_inv ;
wire [0:2] mux_tree_tapbuf_size7_3_sram ;
wire [0:2] mux_tree_tapbuf_size7_3_sram_inv ;
wire [0:0] mux_tree_tapbuf_size7_mem_0_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size7_mem_1_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size7_mem_2_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size7_mem_3_ccff_tail ;

mux_tree_tapbuf_size6_2_1 mux_right_track_0 (
    .in ( { right_top_grid_pin_1_[0] , chany_bottom_in[5] , 
        chany_bottom_in[12] , chany_bottom_in[19] , chanx_left_in[2] , 
        chanx_left_in[12] } ) ,
    .sram ( mux_tree_tapbuf_size6_0_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size6_0_sram_inv ) , 
    .out ( chanx_right_out[0] ) , .p0 ( optlc_net_163 ) ) ;
mux_tree_tapbuf_size6_3_1 mux_right_track_4 (
    .in ( { right_top_grid_pin_1_[0] , chany_bottom_in[3] , 
        chany_bottom_in[10] , chany_bottom_in[17] , chanx_left_in[5] , 
        chanx_left_in[14] } ) ,
    .sram ( mux_tree_tapbuf_size6_1_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size6_1_sram_inv ) , 
    .out ( chanx_right_out[2] ) , .p0 ( optlc_net_163 ) ) ;
mux_tree_tapbuf_size6_7 mux_right_track_8 (
    .in ( { right_top_grid_pin_1_[0] , chany_bottom_in[2] , 
        chany_bottom_in[9] , chany_bottom_in[16] , chanx_left_in[6] , 
        chanx_left_in[16] } ) ,
    .sram ( mux_tree_tapbuf_size6_2_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size6_2_sram_inv ) , 
    .out ( chanx_right_out[4] ) , .p0 ( optlc_net_163 ) ) ;
mux_tree_tapbuf_size6_0_3 mux_left_track_5 (
    .in ( { chanx_right_in[5] , chanx_right_in[14] , chany_bottom_in[1] , 
        chany_bottom_in[8] , chany_bottom_in[15] , left_top_grid_pin_1_[0] } ) ,
    .sram ( mux_tree_tapbuf_size6_3_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size6_3_sram_inv ) , 
    .out ( chanx_left_out[2] ) , .p0 ( optlc_net_162 ) ) ;
mux_tree_tapbuf_size6_1_1 mux_left_track_9 (
    .in ( { chanx_right_in[6] , chanx_right_in[16] , chany_bottom_in[2] , 
        chany_bottom_in[9] , chany_bottom_in[16] , left_top_grid_pin_1_[0] } ) ,
    .sram ( mux_tree_tapbuf_size6_4_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size6_4_sram_inv ) , 
    .out ( chanx_left_out[4] ) , .p0 ( optlc_net_162 ) ) ;
mux_tree_tapbuf_size6_mem_2_1 mem_right_track_0 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( ccff_head ) , 
    .ccff_tail ( mux_tree_tapbuf_size6_mem_0_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size6_0_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size6_0_sram_inv ) ) ;
mux_tree_tapbuf_size6_mem_3_1 mem_right_track_4 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size5_mem_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size6_mem_1_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size6_1_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size6_1_sram_inv ) ) ;
mux_tree_tapbuf_size6_mem_7 mem_right_track_8 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size6_mem_1_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size6_mem_2_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size6_2_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size6_2_sram_inv ) ) ;
mux_tree_tapbuf_size6_mem_0_3 mem_left_track_5 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size5_mem_4_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size6_mem_3_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size6_3_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size6_3_sram_inv ) ) ;
mux_tree_tapbuf_size6_mem_1_1 mem_left_track_9 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size6_mem_3_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size6_mem_4_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size6_4_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size6_4_sram_inv ) ) ;
mux_tree_tapbuf_size5_5 mux_right_track_2 (
    .in ( { chany_bottom_in[4] , chany_bottom_in[11] , chany_bottom_in[18] , 
        chanx_left_in[4] , chanx_left_in[13] } ) ,
    .sram ( mux_tree_tapbuf_size5_0_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size5_0_sram_inv ) ,
    .out ( { ropt_net_172 } ) ,
    .p0 ( optlc_net_163 ) ) ;
mux_tree_tapbuf_size5_4 mux_right_track_16 (
    .in ( { chany_bottom_in[1] , chany_bottom_in[8] , chany_bottom_in[15] , 
        chanx_left_in[8] , chanx_left_in[17] } ) ,
    .sram ( mux_tree_tapbuf_size5_1_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size5_1_sram_inv ) , 
    .out ( chanx_right_out[8] ) , .p0 ( optlc_net_165 ) ) ;
mux_tree_tapbuf_size5_6 mux_right_track_24 (
    .in ( { chany_bottom_in[0] , chany_bottom_in[7] , chany_bottom_in[14] , 
        chanx_left_in[9] , chanx_left_in[18] } ) ,
    .sram ( mux_tree_tapbuf_size5_2_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size5_2_sram_inv ) , 
    .out ( chanx_right_out[12] ) , .p0 ( optlc_net_165 ) ) ;
mux_tree_tapbuf_size5_0_2 mux_left_track_1 (
    .in ( { chanx_right_in[2] , chanx_right_in[12] , chany_bottom_in[6] , 
        chany_bottom_in[13] , left_top_grid_pin_1_[0] } ) ,
    .sram ( mux_tree_tapbuf_size5_3_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size5_3_sram_inv ) , 
    .out ( chanx_left_out[0] ) , .p0 ( optlc_net_162 ) ) ;
mux_tree_tapbuf_size5_3_1 mux_left_track_3 (
    .in ( { chanx_right_in[4] , chanx_right_in[13] , chany_bottom_in[0] , 
        chany_bottom_in[7] , chany_bottom_in[14] } ) ,
    .sram ( mux_tree_tapbuf_size5_4_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size5_4_sram_inv ) , 
    .out ( chanx_left_out[1] ) , .p0 ( optlc_net_162 ) ) ;
mux_tree_tapbuf_size5_1_1 mux_left_track_17 (
    .in ( { chanx_right_in[8] , chanx_right_in[17] , chany_bottom_in[3] , 
        chany_bottom_in[10] , chany_bottom_in[17] } ) ,
    .sram ( mux_tree_tapbuf_size5_5_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size5_5_sram_inv ) , 
    .out ( chanx_left_out[8] ) , .p0 ( optlc_net_164 ) ) ;
mux_tree_tapbuf_size5_2_1 mux_left_track_25 (
    .in ( { chanx_right_in[9] , chanx_right_in[18] , chany_bottom_in[4] , 
        chany_bottom_in[11] , chany_bottom_in[18] } ) ,
    .sram ( mux_tree_tapbuf_size5_6_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size5_6_sram_inv ) , 
    .out ( chanx_left_out[12] ) , .p0 ( optlc_net_164 ) ) ;
mux_tree_tapbuf_size5_mem_5 mem_right_track_2 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size6_mem_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size5_mem_0_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size5_0_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size5_0_sram_inv ) ) ;
mux_tree_tapbuf_size5_mem_4 mem_right_track_16 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size6_mem_2_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size5_mem_1_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size5_1_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size5_1_sram_inv ) ) ;
mux_tree_tapbuf_size5_mem_6 mem_right_track_24 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size5_mem_1_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size5_mem_2_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size5_2_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size5_2_sram_inv ) ) ;
mux_tree_tapbuf_size5_mem_0_2 mem_left_track_1 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_6_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size5_mem_3_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size5_3_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size5_3_sram_inv ) ) ;
mux_tree_tapbuf_size5_mem_3_1 mem_left_track_3 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size5_mem_3_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size5_mem_4_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size5_4_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size5_4_sram_inv ) ) ;
mux_tree_tapbuf_size5_mem_1_1 mem_left_track_17 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size6_mem_4_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size5_mem_5_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size5_5_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size5_5_sram_inv ) ) ;
mux_tree_tapbuf_size5_mem_2_1 mem_left_track_25 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size5_mem_5_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size5_mem_6_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size5_6_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size5_6_sram_inv ) ) ;
mux_tree_tapbuf_size3_8 mux_right_track_32 (
    .in ( { chany_bottom_in[6] , chany_bottom_in[13] , chanx_left_in[10] } ) ,
    .sram ( mux_tree_tapbuf_size3_0_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size3_0_sram_inv ) , 
    .out ( chanx_right_out[16] ) , .p0 ( optlc_net_165 ) ) ;
mux_tree_tapbuf_size3_0_3 mux_bottom_track_13 (
    .in ( { chanx_right_in[10] , bottom_left_grid_pin_36_[0] , 
        chanx_left_in[10] } ) ,
    .sram ( mux_tree_tapbuf_size3_1_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size3_1_sram_inv ) , 
    .out ( chany_bottom_out[6] ) , .p0 ( optlc_net_164 ) ) ;
mux_tree_tapbuf_size3_1_2 mux_bottom_track_15 (
    .in ( { chanx_right_in[12] , bottom_left_grid_pin_37_[0] , 
        chanx_left_in[12] } ) ,
    .sram ( mux_tree_tapbuf_size3_2_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size3_2_sram_inv ) , 
    .out ( chany_bottom_out[7] ) , .p0 ( optlc_net_164 ) ) ;
mux_tree_tapbuf_size3_2_2 mux_bottom_track_17 (
    .in ( { chanx_right_in[13] , bottom_left_grid_pin_38_[0] , 
        chanx_left_in[13] } ) ,
    .sram ( mux_tree_tapbuf_size3_3_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size3_3_sram_inv ) , 
    .out ( chany_bottom_out[8] ) , .p0 ( optlc_net_163 ) ) ;
mux_tree_tapbuf_size3_3_2 mux_bottom_track_19 (
    .in ( { chanx_right_in[14] , bottom_left_grid_pin_39_[0] , 
        chanx_left_in[14] } ) ,
    .sram ( mux_tree_tapbuf_size3_4_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size3_4_sram_inv ) , 
    .out ( chany_bottom_out[9] ) , .p0 ( optlc_net_162 ) ) ;
mux_tree_tapbuf_size3_4_1 mux_bottom_track_21 (
    .in ( { chanx_right_in[16] , bottom_left_grid_pin_40_[0] , 
        chanx_left_in[16] } ) ,
    .sram ( mux_tree_tapbuf_size3_5_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size3_5_sram_inv ) , 
    .out ( chany_bottom_out[10] ) , .p0 ( optlc_net_162 ) ) ;
mux_tree_tapbuf_size3_5_1 mux_bottom_track_23 (
    .in ( { chanx_right_in[17] , bottom_left_grid_pin_41_[0] , 
        chanx_left_in[17] } ) ,
    .sram ( mux_tree_tapbuf_size3_6_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size3_6_sram_inv ) , 
    .out ( chany_bottom_out[11] ) , .p0 ( optlc_net_162 ) ) ;
mux_tree_tapbuf_size3_mem_8 mem_right_track_32 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size5_mem_2_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size3_mem_0_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size3_0_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size3_0_sram_inv ) ) ;
mux_tree_tapbuf_size3_mem_0_3 mem_bottom_track_13 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size4_mem_1_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size3_mem_1_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size3_1_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size3_1_sram_inv ) ) ;
mux_tree_tapbuf_size3_mem_1_2 mem_bottom_track_15 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size3_mem_1_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size3_mem_2_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size3_2_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size3_2_sram_inv ) ) ;
mux_tree_tapbuf_size3_mem_2_2 mem_bottom_track_17 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size3_mem_2_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size3_mem_3_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size3_3_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size3_3_sram_inv ) ) ;
mux_tree_tapbuf_size3_mem_3_2 mem_bottom_track_19 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size3_mem_3_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size3_mem_4_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size3_4_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size3_4_sram_inv ) ) ;
mux_tree_tapbuf_size3_mem_4_1 mem_bottom_track_21 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size3_mem_4_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size3_mem_5_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size3_5_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size3_5_sram_inv ) ) ;
mux_tree_tapbuf_size3_mem_5_1 mem_bottom_track_23 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size3_mem_5_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size3_mem_6_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size3_6_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size3_6_sram_inv ) ) ;
mux_tree_tapbuf_size7_0_3 mux_bottom_track_1 (
    .in ( { chanx_right_in[2] , bottom_left_grid_pin_34_[0] , 
        bottom_left_grid_pin_36_[0] , bottom_left_grid_pin_38_[0] , 
        bottom_left_grid_pin_40_[0] , chanx_left_in[1] , chanx_left_in[2] } ) ,
    .sram ( mux_tree_tapbuf_size7_0_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size7_0_sram_inv ) ,
    .out ( { ropt_net_175 } ) ,
    .p0 ( optlc_net_162 ) ) ;
mux_tree_tapbuf_size7_1_3 mux_bottom_track_3 (
    .in ( { chanx_right_in[4] , bottom_left_grid_pin_35_[0] , 
        bottom_left_grid_pin_37_[0] , bottom_left_grid_pin_39_[0] , 
        bottom_left_grid_pin_41_[0] , chanx_left_in[3] , chanx_left_in[4] } ) ,
    .sram ( mux_tree_tapbuf_size7_1_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size7_1_sram_inv ) , 
    .out ( chany_bottom_out[1] ) , .p0 ( optlc_net_164 ) ) ;
mux_tree_tapbuf_size7_2_2 mux_bottom_track_5 (
    .in ( { chanx_right_in[5] , bottom_left_grid_pin_34_[0] , 
        bottom_left_grid_pin_36_[0] , bottom_left_grid_pin_38_[0] , 
        bottom_left_grid_pin_40_[0] , chanx_left_in[5] , chanx_left_in[7] } ) ,
    .sram ( mux_tree_tapbuf_size7_2_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size7_2_sram_inv ) ,
    .out ( { ropt_net_207 } ) ,
    .p0 ( optlc_net_164 ) ) ;
mux_tree_tapbuf_size7_7 mux_bottom_track_7 (
    .in ( { chanx_right_in[6] , bottom_left_grid_pin_35_[0] , 
        bottom_left_grid_pin_37_[0] , bottom_left_grid_pin_39_[0] , 
        bottom_left_grid_pin_41_[0] , chanx_left_in[6] , chanx_left_in[11] } ) ,
    .sram ( mux_tree_tapbuf_size7_3_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size7_3_sram_inv ) , 
    .out ( chany_bottom_out[3] ) , .p0 ( optlc_net_164 ) ) ;
mux_tree_tapbuf_size7_mem_0_3 mem_bottom_track_1 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size3_mem_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size7_mem_0_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size7_0_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size7_0_sram_inv ) ) ;
mux_tree_tapbuf_size7_mem_1_3 mem_bottom_track_3 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size7_mem_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size7_mem_1_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size7_1_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size7_1_sram_inv ) ) ;
mux_tree_tapbuf_size7_mem_2_2 mem_bottom_track_5 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size7_mem_1_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size7_mem_2_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size7_2_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size7_2_sram_inv ) ) ;
mux_tree_tapbuf_size7_mem_7 mem_bottom_track_7 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size7_mem_2_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size7_mem_3_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size7_3_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size7_3_sram_inv ) ) ;
mux_tree_tapbuf_size4_2_1 mux_bottom_track_9 (
    .in ( { chanx_right_in[8] , bottom_left_grid_pin_34_[0] , 
        chanx_left_in[8] , chanx_left_in[15] } ) ,
    .sram ( mux_tree_tapbuf_size4_0_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size4_0_sram_inv ) , 
    .out ( chany_bottom_out[4] ) , .p0 ( optlc_net_164 ) ) ;
mux_tree_tapbuf_size4_0_2 mux_bottom_track_11 (
    .in ( { chanx_right_in[9] , bottom_left_grid_pin_35_[0] , 
        chanx_left_in[9] , chanx_left_in[19] } ) ,
    .sram ( mux_tree_tapbuf_size4_1_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size4_1_sram_inv ) ,
    .out ( { ropt_net_176 } ) ,
    .p0 ( optlc_net_164 ) ) ;
mux_tree_tapbuf_size4_1_1 mux_bottom_track_25 (
    .in ( { chanx_right_in[18] , chanx_right_in[19] , 
        bottom_left_grid_pin_34_[0] , chanx_left_in[18] } ) ,
    .sram ( mux_tree_tapbuf_size4_2_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size4_2_sram_inv ) , 
    .out ( chany_bottom_out[12] ) , .p0 ( optlc_net_165 ) ) ;
mux_tree_tapbuf_size4_7 mux_left_track_33 (
    .in ( { chanx_right_in[10] , chany_bottom_in[5] , chany_bottom_in[12] , 
        chany_bottom_in[19] } ) ,
    .sram ( mux_tree_tapbuf_size4_3_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size4_3_sram_inv ) , 
    .out ( chanx_left_out[16] ) , .p0 ( optlc_net_164 ) ) ;
mux_tree_tapbuf_size4_mem_2_1 mem_bottom_track_9 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size7_mem_3_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size4_mem_0_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size4_0_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size4_0_sram_inv ) ) ;
mux_tree_tapbuf_size4_mem_0_2 mem_bottom_track_11 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size4_mem_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size4_mem_1_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size4_1_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size4_1_sram_inv ) ) ;
mux_tree_tapbuf_size4_mem_1_1 mem_bottom_track_25 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size3_mem_6_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size4_mem_2_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size4_2_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size4_2_sram_inv ) ) ;
mux_tree_tapbuf_size4_mem_7 mem_left_track_33 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size5_mem_6_ccff_tail ) , 
    .ccff_tail ( ccff_tail ) , .mem_out ( mux_tree_tapbuf_size4_3_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size4_3_sram_inv ) ) ;
mux_tree_tapbuf_size2_0_3 mux_bottom_track_27 (
    .in ( { chanx_right_in[15] , bottom_left_grid_pin_35_[0] } ) ,
    .sram ( mux_tree_tapbuf_size2_0_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_0_sram_inv ) ,
    .out ( { ropt_net_169 } ) ,
    .p0 ( optlc_net_165 ) ) ;
mux_tree_tapbuf_size2_1_3 mux_bottom_track_29 (
    .in ( { chanx_right_in[11] , bottom_left_grid_pin_36_[0] } ) ,
    .sram ( mux_tree_tapbuf_size2_1_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_1_sram_inv ) , 
    .out ( chany_bottom_out[14] ) , .p0 ( optlc_net_165 ) ) ;
mux_tree_tapbuf_size2_2_3 mux_bottom_track_31 (
    .in ( { chanx_right_in[7] , bottom_left_grid_pin_37_[0] } ) ,
    .sram ( mux_tree_tapbuf_size2_2_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_2_sram_inv ) , 
    .out ( chany_bottom_out[15] ) , .p0 ( optlc_net_163 ) ) ;
mux_tree_tapbuf_size2_3_3 mux_bottom_track_33 (
    .in ( { chanx_right_in[3] , bottom_left_grid_pin_38_[0] } ) ,
    .sram ( mux_tree_tapbuf_size2_3_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_3_sram_inv ) , 
    .out ( chany_bottom_out[16] ) , .p0 ( optlc_net_163 ) ) ;
mux_tree_tapbuf_size2_4_2 mux_bottom_track_35 (
    .in ( { chanx_right_in[1] , bottom_left_grid_pin_39_[0] } ) ,
    .sram ( mux_tree_tapbuf_size2_4_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_4_sram_inv ) , 
    .out ( chany_bottom_out[17] ) , .p0 ( optlc_net_163 ) ) ;
mux_tree_tapbuf_size2_5_2 mux_bottom_track_37 (
    .in ( { chanx_right_in[0] , bottom_left_grid_pin_40_[0] } ) ,
    .sram ( mux_tree_tapbuf_size2_5_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_5_sram_inv ) , 
    .out ( chany_bottom_out[18] ) , .p0 ( optlc_net_162 ) ) ;
mux_tree_tapbuf_size2_14 mux_bottom_track_39 (
    .in ( { bottom_left_grid_pin_41_[0] , chanx_left_in[0] } ) ,
    .sram ( mux_tree_tapbuf_size2_6_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_6_sram_inv ) , 
    .out ( chany_bottom_out[19] ) , .p0 ( optlc_net_162 ) ) ;
mux_tree_tapbuf_size2_mem_0_3 mem_bottom_track_27 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size4_mem_2_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_0_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_0_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_0_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem_1_3 mem_bottom_track_29 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_1_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_1_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_1_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem_2_3 mem_bottom_track_31 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_1_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_2_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_2_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_2_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem_3_3 mem_bottom_track_33 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_2_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_3_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_3_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_3_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem_4_2 mem_bottom_track_35 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_3_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_4_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_4_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_4_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem_5_2 mem_bottom_track_37 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_4_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_5_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_5_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_5_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem_14 mem_bottom_track_39 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_5_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_6_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_6_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_6_sram_inv ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_1__0 ( .A ( chanx_right_in[2] ) , 
    .X ( ropt_net_192 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_2__1 ( .A ( chanx_right_in[4] ) , 
    .X ( ropt_net_185 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_3__2 ( .A ( chanx_right_in[5] ) , 
    .X ( ropt_net_189 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_150 ( .LO ( SYNOPSYS_UNCONNECTED_1 ) , 
    .HI ( optlc_net_162 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_152 ( .LO ( SYNOPSYS_UNCONNECTED_2 ) , 
    .HI ( optlc_net_163 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_6__5 ( .A ( chanx_right_in[9] ) , 
    .X ( chanx_left_out[10] ) ) ;
sky130_fd_sc_hd__conb_1 optlc_154 ( .LO ( SYNOPSYS_UNCONNECTED_3 ) , 
    .HI ( optlc_net_164 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_156 ( .LO ( SYNOPSYS_UNCONNECTED_4 ) , 
    .HI ( optlc_net_165 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_9__8 ( .A ( chanx_right_in[13] ) , 
    .X ( chanx_left_out[14] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_751 ( .A ( chanx_right_in[10] ) , 
    .X ( ropt_net_210 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_752 ( .A ( ropt_net_169 ) , 
    .X ( ropt_net_203 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_753 ( .A ( chanx_right_in[16] ) , 
    .X ( ropt_net_197 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_754 ( .A ( chanx_right_in[12] ) , 
    .X ( ropt_net_208 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_755 ( .A ( ropt_net_172 ) , 
    .X ( ropt_net_202 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_779 ( .A ( ropt_net_195 ) , 
    .X ( chany_bottom_out[5] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_16__15 ( .A ( chanx_left_in[5] ) , 
    .X ( aps_rename_2_ ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_756 ( .A ( ropt_net_173 ) , 
    .X ( ropt_net_196 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_757 ( .A ( chanx_left_in[9] ) , 
    .X ( ropt_net_212 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_758 ( .A ( ropt_net_175 ) , 
    .X ( ropt_net_211 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_759 ( .A ( ropt_net_176 ) , 
    .X ( ropt_net_195 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_760 ( .A ( chanx_right_in[14] ) , 
    .X ( chanx_left_out[15] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_761 ( .A ( chanx_left_in[14] ) , 
    .X ( ropt_net_213 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_762 ( .A ( chanx_left_in[12] ) , 
    .X ( ropt_net_209 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_763 ( .A ( chanx_left_in[17] ) , 
    .X ( chanx_right_out[18] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_780 ( .A ( ropt_net_196 ) , 
    .X ( chanx_left_out[18] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_764 ( .A ( chanx_right_in[18] ) , 
    .X ( chanx_left_out[19] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_RR_76 ( .A ( chanx_right_in[8] ) , 
    .X ( ropt_net_184 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_765 ( .A ( chanx_left_in[8] ) , 
    .X ( chanx_right_out[9] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_766 ( .A ( chanx_left_in[10] ) , 
    .X ( ropt_net_214 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_781 ( .A ( ropt_net_197 ) , 
    .X ( chanx_left_out[17] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_782 ( .A ( ropt_net_198 ) , 
    .X ( chanx_left_out[5] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_785 ( .A ( ropt_net_199 ) , 
    .X ( chanx_left_out[3] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_768 ( .A ( ropt_net_184 ) , 
    .X ( chanx_left_out[9] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_83 ( .A ( chanx_left_in[4] ) , 
    .X ( BUF_net_83 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_769 ( .A ( ropt_net_185 ) , 
    .X ( ropt_net_198 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_770 ( .A ( ropt_net_186 ) , 
    .X ( chanx_right_out[3] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_786 ( .A ( ropt_net_200 ) , 
    .X ( chanx_right_out[7] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_787 ( .A ( ropt_net_201 ) , 
    .X ( chanx_right_out[6] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_771 ( .A ( ropt_net_187 ) , 
    .X ( ropt_net_200 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_788 ( .A ( ropt_net_202 ) , 
    .X ( chanx_right_out[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_90 ( .A ( chanx_left_in[13] ) , 
    .X ( ropt_net_188 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_790 ( .A ( ropt_net_203 ) , 
    .X ( chany_bottom_out[13] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_92 ( .A ( chanx_left_in[16] ) , 
    .X ( BUF_net_92 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_RR_93 ( .A ( chanx_left_in[18] ) , 
    .X ( ropt_net_191 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_772 ( .A ( ropt_net_188 ) , 
    .X ( ropt_net_204 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_773 ( .A ( ropt_net_189 ) , 
    .X ( chanx_left_out[6] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_775 ( .A ( ropt_net_190 ) , 
    .X ( chanx_left_out[7] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_777 ( .A ( ropt_net_191 ) , 
    .X ( chanx_right_out[19] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_778 ( .A ( ropt_net_192 ) , 
    .X ( ropt_net_199 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_792 ( .A ( ropt_net_204 ) , 
    .X ( chanx_right_out[14] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 BUFT_RR_114 ( .A ( BUF_net_83 ) , 
    .X ( ropt_net_206 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 BUFT_RR_115 ( .A ( aps_rename_2_ ) , 
    .X ( ropt_net_201 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_116 ( .A ( chanx_left_in[6] ) , 
    .X ( ropt_net_187 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_793 ( .A ( ropt_net_205 ) , 
    .X ( chanx_right_out[17] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_794 ( .A ( ropt_net_206 ) , 
    .X ( chanx_right_out[5] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_796 ( .A ( ropt_net_207 ) , 
    .X ( chany_bottom_out[2] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_P_126 ( .A ( chanx_right_in[6] ) , 
    .X ( ropt_net_190 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_P_127 ( .A ( chanx_left_in[2] ) , 
    .X ( ropt_net_186 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_802 ( .A ( ropt_net_208 ) , 
    .X ( chanx_left_out[13] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_804 ( .A ( ropt_net_209 ) , 
    .X ( chanx_right_out[13] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_805 ( .A ( ropt_net_210 ) , 
    .X ( chanx_left_out[11] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_806 ( .A ( ropt_net_211 ) , 
    .X ( chany_bottom_out[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_P_144 ( .A ( chanx_right_in[17] ) , 
    .X ( ropt_net_173 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_807 ( .A ( ropt_net_212 ) , 
    .X ( chanx_right_out[10] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_808 ( .A ( ropt_net_213 ) , 
    .X ( chanx_right_out[15] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 BUFT_P_147 ( .A ( BUF_net_92 ) , 
    .X ( ropt_net_205 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_809 ( .A ( ropt_net_214 ) , 
    .X ( chanx_right_out[11] ) ) ;
endmodule


module mux_tree_tapbuf_size7_mem_1_2 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 FTB_28__79 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size7_mem_0_2 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_27__78 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size7_mem_2_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_26__77 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size7_mem_6 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_25__76 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_35 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size7_1_2 ( in , sram , sram_inv , out , p0 ) ;
input  [0:6] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;

const1_35 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_3_ ( .A0 ( p0 ) , .A1 ( in[6] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
endmodule


module const1_26_3 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size7_0_2 ( in , sram , sram_inv , out , p0 ) ;
input  [0:6] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;

const1_26_3 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_3_ ( .A0 ( p0 ) , .A1 ( in[6] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
endmodule


module const1_25_3 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size7_2_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:6] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;

const1_25_3 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_3_ ( .A0 ( p0 ) , .A1 ( in[6] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
endmodule


module const1_24_3 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size7_6 ( in , sram , sram_inv , out , p0 ) ;
input  [0:6] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;

const1_24_3 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_3_ ( .A0 ( p0 ) , .A1 ( in[6] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
endmodule


module mux_tree_tapbuf_size10_mem_4 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_24__75 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size10_mem_3 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_23__74 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size10_mem_5 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_22__73 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size10_mem_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_21__72 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size10_mem_0 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_20__71 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size10_mem_2 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_19__70 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size10_mem_7 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_18__69 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size10_mem_6 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_17__68 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size10_mem_8 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_16__67 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size10_mem_10 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_15__66 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size10_mem_9 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_14__65 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size10_mem_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_13__64 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_23_3 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size10_4 ( in , sram , sram_inv , out , p0 ) ;
input  [0:9] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

const1_23_3 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[6] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[8] ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[9] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
endmodule


module const1_22_3 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size10_3 ( in , sram , sram_inv , out , p0 ) ;
input  [0:9] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

const1_22_3 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[6] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[8] ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[9] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
endmodule


module const1_21_3 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size10_5 ( in , sram , sram_inv , out , p0 ) ;
input  [0:9] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

const1_21_3 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[6] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[8] ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[9] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
endmodule


module const1_20_3 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size10_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:9] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

const1_20_3 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[6] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[8] ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[9] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
endmodule


module const1_19_3 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size10_0 ( in , sram , sram_inv , out , p0 ) ;
input  [0:9] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

const1_19_3 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[6] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[8] ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[9] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
endmodule


module const1_18_3 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size10_2 ( in , sram , sram_inv , out , p0 ) ;
input  [0:9] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

const1_18_3 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[6] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[8] ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[9] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
endmodule


module const1_17_3 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size10_7 ( in , sram , sram_inv , out , p0 ) ;
input  [0:9] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

const1_17_3 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[6] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[8] ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[9] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
endmodule


module const1_16_4 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size10_6 ( in , sram , sram_inv , out , p0 ) ;
input  [0:9] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

const1_16_4 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[6] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[8] ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[9] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
endmodule


module const1_15_4 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size10_8 ( in , sram , sram_inv , out , p0 ) ;
input  [0:9] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

const1_15_4 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[6] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[8] ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[9] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
endmodule


module const1_14_4 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size10_10 ( in , sram , sram_inv , out , p0 ) ;
input  [0:9] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

const1_14_4 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[6] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[8] ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[9] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
endmodule


module const1_13_4 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size10_9 ( in , sram , sram_inv , out , p0 ) ;
input  [0:9] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

const1_13_4 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[6] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[8] ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[9] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
endmodule


module const1_12_4 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size10_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:9] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

const1_12_4 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[6] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[8] ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[9] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
endmodule


module mux_tree_tapbuf_size16_mem_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:4] mem_out ;
output [0:4] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_4_ ( .D ( mem_out[3] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[4] ) , .Q_N ( mem_outb[4] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_12__63 ( .A ( mem_out[4] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size16_mem_0 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:4] mem_out ;
output [0:4] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_4_ ( .D ( mem_out[3] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[4] ) , .Q_N ( mem_outb[4] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_11__62 ( .A ( mem_out[4] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size16_mem_2 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:4] mem_out ;
output [0:4] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_4_ ( .D ( mem_out[3] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[4] ) , .Q_N ( mem_outb[4] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_10__61 ( .A ( mem_out[4] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size16_mem ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:4] mem_out ;
output [0:4] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_4_ ( .D ( mem_out[3] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[4] ) , .Q_N ( mem_outb[4] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_9__60 ( .A ( mem_out[4] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_11_4 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size16_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:15] in ;
input  [0:4] sram ;
input  [0:4] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_10_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_11_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_12_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_13_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_14_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_15_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

const1_11_4 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_15_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( in[2] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[4] ) , .A1 ( in[3] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[6] ) , .A1 ( in[5] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( in[8] ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_4_ ( .A0 ( in[10] ) , .A1 ( in[9] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_5_ ( .A0 ( in[12] ) , .A1 ( in[11] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_6_ ( .A0 ( in[14] ) , .A1 ( in[13] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_7_ ( .A0 ( p0 ) , .A1 ( in[15] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_10_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_2_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_11_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_3_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_12_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_10_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_13_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_12_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_11_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_14_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l5_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_14_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_13_X[0] ) , .S ( sram[4] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_15_X[0] ) ) ;
endmodule


module const1_10_4 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size16_0 ( in , sram , sram_inv , out , p0 ) ;
input  [0:15] in ;
input  [0:4] sram ;
input  [0:4] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_10_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_11_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_12_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_13_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_14_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

const1_10_4 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( in[2] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[4] ) , .A1 ( in[3] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[6] ) , .A1 ( in[5] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( in[8] ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_4_ ( .A0 ( in[10] ) , .A1 ( in[9] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_5_ ( .A0 ( in[12] ) , .A1 ( in[11] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_6_ ( .A0 ( in[14] ) , .A1 ( in[13] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_7_ ( .A0 ( p0 ) , .A1 ( in[15] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_10_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_2_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_11_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_3_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_12_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_10_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_13_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_12_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_11_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_14_X[0] ) ) ;
sky130_fd_sc_hd__mux2_4 mux_l5_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_14_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_13_X[0] ) , .S ( sram[4] ) , .X ( out[0] ) ) ;
endmodule


module const1_9_4 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size16_2 ( in , sram , sram_inv , out , p0 ) ;
input  [0:15] in ;
input  [0:4] sram ;
input  [0:4] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_10_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_11_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_12_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_13_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_14_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_15_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

const1_9_4 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_15_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( in[2] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[4] ) , .A1 ( in[3] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[6] ) , .A1 ( in[5] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( in[8] ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_4_ ( .A0 ( in[10] ) , .A1 ( in[9] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_5_ ( .A0 ( in[12] ) , .A1 ( in[11] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_6_ ( .A0 ( in[14] ) , .A1 ( in[13] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_7_ ( .A0 ( p0 ) , .A1 ( in[15] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_10_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_2_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_11_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_3_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_12_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_10_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_13_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_12_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_11_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_14_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l5_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_14_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_13_X[0] ) , .S ( sram[4] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_15_X[0] ) ) ;
endmodule


module const1_8_4 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size16 ( in , sram , sram_inv , out , p0 ) ;
input  [0:15] in ;
input  [0:4] sram ;
input  [0:4] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_10_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_11_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_12_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_13_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_14_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_15_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

const1_8_4 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_15_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( in[2] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[4] ) , .A1 ( in[3] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[6] ) , .A1 ( in[5] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( in[8] ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_4_ ( .A0 ( in[10] ) , .A1 ( in[9] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_5_ ( .A0 ( in[12] ) , .A1 ( in[11] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_6_ ( .A0 ( in[14] ) , .A1 ( in[13] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_7_ ( .A0 ( p0 ) , .A1 ( in[15] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_10_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_2_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_11_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_3_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_12_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_10_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_13_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_12_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_11_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_14_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l5_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_14_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_13_X[0] ) , .S ( sram[4] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_15_X[0] ) ) ;
endmodule


module mux_tree_tapbuf_size12_mem_3 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_8__59 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size12_mem_2 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_7__58 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size12_mem_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_6__57 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size12_mem_0 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_5__56 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size12_mem_5 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_4__55 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size12_mem_4 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_3__54 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size12_mem ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_2__53 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size12_mem_6 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_1__52 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_7_4 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size12_3 ( in , sram , sram_inv , out , p0 ) ;
input  [0:11] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_10_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_11_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

const1_7_4 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_11_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_3_ ( .A0 ( in[7] ) , .A1 ( in[6] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_4_ ( .A0 ( in[9] ) , .A1 ( in[8] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[10] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[11] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_10_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_10_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_11_X[0] ) ) ;
endmodule


module const1_6_5 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size12_2 ( in , sram , sram_inv , out , p0 ) ;
input  [0:11] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_10_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_11_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

const1_6_5 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_11_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_3_ ( .A0 ( in[7] ) , .A1 ( in[6] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_4_ ( .A0 ( in[9] ) , .A1 ( in[8] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[10] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[11] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_10_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_10_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_11_X[0] ) ) ;
endmodule


module const1_5_5 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size12_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:11] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_10_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_11_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

const1_5_5 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_11_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_3_ ( .A0 ( in[7] ) , .A1 ( in[6] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_4_ ( .A0 ( in[9] ) , .A1 ( in[8] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[10] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[11] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_10_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_10_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_11_X[0] ) ) ;
endmodule


module const1_4_5 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size12_0 ( in , sram , sram_inv , out , p0 ) ;
input  [0:11] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_10_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_11_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

const1_4_5 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_11_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_3_ ( .A0 ( in[7] ) , .A1 ( in[6] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_4_ ( .A0 ( in[9] ) , .A1 ( in[8] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[10] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[11] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_10_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_10_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_11_X[0] ) ) ;
endmodule


module const1_3_5 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size12_5 ( in , sram , sram_inv , out , p0 ) ;
input  [0:11] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_10_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_11_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

const1_3_5 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_11_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_3_ ( .A0 ( in[7] ) , .A1 ( in[6] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_4_ ( .A0 ( in[9] ) , .A1 ( in[8] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[10] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[11] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_10_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_10_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_11_X[0] ) ) ;
endmodule


module const1_2_5 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size12_4 ( in , sram , sram_inv , out , p0 ) ;
input  [0:11] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_10_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_11_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

const1_2_5 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_11_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_3_ ( .A0 ( in[7] ) , .A1 ( in[6] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_4_ ( .A0 ( in[9] ) , .A1 ( in[8] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[10] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[11] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_10_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_10_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_11_X[0] ) ) ;
endmodule


module const1_1_5 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size12 ( in , sram , sram_inv , out , p0 ) ;
input  [0:11] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_10_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

const1_1_5 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_3_ ( .A0 ( in[7] ) , .A1 ( in[6] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_4_ ( .A0 ( in[9] ) , .A1 ( in[8] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[10] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[11] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_10_X[0] ) ) ;
sky130_fd_sc_hd__mux2_8 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_10_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , .S ( sram[3] ) , .X ( out[0] ) ) ;
endmodule


module const1_0_5 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size12_6 ( in , sram , sram_inv , out , p0 ) ;
input  [0:11] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_10_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_11_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

const1_0_5 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_11_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_3_ ( .A0 ( in[7] ) , .A1 ( in[6] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_4_ ( .A0 ( in[9] ) , .A1 ( in[8] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[10] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[11] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_10_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_10_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_11_X[0] ) ) ;
endmodule


module sb_1__1_ ( prog_clk , chany_top_in , top_left_grid_pin_34_ , 
    top_left_grid_pin_35_ , top_left_grid_pin_36_ , top_left_grid_pin_37_ , 
    top_left_grid_pin_38_ , top_left_grid_pin_39_ , top_left_grid_pin_40_ , 
    top_left_grid_pin_41_ , chanx_right_in , right_top_grid_pin_42_ , 
    right_top_grid_pin_43_ , right_top_grid_pin_44_ , right_top_grid_pin_45_ , 
    right_top_grid_pin_46_ , right_top_grid_pin_47_ , right_top_grid_pin_48_ , 
    right_top_grid_pin_49_ , chany_bottom_in , bottom_left_grid_pin_34_ , 
    bottom_left_grid_pin_35_ , bottom_left_grid_pin_36_ , 
    bottom_left_grid_pin_37_ , bottom_left_grid_pin_38_ , 
    bottom_left_grid_pin_39_ , bottom_left_grid_pin_40_ , 
    bottom_left_grid_pin_41_ , chanx_left_in , left_top_grid_pin_42_ , 
    left_top_grid_pin_43_ , left_top_grid_pin_44_ , left_top_grid_pin_45_ , 
    left_top_grid_pin_46_ , left_top_grid_pin_47_ , left_top_grid_pin_48_ , 
    left_top_grid_pin_49_ , ccff_head , chany_top_out , chanx_right_out , 
    chany_bottom_out , chanx_left_out , ccff_tail ) ;
input  [0:0] prog_clk ;
input  [0:19] chany_top_in ;
input  [0:0] top_left_grid_pin_34_ ;
input  [0:0] top_left_grid_pin_35_ ;
input  [0:0] top_left_grid_pin_36_ ;
input  [0:0] top_left_grid_pin_37_ ;
input  [0:0] top_left_grid_pin_38_ ;
input  [0:0] top_left_grid_pin_39_ ;
input  [0:0] top_left_grid_pin_40_ ;
input  [0:0] top_left_grid_pin_41_ ;
input  [0:19] chanx_right_in ;
input  [0:0] right_top_grid_pin_42_ ;
input  [0:0] right_top_grid_pin_43_ ;
input  [0:0] right_top_grid_pin_44_ ;
input  [0:0] right_top_grid_pin_45_ ;
input  [0:0] right_top_grid_pin_46_ ;
input  [0:0] right_top_grid_pin_47_ ;
input  [0:0] right_top_grid_pin_48_ ;
input  [0:0] right_top_grid_pin_49_ ;
input  [0:19] chany_bottom_in ;
input  [0:0] bottom_left_grid_pin_34_ ;
input  [0:0] bottom_left_grid_pin_35_ ;
input  [0:0] bottom_left_grid_pin_36_ ;
input  [0:0] bottom_left_grid_pin_37_ ;
input  [0:0] bottom_left_grid_pin_38_ ;
input  [0:0] bottom_left_grid_pin_39_ ;
input  [0:0] bottom_left_grid_pin_40_ ;
input  [0:0] bottom_left_grid_pin_41_ ;
input  [0:19] chanx_left_in ;
input  [0:0] left_top_grid_pin_42_ ;
input  [0:0] left_top_grid_pin_43_ ;
input  [0:0] left_top_grid_pin_44_ ;
input  [0:0] left_top_grid_pin_45_ ;
input  [0:0] left_top_grid_pin_46_ ;
input  [0:0] left_top_grid_pin_47_ ;
input  [0:0] left_top_grid_pin_48_ ;
input  [0:0] left_top_grid_pin_49_ ;
input  [0:0] ccff_head ;
output [0:19] chany_top_out ;
output [0:19] chanx_right_out ;
output [0:19] chany_bottom_out ;
output [0:19] chanx_left_out ;
output [0:0] ccff_tail ;

wire [0:3] mux_tree_tapbuf_size10_0_sram ;
wire [0:3] mux_tree_tapbuf_size10_0_sram_inv ;
wire [0:3] mux_tree_tapbuf_size10_10_sram ;
wire [0:3] mux_tree_tapbuf_size10_10_sram_inv ;
wire [0:3] mux_tree_tapbuf_size10_11_sram ;
wire [0:3] mux_tree_tapbuf_size10_11_sram_inv ;
wire [0:3] mux_tree_tapbuf_size10_1_sram ;
wire [0:3] mux_tree_tapbuf_size10_1_sram_inv ;
wire [0:3] mux_tree_tapbuf_size10_2_sram ;
wire [0:3] mux_tree_tapbuf_size10_2_sram_inv ;
wire [0:3] mux_tree_tapbuf_size10_3_sram ;
wire [0:3] mux_tree_tapbuf_size10_3_sram_inv ;
wire [0:3] mux_tree_tapbuf_size10_4_sram ;
wire [0:3] mux_tree_tapbuf_size10_4_sram_inv ;
wire [0:3] mux_tree_tapbuf_size10_5_sram ;
wire [0:3] mux_tree_tapbuf_size10_5_sram_inv ;
wire [0:3] mux_tree_tapbuf_size10_6_sram ;
wire [0:3] mux_tree_tapbuf_size10_6_sram_inv ;
wire [0:3] mux_tree_tapbuf_size10_7_sram ;
wire [0:3] mux_tree_tapbuf_size10_7_sram_inv ;
wire [0:3] mux_tree_tapbuf_size10_8_sram ;
wire [0:3] mux_tree_tapbuf_size10_8_sram_inv ;
wire [0:3] mux_tree_tapbuf_size10_9_sram ;
wire [0:3] mux_tree_tapbuf_size10_9_sram_inv ;
wire [0:0] mux_tree_tapbuf_size10_mem_0_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size10_mem_10_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size10_mem_11_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size10_mem_1_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size10_mem_2_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size10_mem_3_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size10_mem_4_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size10_mem_5_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size10_mem_6_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size10_mem_7_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size10_mem_8_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size10_mem_9_ccff_tail ;
wire [0:3] mux_tree_tapbuf_size12_0_sram ;
wire [0:3] mux_tree_tapbuf_size12_0_sram_inv ;
wire [0:3] mux_tree_tapbuf_size12_1_sram ;
wire [0:3] mux_tree_tapbuf_size12_1_sram_inv ;
wire [0:3] mux_tree_tapbuf_size12_2_sram ;
wire [0:3] mux_tree_tapbuf_size12_2_sram_inv ;
wire [0:3] mux_tree_tapbuf_size12_3_sram ;
wire [0:3] mux_tree_tapbuf_size12_3_sram_inv ;
wire [0:3] mux_tree_tapbuf_size12_4_sram ;
wire [0:3] mux_tree_tapbuf_size12_4_sram_inv ;
wire [0:3] mux_tree_tapbuf_size12_5_sram ;
wire [0:3] mux_tree_tapbuf_size12_5_sram_inv ;
wire [0:3] mux_tree_tapbuf_size12_6_sram ;
wire [0:3] mux_tree_tapbuf_size12_6_sram_inv ;
wire [0:3] mux_tree_tapbuf_size12_7_sram ;
wire [0:3] mux_tree_tapbuf_size12_7_sram_inv ;
wire [0:0] mux_tree_tapbuf_size12_mem_0_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size12_mem_1_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size12_mem_2_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size12_mem_3_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size12_mem_4_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size12_mem_5_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size12_mem_6_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size12_mem_7_ccff_tail ;
wire [0:4] mux_tree_tapbuf_size16_0_sram ;
wire [0:4] mux_tree_tapbuf_size16_0_sram_inv ;
wire [0:4] mux_tree_tapbuf_size16_1_sram ;
wire [0:4] mux_tree_tapbuf_size16_1_sram_inv ;
wire [0:4] mux_tree_tapbuf_size16_2_sram ;
wire [0:4] mux_tree_tapbuf_size16_2_sram_inv ;
wire [0:4] mux_tree_tapbuf_size16_3_sram ;
wire [0:4] mux_tree_tapbuf_size16_3_sram_inv ;
wire [0:0] mux_tree_tapbuf_size16_mem_0_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size16_mem_1_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size16_mem_2_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size16_mem_3_ccff_tail ;
wire [0:2] mux_tree_tapbuf_size7_0_sram ;
wire [0:2] mux_tree_tapbuf_size7_0_sram_inv ;
wire [0:2] mux_tree_tapbuf_size7_1_sram ;
wire [0:2] mux_tree_tapbuf_size7_1_sram_inv ;
wire [0:2] mux_tree_tapbuf_size7_2_sram ;
wire [0:2] mux_tree_tapbuf_size7_2_sram_inv ;
wire [0:2] mux_tree_tapbuf_size7_3_sram ;
wire [0:2] mux_tree_tapbuf_size7_3_sram_inv ;
wire [0:0] mux_tree_tapbuf_size7_mem_0_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size7_mem_1_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size7_mem_2_ccff_tail ;

mux_tree_tapbuf_size12_6 mux_top_track_0 (
    .in ( { top_left_grid_pin_34_[0] , top_left_grid_pin_36_[0] , 
        top_left_grid_pin_38_[0] , top_left_grid_pin_40_[0] , 
        chanx_right_in[1] , chanx_right_in[2] , chanx_right_in[12] , 
        chany_bottom_in[2] , chany_bottom_in[12] , chanx_left_in[0] , 
        chanx_left_in[2] , chanx_left_in[12] } ) ,
    .sram ( mux_tree_tapbuf_size12_0_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size12_0_sram_inv ) , 
    .out ( chany_top_out[0] ) , .p0 ( optlc_net_147 ) ) ;
mux_tree_tapbuf_size12 mux_top_track_2 (
    .in ( { top_left_grid_pin_35_[0] , top_left_grid_pin_37_[0] , 
        top_left_grid_pin_39_[0] , top_left_grid_pin_41_[0] , 
        chanx_right_in[3] , chanx_right_in[4] , chanx_right_in[13] , 
        chany_bottom_in[4] , chany_bottom_in[13] , chanx_left_in[4] , 
        chanx_left_in[13] , chanx_left_in[19] } ) ,
    .sram ( mux_tree_tapbuf_size12_1_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size12_1_sram_inv ) , 
    .out ( chany_top_out[1] ) , .p0 ( optlc_net_145 ) ) ;
mux_tree_tapbuf_size12_4 mux_right_track_0 (
    .in ( { chany_top_in[2] , chany_top_in[12] , chany_top_in[19] , 
        right_top_grid_pin_42_[0] , right_top_grid_pin_44_[0] , 
        right_top_grid_pin_46_[0] , right_top_grid_pin_48_[0] , 
        chany_bottom_in[2] , chany_bottom_in[12] , chany_bottom_in[15] , 
        chanx_left_in[2] , chanx_left_in[12] } ) ,
    .sram ( mux_tree_tapbuf_size12_2_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size12_2_sram_inv ) , 
    .out ( chanx_right_out[0] ) , .p0 ( optlc_net_145 ) ) ;
mux_tree_tapbuf_size12_5 mux_right_track_2 (
    .in ( { chany_top_in[0] , chany_top_in[4] , chany_top_in[13] , 
        right_top_grid_pin_43_[0] , right_top_grid_pin_45_[0] , 
        right_top_grid_pin_47_[0] , right_top_grid_pin_49_[0] , 
        chany_bottom_in[4] , chany_bottom_in[11] , chany_bottom_in[13] , 
        chanx_left_in[4] , chanx_left_in[13] } ) ,
    .sram ( mux_tree_tapbuf_size12_3_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size12_3_sram_inv ) , 
    .out ( chanx_right_out[1] ) , .p0 ( optlc_net_145 ) ) ;
mux_tree_tapbuf_size12_0 mux_bottom_track_1 (
    .in ( { chany_top_in[2] , chany_top_in[12] , chanx_right_in[2] , 
        chanx_right_in[12] , chanx_right_in[15] , 
        bottom_left_grid_pin_34_[0] , bottom_left_grid_pin_36_[0] , 
        bottom_left_grid_pin_38_[0] , bottom_left_grid_pin_40_[0] , 
        chanx_left_in[1] , chanx_left_in[2] , chanx_left_in[12] } ) ,
    .sram ( mux_tree_tapbuf_size12_4_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size12_4_sram_inv ) , 
    .out ( chany_bottom_out[0] ) , .p0 ( optlc_net_144 ) ) ;
mux_tree_tapbuf_size12_1 mux_bottom_track_3 (
    .in ( { chany_top_in[4] , chany_top_in[13] , chanx_right_in[4] , 
        chanx_right_in[11] , chanx_right_in[13] , 
        bottom_left_grid_pin_35_[0] , bottom_left_grid_pin_37_[0] , 
        bottom_left_grid_pin_39_[0] , bottom_left_grid_pin_41_[0] , 
        chanx_left_in[3] , chanx_left_in[4] , chanx_left_in[13] } ) ,
    .sram ( mux_tree_tapbuf_size12_5_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size12_5_sram_inv ) , 
    .out ( chany_bottom_out[1] ) , .p0 ( optlc_net_146 ) ) ;
mux_tree_tapbuf_size12_2 mux_left_track_1 (
    .in ( { chany_top_in[0] , chany_top_in[2] , chany_top_in[12] , 
        chanx_right_in[2] , chanx_right_in[12] , chany_bottom_in[2] , 
        chany_bottom_in[12] , chany_bottom_in[19] , left_top_grid_pin_42_[0] , 
        left_top_grid_pin_44_[0] , left_top_grid_pin_46_[0] , 
        left_top_grid_pin_48_[0] } ) ,
    .sram ( mux_tree_tapbuf_size12_6_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size12_6_sram_inv ) , 
    .out ( chanx_left_out[0] ) , .p0 ( optlc_net_147 ) ) ;
mux_tree_tapbuf_size12_3 mux_left_track_3 (
    .in ( { chany_top_in[4] , chany_top_in[13] , chany_top_in[19] , 
        chanx_right_in[4] , chanx_right_in[13] , chany_bottom_in[0] , 
        chany_bottom_in[4] , chany_bottom_in[13] , left_top_grid_pin_43_[0] , 
        left_top_grid_pin_45_[0] , left_top_grid_pin_47_[0] , 
        left_top_grid_pin_49_[0] } ) ,
    .sram ( mux_tree_tapbuf_size12_7_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size12_7_sram_inv ) , 
    .out ( chanx_left_out[1] ) , .p0 ( optlc_net_147 ) ) ;
mux_tree_tapbuf_size12_mem_6 mem_top_track_0 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( ccff_head ) , 
    .ccff_tail ( mux_tree_tapbuf_size12_mem_0_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size12_0_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size12_0_sram_inv ) ) ;
mux_tree_tapbuf_size12_mem mem_top_track_2 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size12_mem_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size12_mem_1_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size12_1_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size12_1_sram_inv ) ) ;
mux_tree_tapbuf_size12_mem_4 mem_right_track_0 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size7_mem_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size12_mem_2_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size12_2_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size12_2_sram_inv ) ) ;
mux_tree_tapbuf_size12_mem_5 mem_right_track_2 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size12_mem_2_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size12_mem_3_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size12_3_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size12_3_sram_inv ) ) ;
mux_tree_tapbuf_size12_mem_0 mem_bottom_track_1 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size7_mem_1_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size12_mem_4_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size12_4_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size12_4_sram_inv ) ) ;
mux_tree_tapbuf_size12_mem_1 mem_bottom_track_3 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size12_mem_4_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size12_mem_5_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size12_5_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size12_5_sram_inv ) ) ;
mux_tree_tapbuf_size12_mem_2 mem_left_track_1 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size7_mem_2_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size12_mem_6_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size12_6_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size12_6_sram_inv ) ) ;
mux_tree_tapbuf_size12_mem_3 mem_left_track_3 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size12_mem_6_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size12_mem_7_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size12_7_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size12_7_sram_inv ) ) ;
mux_tree_tapbuf_size16 mux_top_track_4 (
    .in ( { top_left_grid_pin_34_[0] , top_left_grid_pin_35_[0] , 
        top_left_grid_pin_36_[0] , top_left_grid_pin_37_[0] , 
        top_left_grid_pin_38_[0] , top_left_grid_pin_39_[0] , 
        top_left_grid_pin_40_[0] , top_left_grid_pin_41_[0] , 
        chanx_right_in[5] , chanx_right_in[7] , chanx_right_in[14] , 
        chany_bottom_in[5] , chany_bottom_in[14] , chanx_left_in[5] , 
        chanx_left_in[14] , chanx_left_in[15] } ) ,
    .sram ( mux_tree_tapbuf_size16_0_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size16_0_sram_inv ) , 
    .out ( chany_top_out[2] ) , .p0 ( optlc_net_147 ) ) ;
mux_tree_tapbuf_size16_2 mux_right_track_4 (
    .in ( { chany_top_in[1] , chany_top_in[5] , chany_top_in[14] , 
        right_top_grid_pin_42_[0] , right_top_grid_pin_43_[0] , 
        right_top_grid_pin_44_[0] , right_top_grid_pin_45_[0] , 
        right_top_grid_pin_46_[0] , right_top_grid_pin_47_[0] , 
        right_top_grid_pin_48_[0] , right_top_grid_pin_49_[0] , 
        chany_bottom_in[5] , chany_bottom_in[7] , chany_bottom_in[14] , 
        chanx_left_in[5] , chanx_left_in[14] } ) ,
    .sram ( mux_tree_tapbuf_size16_1_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size16_1_sram_inv ) , 
    .out ( chanx_right_out[2] ) , .p0 ( optlc_net_145 ) ) ;
mux_tree_tapbuf_size16_0 mux_bottom_track_5 (
    .in ( { chany_top_in[5] , chany_top_in[14] , chanx_right_in[5] , 
        chanx_right_in[7] , chanx_right_in[14] , bottom_left_grid_pin_34_[0] , 
        bottom_left_grid_pin_35_[0] , bottom_left_grid_pin_36_[0] , 
        bottom_left_grid_pin_37_[0] , bottom_left_grid_pin_38_[0] , 
        bottom_left_grid_pin_39_[0] , bottom_left_grid_pin_40_[0] , 
        bottom_left_grid_pin_41_[0] , chanx_left_in[5] , chanx_left_in[7] , 
        chanx_left_in[14] } ) ,
    .sram ( mux_tree_tapbuf_size16_2_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size16_2_sram_inv ) , 
    .out ( chany_bottom_out[2] ) , .p0 ( optlc_net_144 ) ) ;
mux_tree_tapbuf_size16_1 mux_left_track_5 (
    .in ( { chany_top_in[5] , chany_top_in[14] , chany_top_in[15] , 
        chanx_right_in[5] , chanx_right_in[14] , chany_bottom_in[1] , 
        chany_bottom_in[5] , chany_bottom_in[14] , left_top_grid_pin_42_[0] , 
        left_top_grid_pin_43_[0] , left_top_grid_pin_44_[0] , 
        left_top_grid_pin_45_[0] , left_top_grid_pin_46_[0] , 
        left_top_grid_pin_47_[0] , left_top_grid_pin_48_[0] , 
        left_top_grid_pin_49_[0] } ) ,
    .sram ( mux_tree_tapbuf_size16_3_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size16_3_sram_inv ) , 
    .out ( chanx_left_out[2] ) , .p0 ( optlc_net_147 ) ) ;
mux_tree_tapbuf_size16_mem mem_top_track_4 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size12_mem_1_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size16_mem_0_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size16_0_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size16_0_sram_inv ) ) ;
mux_tree_tapbuf_size16_mem_2 mem_right_track_4 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size12_mem_3_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size16_mem_1_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size16_1_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size16_1_sram_inv ) ) ;
mux_tree_tapbuf_size16_mem_0 mem_bottom_track_5 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size12_mem_5_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size16_mem_2_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size16_2_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size16_2_sram_inv ) ) ;
mux_tree_tapbuf_size16_mem_1 mem_left_track_5 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size12_mem_7_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size16_mem_3_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size16_3_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size16_3_sram_inv ) ) ;
mux_tree_tapbuf_size10_1 mux_top_track_8 (
    .in ( { top_left_grid_pin_34_[0] , top_left_grid_pin_38_[0] , 
        chanx_right_in[6] , chanx_right_in[11] , chanx_right_in[16] , 
        chany_bottom_in[6] , chany_bottom_in[16] , chanx_left_in[6] , 
        chanx_left_in[11] , chanx_left_in[16] } ) ,
    .sram ( mux_tree_tapbuf_size10_0_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size10_0_sram_inv ) , 
    .out ( chany_top_out[4] ) , .p0 ( optlc_net_144 ) ) ;
mux_tree_tapbuf_size10_9 mux_top_track_16 (
    .in ( { top_left_grid_pin_35_[0] , top_left_grid_pin_39_[0] , 
        chanx_right_in[8] , chanx_right_in[15] , chanx_right_in[17] , 
        chany_bottom_in[8] , chany_bottom_in[17] , chanx_left_in[7] , 
        chanx_left_in[8] , chanx_left_in[17] } ) ,
    .sram ( mux_tree_tapbuf_size10_1_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size10_1_sram_inv ) , 
    .out ( chany_top_out[8] ) , .p0 ( optlc_net_144 ) ) ;
mux_tree_tapbuf_size10_10 mux_top_track_24 (
    .in ( { top_left_grid_pin_36_[0] , top_left_grid_pin_40_[0] , 
        chanx_right_in[9] , chanx_right_in[18] , chanx_right_in[19] , 
        chany_bottom_in[9] , chany_bottom_in[18] , chanx_left_in[3] , 
        chanx_left_in[9] , chanx_left_in[18] } ) ,
    .sram ( mux_tree_tapbuf_size10_2_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size10_2_sram_inv ) , 
    .out ( chany_top_out[12] ) , .p0 ( optlc_net_145 ) ) ;
mux_tree_tapbuf_size10_8 mux_right_track_8 (
    .in ( { chany_top_in[3] , chany_top_in[6] , chany_top_in[16] , 
        right_top_grid_pin_42_[0] , right_top_grid_pin_46_[0] , 
        chany_bottom_in[3] , chany_bottom_in[6] , chany_bottom_in[16] , 
        chanx_left_in[6] , chanx_left_in[16] } ) ,
    .sram ( mux_tree_tapbuf_size10_3_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size10_3_sram_inv ) , 
    .out ( chanx_right_out[4] ) , .p0 ( optlc_net_144 ) ) ;
mux_tree_tapbuf_size10_6 mux_right_track_16 (
    .in ( { chany_top_in[7] , chany_top_in[8] , chany_top_in[17] , 
        right_top_grid_pin_43_[0] , right_top_grid_pin_47_[0] , 
        chany_bottom_in[1] , chany_bottom_in[8] , chany_bottom_in[17] , 
        chanx_left_in[8] , chanx_left_in[17] } ) ,
    .sram ( mux_tree_tapbuf_size10_4_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size10_4_sram_inv ) , 
    .out ( chanx_right_out[8] ) , .p0 ( optlc_net_144 ) ) ;
mux_tree_tapbuf_size10_7 mux_right_track_24 (
    .in ( { chany_top_in[9] , chany_top_in[11] , chany_top_in[18] , 
        right_top_grid_pin_44_[0] , right_top_grid_pin_48_[0] , 
        chany_bottom_in[0] , chany_bottom_in[9] , chany_bottom_in[18] , 
        chanx_left_in[9] , chanx_left_in[18] } ) ,
    .sram ( mux_tree_tapbuf_size10_5_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size10_5_sram_inv ) , 
    .out ( chanx_right_out[12] ) , .p0 ( optlc_net_145 ) ) ;
mux_tree_tapbuf_size10_2 mux_bottom_track_9 (
    .in ( { chany_top_in[6] , chany_top_in[16] , chanx_right_in[3] , 
        chanx_right_in[6] , chanx_right_in[16] , bottom_left_grid_pin_34_[0] , 
        bottom_left_grid_pin_38_[0] , chanx_left_in[6] , chanx_left_in[11] , 
        chanx_left_in[16] } ) ,
    .sram ( mux_tree_tapbuf_size10_6_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size10_6_sram_inv ) , 
    .out ( chany_bottom_out[4] ) , .p0 ( optlc_net_144 ) ) ;
mux_tree_tapbuf_size10_0 mux_bottom_track_17 (
    .in ( { chany_top_in[8] , chany_top_in[17] , chanx_right_in[1] , 
        chanx_right_in[8] , chanx_right_in[17] , bottom_left_grid_pin_35_[0] , 
        bottom_left_grid_pin_39_[0] , chanx_left_in[8] , chanx_left_in[15] , 
        chanx_left_in[17] } ) ,
    .sram ( mux_tree_tapbuf_size10_7_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size10_7_sram_inv ) , 
    .out ( chany_bottom_out[8] ) , .p0 ( optlc_net_146 ) ) ;
mux_tree_tapbuf_size10_1 mux_bottom_track_25 (
    .in ( { chany_top_in[9] , chany_top_in[18] , chanx_right_in[0] , 
        chanx_right_in[9] , chanx_right_in[18] , bottom_left_grid_pin_36_[0] , 
        bottom_left_grid_pin_40_[0] , chanx_left_in[9] , chanx_left_in[18] , 
        chanx_left_in[19] } ) ,
    .sram ( mux_tree_tapbuf_size10_8_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size10_8_sram_inv ) , 
    .out ( chany_bottom_out[12] ) , .p0 ( optlc_net_145 ) ) ;
mux_tree_tapbuf_size10_5 mux_left_track_9 (
    .in ( { chany_top_in[6] , chany_top_in[11] , chany_top_in[16] , 
        chanx_right_in[6] , chanx_right_in[16] , chany_bottom_in[3] , 
        chany_bottom_in[6] , chany_bottom_in[16] , left_top_grid_pin_42_[0] , 
        left_top_grid_pin_46_[0] } ) ,
    .sram ( mux_tree_tapbuf_size10_9_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size10_9_sram_inv ) , 
    .out ( chanx_left_out[4] ) , .p0 ( optlc_net_147 ) ) ;
mux_tree_tapbuf_size10_3 mux_left_track_17 (
    .in ( { chany_top_in[7] , chany_top_in[8] , chany_top_in[17] , 
        chanx_right_in[8] , chanx_right_in[17] , chany_bottom_in[7] , 
        chany_bottom_in[8] , chany_bottom_in[17] , left_top_grid_pin_43_[0] , 
        left_top_grid_pin_47_[0] } ) ,
    .sram ( mux_tree_tapbuf_size10_10_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size10_10_sram_inv ) , 
    .out ( chanx_left_out[8] ) , .p0 ( optlc_net_146 ) ) ;
mux_tree_tapbuf_size10_4 mux_left_track_25 (
    .in ( { chany_top_in[3] , chany_top_in[9] , chany_top_in[18] , 
        chanx_right_in[9] , chanx_right_in[18] , chany_bottom_in[9] , 
        chany_bottom_in[11] , chany_bottom_in[18] , left_top_grid_pin_44_[0] , 
        left_top_grid_pin_48_[0] } ) ,
    .sram ( mux_tree_tapbuf_size10_11_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size10_11_sram_inv ) , 
    .out ( chanx_left_out[12] ) , .p0 ( optlc_net_147 ) ) ;
mux_tree_tapbuf_size10_mem_1 mem_top_track_8 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size16_mem_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size10_mem_0_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size10_0_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size10_0_sram_inv ) ) ;
mux_tree_tapbuf_size10_mem_9 mem_top_track_16 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size10_mem_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size10_mem_1_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size10_1_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size10_1_sram_inv ) ) ;
mux_tree_tapbuf_size10_mem_10 mem_top_track_24 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size10_mem_1_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size10_mem_2_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size10_2_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size10_2_sram_inv ) ) ;
mux_tree_tapbuf_size10_mem_8 mem_right_track_8 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size16_mem_1_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size10_mem_3_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size10_3_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size10_3_sram_inv ) ) ;
mux_tree_tapbuf_size10_mem_6 mem_right_track_16 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size10_mem_3_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size10_mem_4_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size10_4_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size10_4_sram_inv ) ) ;
mux_tree_tapbuf_size10_mem_7 mem_right_track_24 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size10_mem_4_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size10_mem_5_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size10_5_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size10_5_sram_inv ) ) ;
mux_tree_tapbuf_size10_mem_2 mem_bottom_track_9 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size16_mem_2_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size10_mem_6_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size10_6_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size10_6_sram_inv ) ) ;
mux_tree_tapbuf_size10_mem_0 mem_bottom_track_17 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size10_mem_6_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size10_mem_7_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size10_7_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size10_7_sram_inv ) ) ;
mux_tree_tapbuf_size10_mem_1 mem_bottom_track_25 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size10_mem_7_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size10_mem_8_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size10_8_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size10_8_sram_inv ) ) ;
mux_tree_tapbuf_size10_mem_5 mem_left_track_9 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size16_mem_3_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size10_mem_9_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size10_9_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size10_9_sram_inv ) ) ;
mux_tree_tapbuf_size10_mem_3 mem_left_track_17 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size10_mem_9_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size10_mem_10_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size10_10_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size10_10_sram_inv ) ) ;
mux_tree_tapbuf_size10_mem_4 mem_left_track_25 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size10_mem_10_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size10_mem_11_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size10_11_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size10_11_sram_inv ) ) ;
mux_tree_tapbuf_size7_6 mux_top_track_32 (
    .in ( { top_left_grid_pin_37_[0] , top_left_grid_pin_41_[0] , 
        chanx_right_in[0] , chanx_right_in[10] , chany_bottom_in[10] , 
        chanx_left_in[1] , chanx_left_in[10] } ) ,
    .sram ( mux_tree_tapbuf_size7_0_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size7_0_sram_inv ) , 
    .out ( chany_top_out[16] ) , .p0 ( optlc_net_145 ) ) ;
mux_tree_tapbuf_size7_2_1 mux_right_track_32 (
    .in ( { chany_top_in[10] , chany_top_in[15] , right_top_grid_pin_45_[0] , 
        right_top_grid_pin_49_[0] , chany_bottom_in[10] , 
        chany_bottom_in[19] , chanx_left_in[10] } ) ,
    .sram ( mux_tree_tapbuf_size7_1_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size7_1_sram_inv ) , 
    .out ( chanx_right_out[16] ) , .p0 ( optlc_net_145 ) ) ;
mux_tree_tapbuf_size7_0_2 mux_bottom_track_33 (
    .in ( { chany_top_in[10] , chanx_right_in[10] , chanx_right_in[19] , 
        bottom_left_grid_pin_37_[0] , bottom_left_grid_pin_41_[0] , 
        chanx_left_in[0] , chanx_left_in[10] } ) ,
    .sram ( mux_tree_tapbuf_size7_2_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size7_2_sram_inv ) , 
    .out ( chany_bottom_out[16] ) , .p0 ( optlc_net_146 ) ) ;
mux_tree_tapbuf_size7_1_2 mux_left_track_33 (
    .in ( { chany_top_in[1] , chany_top_in[10] , chanx_right_in[10] , 
        chany_bottom_in[10] , chany_bottom_in[15] , left_top_grid_pin_45_[0] , 
        left_top_grid_pin_49_[0] } ) ,
    .sram ( mux_tree_tapbuf_size7_3_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size7_3_sram_inv ) , 
    .out ( chanx_left_out[16] ) , .p0 ( optlc_net_146 ) ) ;
mux_tree_tapbuf_size7_mem_6 mem_top_track_32 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size10_mem_2_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size7_mem_0_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size7_0_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size7_0_sram_inv ) ) ;
mux_tree_tapbuf_size7_mem_2_1 mem_right_track_32 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size10_mem_5_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size7_mem_1_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size7_1_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size7_1_sram_inv ) ) ;
mux_tree_tapbuf_size7_mem_0_2 mem_bottom_track_33 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size10_mem_8_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size7_mem_2_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size7_2_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size7_2_sram_inv ) ) ;
mux_tree_tapbuf_size7_mem_1_2 mem_left_track_33 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size10_mem_11_ccff_tail ) , 
    .ccff_tail ( ccff_tail ) , .mem_out ( mux_tree_tapbuf_size7_3_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size7_3_sram_inv ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_1__0 ( .A ( chany_top_in[2] ) , 
    .X ( chany_bottom_out[3] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_2__1 ( .A ( chany_top_in[4] ) , 
    .X ( chany_bottom_out[5] ) ) ;
sky130_fd_sc_hd__dlygate4sd1_1 FTB_3__2 ( .A ( chany_top_in[5] ) , 
    .X ( chany_bottom_out[6] ) ) ;
sky130_fd_sc_hd__conb_1 optlc_133 ( .LO ( SYNOPSYS_UNCONNECTED_1 ) , 
    .HI ( optlc_net_144 ) ) ;
sky130_fd_sc_hd__dlygate4sd1_1 FTB_5__4 ( .A ( chany_top_in[8] ) , 
    .X ( ropt_net_148 ) ) ;
sky130_fd_sc_hd__dlygate4sd1_1 FTB_6__5 ( .A ( chany_top_in[9] ) , 
    .X ( chany_bottom_out[10] ) ) ;
sky130_fd_sc_hd__dlygate4sd1_1 FTB_7__6 ( .A ( chany_top_in[10] ) , 
    .X ( chany_bottom_out[11] ) ) ;
sky130_fd_sc_hd__conb_1 optlc_135 ( .LO ( SYNOPSYS_UNCONNECTED_2 ) , 
    .HI ( optlc_net_145 ) ) ;
sky130_fd_sc_hd__dlygate4sd1_1 FTB_9__8 ( .A ( chany_top_in[13] ) , 
    .X ( chany_bottom_out[14] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_10__9 ( .A ( chany_top_in[14] ) , 
    .X ( chany_bottom_out[15] ) ) ;
sky130_fd_sc_hd__dlygate4sd1_1 FTB_11__10 ( .A ( chany_top_in[16] ) , 
    .X ( chany_bottom_out[17] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_12__11 ( .A ( chany_top_in[17] ) , 
    .X ( chany_bottom_out[18] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_746 ( .A ( ropt_net_148 ) , 
    .X ( chany_bottom_out[9] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_14__13 ( .A ( chanx_right_in[2] ) , 
    .X ( chanx_left_out[3] ) ) ;
sky130_fd_sc_hd__conb_1 optlc_137 ( .LO ( SYNOPSYS_UNCONNECTED_3 ) , 
    .HI ( optlc_net_146 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_16__15 ( .A ( chanx_right_in[5] ) , 
    .X ( chanx_left_out[6] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_17__16 ( .A ( chanx_right_in[6] ) , 
    .X ( aps_rename_2_ ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_18__17 ( .A ( chanx_right_in[8] ) , 
    .X ( aps_rename_3_ ) ) ;
sky130_fd_sc_hd__dlygate4sd1_1 FTB_19__18 ( .A ( chanx_right_in[9] ) , 
    .X ( chanx_left_out[10] ) ) ;
sky130_fd_sc_hd__dlygate4sd1_1 FTB_20__19 ( .A ( chanx_right_in[10] ) , 
    .X ( chanx_left_out[11] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_21__20 ( .A ( chanx_right_in[12] ) , 
    .X ( chanx_left_out[13] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_22__21 ( .A ( chanx_right_in[13] ) , 
    .X ( chanx_left_out[14] ) ) ;
sky130_fd_sc_hd__dlygate4sd1_1 FTB_23__22 ( .A ( chanx_right_in[14] ) , 
    .X ( chanx_left_out[15] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_748 ( .A ( ropt_net_149 ) , 
    .X ( chanx_left_out[19] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_753 ( .A ( chanx_left_in[16] ) , 
    .X ( chanx_right_out[17] ) ) ;
sky130_fd_sc_hd__dlygate4sd1_1 FTB_26__25 ( .A ( chanx_right_in[18] ) , 
    .X ( ropt_net_149 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_139 ( .LO ( SYNOPSYS_UNCONNECTED_4 ) , 
    .HI ( optlc_net_147 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_28__27 ( .A ( chany_bottom_in[4] ) , 
    .X ( chany_top_out[5] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_754 ( .A ( chanx_left_in[8] ) , 
    .X ( ropt_net_159 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_30__29 ( .A ( chany_bottom_in[6] ) , 
    .X ( chany_top_out[7] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_31__30 ( .A ( chany_bottom_in[8] ) , 
    .X ( chany_top_out[9] ) ) ;
sky130_fd_sc_hd__dlygate4sd1_1 FTB_32__31 ( .A ( chany_bottom_in[9] ) , 
    .X ( chany_top_out[10] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_33__32 ( .A ( chany_bottom_in[10] ) , 
    .X ( chany_top_out[11] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_761 ( .A ( ropt_net_152 ) , 
    .X ( ropt_net_157 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_35__34 ( .A ( chany_bottom_in[13] ) , 
    .X ( chany_top_out[14] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_762 ( .A ( ropt_net_153 ) , 
    .X ( ropt_net_155 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_763 ( .A ( ropt_net_154 ) , 
    .X ( chanx_right_out[15] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_767 ( .A ( ropt_net_155 ) , 
    .X ( chanx_right_out[18] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_39__38 ( .A ( chany_bottom_in[18] ) , 
    .X ( chany_top_out[19] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_768 ( .A ( ropt_net_156 ) , 
    .X ( chanx_right_out[7] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_769 ( .A ( ropt_net_157 ) , 
    .X ( chanx_right_out[11] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_42__41 ( .A ( chanx_left_in[5] ) , 
    .X ( chanx_right_out[6] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_774 ( .A ( ropt_net_158 ) , 
    .X ( chanx_right_out[5] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_775 ( .A ( ropt_net_159 ) , 
    .X ( chanx_right_out[9] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_45__44 ( .A ( chanx_left_in[9] ) , 
    .X ( chanx_right_out[10] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_46__45 ( .A ( chanx_left_in[10] ) , 
    .X ( ropt_net_152 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_48__47 ( .A ( chanx_left_in[13] ) , 
    .X ( chanx_right_out[14] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_49__48 ( .A ( chanx_left_in[14] ) , 
    .X ( ropt_net_154 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_RR_87 ( .A ( chanx_right_in[16] ) , 
    .X ( chanx_left_out[17] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_RR_89 ( .A ( chany_bottom_in[17] ) , 
    .X ( chany_top_out[18] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_90 ( .A ( chanx_left_in[6] ) , 
    .X ( BUF_net_90 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_RR_92 ( .A ( chanx_left_in[12] ) , 
    .X ( chanx_right_out[13] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_RR_95 ( .A ( chanx_left_in[18] ) , 
    .X ( chanx_right_out[19] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_RR_100 ( .A ( chany_top_in[6] ) , 
    .X ( chany_bottom_out[7] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_RR_101 ( .A ( chanx_left_in[2] ) , 
    .X ( chanx_right_out[3] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_RR_105 ( .A ( chany_top_in[18] ) , 
    .X ( chany_bottom_out[19] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 BUFT_RR_106 ( .A ( BUF_net_90 ) , 
    .X ( ropt_net_156 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_109 ( .A ( chanx_left_in[17] ) , 
    .X ( ropt_net_153 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_P_115 ( .A ( chany_top_in[12] ) , 
    .X ( chany_bottom_out[13] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_P_116 ( .A ( chanx_right_in[4] ) , 
    .X ( chanx_left_out[5] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_P_117 ( .A ( chany_bottom_in[2] ) , 
    .X ( chany_top_out[3] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_P_118 ( .A ( chany_bottom_in[5] ) , 
    .X ( chany_top_out[6] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_P_119 ( .A ( chany_bottom_in[12] ) , 
    .X ( chany_top_out[13] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_P_120 ( .A ( chany_bottom_in[14] ) , 
    .X ( chany_top_out[15] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_P_121 ( .A ( chany_bottom_in[16] ) , 
    .X ( chany_top_out[17] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 BUFT_P_122 ( .A ( aps_rename_2_ ) , 
    .X ( chanx_left_out[7] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 BUFT_P_123 ( .A ( aps_rename_3_ ) , 
    .X ( chanx_left_out[9] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_P_125 ( .A ( chanx_right_in[17] ) , 
    .X ( chanx_left_out[18] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_P_127 ( .A ( chanx_left_in[4] ) , 
    .X ( ropt_net_158 ) ) ;
endmodule


module mux_tree_tapbuf_size10_mem ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_33__59 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_34 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size10 ( in , sram , sram_inv , out , p0 ) ;
input  [0:9] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

const1_34 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[6] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[8] ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[9] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
endmodule


module mux_tree_tapbuf_size6_mem_0_2 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd1_1 FTB_32__58 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size6_mem_6 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_31__57 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_31 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size6_0_2 ( in , sram , sram_inv , out , p0 ) ;
input  [0:5] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;

const1_31 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
endmodule


module const1_30_1 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size6_6 ( in , sram , sram_inv , out , p0 ) ;
input  [0:5] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;

const1_30_1 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_69 ( 
    .A ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .X ( out[0] ) ) ;
endmodule


module mux_tree_tapbuf_size14_mem_0 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_30__56 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size14_mem ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_29__55 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_29_1 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size14_0 ( in , sram , sram_inv , out , p0 ) ;
input  [0:13] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_10_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_11_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_12_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_13_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

const1_29_1 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_13_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_3_ ( .A0 ( in[7] ) , .A1 ( in[6] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_4_ ( .A0 ( in[9] ) , .A1 ( in[8] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_5_ ( .A0 ( in[11] ) , .A1 ( in[10] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_6_ ( .A0 ( in[13] ) , .A1 ( in[12] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_10_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_11_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_10_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_12_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_12_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_11_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_13_X[0] ) ) ;
endmodule


module const1_28_1 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size14 ( in , sram , sram_inv , out , p0 ) ;
input  [0:13] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_10_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_11_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_12_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

const1_28_1 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_3_ ( .A0 ( in[7] ) , .A1 ( in[6] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_4_ ( .A0 ( in[9] ) , .A1 ( in[8] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_5_ ( .A0 ( in[11] ) , .A1 ( in[10] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_6_ ( .A0 ( in[13] ) , .A1 ( in[12] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_10_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_11_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_10_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_12_X[0] ) ) ;
sky130_fd_sc_hd__mux2_8 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_12_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_11_X[0] ) , .S ( sram[3] ) , .X ( out[0] ) ) ;
endmodule


module mux_tree_tapbuf_size9_mem ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_28__54 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size9_mem_0 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_27__53 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_27_1 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size9 ( in , sram , sram_inv , out , p0 ) ;
input  [0:8] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;

const1_27_1 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[7] ) , .A1 ( in[6] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[8] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
endmodule


module const1_26_2 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size9_0 ( in , sram , sram_inv , out , p0 ) ;
input  [0:8] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;

const1_26_2 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[7] ) , .A1 ( in[6] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[8] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_13 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_26__52 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_3_2 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_25__51 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_2_2 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_24__50 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_1_2 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_23__49 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_0_2 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_22__48 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_25_2 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_13 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_25_2 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
endmodule


module const1_24_2 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_3_2 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_24_2 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
endmodule


module const1_23_2 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_2_2 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_23_2 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_66 ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
endmodule


module const1_22_2 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_1_2 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_22_2 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
endmodule


module const1_21_2 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_0_2 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_21_2 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
endmodule


module mux_tree_tapbuf_size3_mem_7 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_21__47 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size3_mem_6 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_20__46 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size3_mem_5 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_19__45 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size3_mem_4 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_18__44 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size3_mem_3_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_17__43 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size3_mem_2_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_16__42 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size3_mem_1_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_15__41 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size3_mem_0_2 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_14__40 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_20_2 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size3_7 ( in , sram , sram_inv , out , p0 ) ;
input  [0:2] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;

const1_20_2 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( p0 ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
endmodule


module const1_19_2 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size3_6 ( in , sram , sram_inv , out , p0 ) ;
input  [0:2] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;

const1_19_2 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( p0 ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
endmodule


module const1_18_2 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size3_5 ( in , sram , sram_inv , out , p0 ) ;
input  [0:2] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;

const1_18_2 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( p0 ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
endmodule


module const1_17_2 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size3_4 ( in , sram , sram_inv , out , p0 ) ;
input  [0:2] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;

const1_17_2 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( p0 ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_105 ( 
    .A ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .X ( out[0] ) ) ;
endmodule


module const1_16_3 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size3_3_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:2] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;

const1_16_3 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( p0 ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
endmodule


module const1_15_3 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size3_2_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:2] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;

const1_15_3 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( p0 ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
endmodule


module const1_14_3 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size3_1_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:2] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;

const1_14_3 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( p0 ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
endmodule


module const1_13_3 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size3_0_2 ( in , sram , sram_inv , out , p0 ) ;
input  [0:2] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;

const1_13_3 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( p0 ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
endmodule


module mux_tree_tapbuf_size4_mem_0_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_13__39 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size4_mem_6 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_12__38 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_12_3 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size4_0_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:3] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;

const1_12_3 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( in[2] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , .A1 ( in[3] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
endmodule


module const1_11_3 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size4_6 ( in , sram , sram_inv , out , p0 ) ;
input  [0:3] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;

const1_11_3 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( in[2] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , .A1 ( in[3] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
endmodule


module mux_tree_tapbuf_size7_mem_1_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_11__37 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size7_mem_0_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_10__36 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size7_mem_3 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_9__35 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size7_mem_2 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_8__34 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size7_mem_2 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_7__33 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size7_mem_5 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_6__32 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size7_mem_4 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_5__31 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_10_3 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size7_1_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:6] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;

const1_10_3 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_3_ ( .A0 ( p0 ) , .A1 ( in[6] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
endmodule


module const1_9_3 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size7_0_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:6] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;

const1_9_3 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_3_ ( .A0 ( p0 ) , .A1 ( in[6] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
endmodule


module const1_8_3 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size7_3 ( in , sram , sram_inv , out , p0 ) ;
input  [0:6] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;

const1_8_3 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_3_ ( .A0 ( p0 ) , .A1 ( in[6] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
endmodule


module const1_7_3 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size7_2 ( in , sram , sram_inv , out , p0 ) ;
input  [0:6] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;

const1_7_3 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_3_ ( .A0 ( p0 ) , .A1 ( in[6] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
endmodule


module const1_6_4 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size7_2 ( in , sram , sram_inv , out , p0 ) ;
input  [0:6] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;

const1_6_4 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_3_ ( .A0 ( p0 ) , .A1 ( in[6] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_61 ( 
    .A ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , .X ( BUF_net_61 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 BUFT_P_104 ( .A ( BUF_net_61 ) , 
    .X ( out[0] ) ) ;
endmodule


module const1_5_4 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size7_5 ( in , sram , sram_inv , out , p0 ) ;
input  [0:6] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;

const1_5_4 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_3_ ( .A0 ( p0 ) , .A1 ( in[6] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
endmodule


module const1_4_4 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size7_4 ( in , sram , sram_inv , out , p0 ) ;
input  [0:6] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;

const1_4_4 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_3_ ( .A0 ( p0 ) , .A1 ( in[6] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
endmodule


module mux_tree_tapbuf_size8_mem_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_4__30 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size8_mem_0 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_3__29 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size8_mem_2 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_2__28 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size8_mem ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:3] mem_out ;
output [0:3] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_1__27 ( .A ( mem_out[3] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_3_4 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size8_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:7] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;

const1_3_4 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( in[2] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[4] ) , .A1 ( in[3] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[6] ) , .A1 ( in[5] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
endmodule


module const1_2_4 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size8_0 ( in , sram , sram_inv , out , p0 ) ;
input  [0:7] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;

const1_2_4 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( in[2] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[4] ) , .A1 ( in[3] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[6] ) , .A1 ( in[5] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
endmodule


module const1_1_4 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size8_2 ( in , sram , sram_inv , out , p0 ) ;
input  [0:7] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;

const1_1_4 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( in[2] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[4] ) , .A1 ( in[3] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[6] ) , .A1 ( in[5] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
endmodule


module const1_0_4 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size8 ( in , sram , sram_inv , out , p0 ) ;
input  [0:7] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;

const1_0_4 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( in[2] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( in[4] ) , .A1 ( in[3] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( .A0 ( in[6] ) , .A1 ( in[5] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( .A0 ( p0 ) , .A1 ( in[7] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
endmodule


module sb_1__0_ ( prog_clk , chany_top_in , top_left_grid_pin_34_ , 
    top_left_grid_pin_35_ , top_left_grid_pin_36_ , top_left_grid_pin_37_ , 
    top_left_grid_pin_38_ , top_left_grid_pin_39_ , top_left_grid_pin_40_ , 
    top_left_grid_pin_41_ , chanx_right_in , right_top_grid_pin_42_ , 
    right_top_grid_pin_43_ , right_top_grid_pin_44_ , right_top_grid_pin_45_ , 
    right_top_grid_pin_46_ , right_top_grid_pin_47_ , right_top_grid_pin_48_ , 
    right_top_grid_pin_49_ , right_bottom_grid_pin_1_ , chanx_left_in , 
    left_top_grid_pin_42_ , left_top_grid_pin_43_ , left_top_grid_pin_44_ , 
    left_top_grid_pin_45_ , left_top_grid_pin_46_ , left_top_grid_pin_47_ , 
    left_top_grid_pin_48_ , left_top_grid_pin_49_ , left_bottom_grid_pin_1_ , 
    ccff_head , chany_top_out , chanx_right_out , chanx_left_out , ccff_tail ) ;
input  [0:0] prog_clk ;
input  [0:19] chany_top_in ;
input  [0:0] top_left_grid_pin_34_ ;
input  [0:0] top_left_grid_pin_35_ ;
input  [0:0] top_left_grid_pin_36_ ;
input  [0:0] top_left_grid_pin_37_ ;
input  [0:0] top_left_grid_pin_38_ ;
input  [0:0] top_left_grid_pin_39_ ;
input  [0:0] top_left_grid_pin_40_ ;
input  [0:0] top_left_grid_pin_41_ ;
input  [0:19] chanx_right_in ;
input  [0:0] right_top_grid_pin_42_ ;
input  [0:0] right_top_grid_pin_43_ ;
input  [0:0] right_top_grid_pin_44_ ;
input  [0:0] right_top_grid_pin_45_ ;
input  [0:0] right_top_grid_pin_46_ ;
input  [0:0] right_top_grid_pin_47_ ;
input  [0:0] right_top_grid_pin_48_ ;
input  [0:0] right_top_grid_pin_49_ ;
input  [0:0] right_bottom_grid_pin_1_ ;
input  [0:19] chanx_left_in ;
input  [0:0] left_top_grid_pin_42_ ;
input  [0:0] left_top_grid_pin_43_ ;
input  [0:0] left_top_grid_pin_44_ ;
input  [0:0] left_top_grid_pin_45_ ;
input  [0:0] left_top_grid_pin_46_ ;
input  [0:0] left_top_grid_pin_47_ ;
input  [0:0] left_top_grid_pin_48_ ;
input  [0:0] left_top_grid_pin_49_ ;
input  [0:0] left_bottom_grid_pin_1_ ;
input  [0:0] ccff_head ;
output [0:19] chany_top_out ;
output [0:19] chanx_right_out ;
output [0:19] chanx_left_out ;
output [0:0] ccff_tail ;

wire [0:3] mux_tree_tapbuf_size10_0_sram ;
wire [0:3] mux_tree_tapbuf_size10_0_sram_inv ;
wire [0:0] mux_tree_tapbuf_size10_mem_0_ccff_tail ;
wire [0:3] mux_tree_tapbuf_size14_0_sram ;
wire [0:3] mux_tree_tapbuf_size14_0_sram_inv ;
wire [0:3] mux_tree_tapbuf_size14_1_sram ;
wire [0:3] mux_tree_tapbuf_size14_1_sram_inv ;
wire [0:0] mux_tree_tapbuf_size14_mem_0_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size14_mem_1_ccff_tail ;
wire [0:1] mux_tree_tapbuf_size2_0_sram ;
wire [0:1] mux_tree_tapbuf_size2_0_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_1_sram ;
wire [0:1] mux_tree_tapbuf_size2_1_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_2_sram ;
wire [0:1] mux_tree_tapbuf_size2_2_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_3_sram ;
wire [0:1] mux_tree_tapbuf_size2_3_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_4_sram ;
wire [0:1] mux_tree_tapbuf_size2_4_sram_inv ;
wire [0:0] mux_tree_tapbuf_size2_mem_0_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_1_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_2_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_3_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_4_ccff_tail ;
wire [0:1] mux_tree_tapbuf_size3_0_sram ;
wire [0:1] mux_tree_tapbuf_size3_0_sram_inv ;
wire [0:1] mux_tree_tapbuf_size3_1_sram ;
wire [0:1] mux_tree_tapbuf_size3_1_sram_inv ;
wire [0:1] mux_tree_tapbuf_size3_2_sram ;
wire [0:1] mux_tree_tapbuf_size3_2_sram_inv ;
wire [0:1] mux_tree_tapbuf_size3_3_sram ;
wire [0:1] mux_tree_tapbuf_size3_3_sram_inv ;
wire [0:1] mux_tree_tapbuf_size3_4_sram ;
wire [0:1] mux_tree_tapbuf_size3_4_sram_inv ;
wire [0:1] mux_tree_tapbuf_size3_5_sram ;
wire [0:1] mux_tree_tapbuf_size3_5_sram_inv ;
wire [0:1] mux_tree_tapbuf_size3_6_sram ;
wire [0:1] mux_tree_tapbuf_size3_6_sram_inv ;
wire [0:1] mux_tree_tapbuf_size3_7_sram ;
wire [0:1] mux_tree_tapbuf_size3_7_sram_inv ;
wire [0:0] mux_tree_tapbuf_size3_mem_0_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size3_mem_1_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size3_mem_2_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size3_mem_3_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size3_mem_4_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size3_mem_5_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size3_mem_6_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size3_mem_7_ccff_tail ;
wire [0:2] mux_tree_tapbuf_size4_0_sram ;
wire [0:2] mux_tree_tapbuf_size4_0_sram_inv ;
wire [0:2] mux_tree_tapbuf_size4_1_sram ;
wire [0:2] mux_tree_tapbuf_size4_1_sram_inv ;
wire [0:0] mux_tree_tapbuf_size4_mem_0_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size4_mem_1_ccff_tail ;
wire [0:2] mux_tree_tapbuf_size6_0_sram ;
wire [0:2] mux_tree_tapbuf_size6_0_sram_inv ;
wire [0:2] mux_tree_tapbuf_size6_1_sram ;
wire [0:2] mux_tree_tapbuf_size6_1_sram_inv ;
wire [0:0] mux_tree_tapbuf_size6_mem_0_ccff_tail ;
wire [0:2] mux_tree_tapbuf_size7_0_sram ;
wire [0:2] mux_tree_tapbuf_size7_0_sram_inv ;
wire [0:2] mux_tree_tapbuf_size7_1_sram ;
wire [0:2] mux_tree_tapbuf_size7_1_sram_inv ;
wire [0:2] mux_tree_tapbuf_size7_2_sram ;
wire [0:2] mux_tree_tapbuf_size7_2_sram_inv ;
wire [0:2] mux_tree_tapbuf_size7_3_sram ;
wire [0:2] mux_tree_tapbuf_size7_3_sram_inv ;
wire [0:2] mux_tree_tapbuf_size7_4_sram ;
wire [0:2] mux_tree_tapbuf_size7_4_sram_inv ;
wire [0:2] mux_tree_tapbuf_size7_5_sram ;
wire [0:2] mux_tree_tapbuf_size7_5_sram_inv ;
wire [0:2] mux_tree_tapbuf_size7_6_sram ;
wire [0:2] mux_tree_tapbuf_size7_6_sram_inv ;
wire [0:0] mux_tree_tapbuf_size7_mem_0_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size7_mem_1_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size7_mem_2_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size7_mem_3_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size7_mem_4_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size7_mem_5_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size7_mem_6_ccff_tail ;
wire [0:3] mux_tree_tapbuf_size8_0_sram ;
wire [0:3] mux_tree_tapbuf_size8_0_sram_inv ;
wire [0:3] mux_tree_tapbuf_size8_1_sram ;
wire [0:3] mux_tree_tapbuf_size8_1_sram_inv ;
wire [0:3] mux_tree_tapbuf_size8_2_sram ;
wire [0:3] mux_tree_tapbuf_size8_2_sram_inv ;
wire [0:3] mux_tree_tapbuf_size8_3_sram ;
wire [0:3] mux_tree_tapbuf_size8_3_sram_inv ;
wire [0:0] mux_tree_tapbuf_size8_mem_0_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size8_mem_1_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size8_mem_2_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size8_mem_3_ccff_tail ;
wire [0:3] mux_tree_tapbuf_size9_0_sram ;
wire [0:3] mux_tree_tapbuf_size9_0_sram_inv ;
wire [0:3] mux_tree_tapbuf_size9_1_sram ;
wire [0:3] mux_tree_tapbuf_size9_1_sram_inv ;
wire [0:0] mux_tree_tapbuf_size9_mem_0_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size9_mem_1_ccff_tail ;

mux_tree_tapbuf_size8 mux_top_track_0 (
    .in ( { top_left_grid_pin_34_[0] , top_left_grid_pin_36_[0] , 
        top_left_grid_pin_38_[0] , top_left_grid_pin_40_[0] , 
        chanx_right_in[1] , chanx_right_in[2] , chanx_left_in[0] , 
        chanx_left_in[2] } ) ,
    .sram ( mux_tree_tapbuf_size8_0_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size8_0_sram_inv ) , 
    .out ( chany_top_out[0] ) , .p0 ( optlc_net_124 ) ) ;
mux_tree_tapbuf_size8_2 mux_right_track_8 (
    .in ( { chany_top_in[2] , chany_top_in[9] , chany_top_in[16] , 
        right_top_grid_pin_42_[0] , right_top_grid_pin_46_[0] , 
        right_bottom_grid_pin_1_[0] , chanx_left_in[6] , chanx_left_in[16] } ) ,
    .sram ( mux_tree_tapbuf_size8_1_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size8_1_sram_inv ) , 
    .out ( chanx_right_out[4] ) , .p0 ( optlc_net_127 ) ) ;
mux_tree_tapbuf_size8_0 mux_left_track_3 (
    .in ( { chany_top_in[6] , chany_top_in[13] , chanx_right_in[4] , 
        chanx_right_in[13] , left_top_grid_pin_43_[0] , 
        left_top_grid_pin_45_[0] , left_top_grid_pin_47_[0] , 
        left_top_grid_pin_49_[0] } ) ,
    .sram ( mux_tree_tapbuf_size8_2_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size8_2_sram_inv ) , 
    .out ( chanx_left_out[1] ) , .p0 ( optlc_net_126 ) ) ;
mux_tree_tapbuf_size8_1 mux_left_track_9 (
    .in ( { chany_top_in[4] , chany_top_in[11] , chany_top_in[18] , 
        chanx_right_in[6] , chanx_right_in[16] , left_top_grid_pin_42_[0] , 
        left_top_grid_pin_46_[0] , left_bottom_grid_pin_1_[0] } ) ,
    .sram ( mux_tree_tapbuf_size8_3_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size8_3_sram_inv ) , 
    .out ( chanx_left_out[4] ) , .p0 ( optlc_net_126 ) ) ;
mux_tree_tapbuf_size8_mem mem_top_track_0 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( ccff_head ) , 
    .ccff_tail ( mux_tree_tapbuf_size8_mem_0_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size8_0_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size8_0_sram_inv ) ) ;
mux_tree_tapbuf_size8_mem_2 mem_right_track_8 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size14_mem_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size8_mem_1_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size8_1_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size8_1_sram_inv ) ) ;
mux_tree_tapbuf_size8_mem_0 mem_left_track_3 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size10_mem_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size8_mem_2_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size8_2_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size8_2_sram_inv ) ) ;
mux_tree_tapbuf_size8_mem_1 mem_left_track_9 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size14_mem_1_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size8_mem_3_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size8_3_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size8_3_sram_inv ) ) ;
mux_tree_tapbuf_size7_4 mux_top_track_2 (
    .in ( { top_left_grid_pin_35_[0] , top_left_grid_pin_37_[0] , 
        top_left_grid_pin_39_[0] , top_left_grid_pin_41_[0] , 
        chanx_right_in[3] , chanx_right_in[4] , chanx_left_in[4] } ) ,
    .sram ( mux_tree_tapbuf_size7_0_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size7_0_sram_inv ) , 
    .out ( chany_top_out[1] ) , .p0 ( optlc_net_124 ) ) ;
mux_tree_tapbuf_size7_5 mux_top_track_4 (
    .in ( { top_left_grid_pin_34_[0] , top_left_grid_pin_36_[0] , 
        top_left_grid_pin_38_[0] , top_left_grid_pin_40_[0] , 
        chanx_right_in[5] , chanx_right_in[7] , chanx_left_in[5] } ) ,
    .sram ( mux_tree_tapbuf_size7_1_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size7_1_sram_inv ) , 
    .out ( chany_top_out[2] ) , .p0 ( optlc_net_124 ) ) ;
mux_tree_tapbuf_size7_2 mux_top_track_6 (
    .in ( { top_left_grid_pin_35_[0] , top_left_grid_pin_37_[0] , 
        top_left_grid_pin_39_[0] , top_left_grid_pin_41_[0] , 
        chanx_right_in[6] , chanx_right_in[11] , chanx_left_in[6] } ) ,
    .sram ( mux_tree_tapbuf_size7_2_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size7_2_sram_inv ) ,
    .out ( { ropt_net_169 } ) ,
    .p0 ( optlc_net_127 ) ) ;
mux_tree_tapbuf_size7_2 mux_right_track_16 (
    .in ( { chany_top_in[3] , chany_top_in[10] , chany_top_in[17] , 
        right_top_grid_pin_43_[0] , right_top_grid_pin_47_[0] , 
        chanx_left_in[8] , chanx_left_in[17] } ) ,
    .sram ( mux_tree_tapbuf_size7_3_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size7_3_sram_inv ) , 
    .out ( chanx_right_out[8] ) , .p0 ( optlc_net_127 ) ) ;
mux_tree_tapbuf_size7_3 mux_right_track_24 (
    .in ( { chany_top_in[4] , chany_top_in[11] , chany_top_in[18] , 
        right_top_grid_pin_44_[0] , right_top_grid_pin_48_[0] , 
        chanx_left_in[9] , chanx_left_in[18] } ) ,
    .sram ( mux_tree_tapbuf_size7_4_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size7_4_sram_inv ) , 
    .out ( chanx_right_out[12] ) , .p0 ( optlc_net_127 ) ) ;
mux_tree_tapbuf_size7_0_1 mux_left_track_17 (
    .in ( { chany_top_in[3] , chany_top_in[10] , chany_top_in[17] , 
        chanx_right_in[8] , chanx_right_in[17] , left_top_grid_pin_43_[0] , 
        left_top_grid_pin_47_[0] } ) ,
    .sram ( mux_tree_tapbuf_size7_5_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size7_5_sram_inv ) , 
    .out ( chanx_left_out[8] ) , .p0 ( optlc_net_126 ) ) ;
mux_tree_tapbuf_size7_1_1 mux_left_track_25 (
    .in ( { chany_top_in[2] , chany_top_in[9] , chany_top_in[16] , 
        chanx_right_in[9] , chanx_right_in[18] , left_top_grid_pin_44_[0] , 
        left_top_grid_pin_48_[0] } ) ,
    .sram ( mux_tree_tapbuf_size7_6_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size7_6_sram_inv ) , 
    .out ( chanx_left_out[12] ) , .p0 ( optlc_net_126 ) ) ;
mux_tree_tapbuf_size7_mem_4 mem_top_track_2 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size8_mem_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size7_mem_0_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size7_0_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size7_0_sram_inv ) ) ;
mux_tree_tapbuf_size7_mem_5 mem_top_track_4 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size7_mem_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size7_mem_1_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size7_1_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size7_1_sram_inv ) ) ;
mux_tree_tapbuf_size7_mem_2 mem_top_track_6 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size7_mem_1_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size7_mem_2_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size7_2_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size7_2_sram_inv ) ) ;
mux_tree_tapbuf_size7_mem_2 mem_right_track_16 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size8_mem_1_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size7_mem_3_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size7_3_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size7_3_sram_inv ) ) ;
mux_tree_tapbuf_size7_mem_3 mem_right_track_24 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size7_mem_3_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size7_mem_4_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size7_4_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size7_4_sram_inv ) ) ;
mux_tree_tapbuf_size7_mem_0_1 mem_left_track_17 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size8_mem_3_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size7_mem_5_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size7_5_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size7_5_sram_inv ) ) ;
mux_tree_tapbuf_size7_mem_1_1 mem_left_track_25 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size7_mem_5_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size7_mem_6_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size7_6_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size7_6_sram_inv ) ) ;
mux_tree_tapbuf_size4_6 mux_top_track_8 (
    .in ( { top_left_grid_pin_34_[0] , chanx_right_in[8] , 
        chanx_right_in[15] , chanx_left_in[8] } ) ,
    .sram ( mux_tree_tapbuf_size4_0_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size4_0_sram_inv ) , 
    .out ( chany_top_out[4] ) , .p0 ( optlc_net_127 ) ) ;
mux_tree_tapbuf_size4_0_1 mux_top_track_10 (
    .in ( { top_left_grid_pin_35_[0] , chanx_right_in[9] , 
        chanx_right_in[19] , chanx_left_in[9] } ) ,
    .sram ( mux_tree_tapbuf_size4_1_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size4_1_sram_inv ) , 
    .out ( chany_top_out[5] ) , .p0 ( optlc_net_127 ) ) ;
mux_tree_tapbuf_size4_mem_6 mem_top_track_8 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size7_mem_2_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size4_mem_0_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size4_0_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size4_0_sram_inv ) ) ;
mux_tree_tapbuf_size4_mem_0_1 mem_top_track_10 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size4_mem_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size4_mem_1_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size4_1_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size4_1_sram_inv ) ) ;
mux_tree_tapbuf_size3_0_2 mux_top_track_12 (
    .in ( { top_left_grid_pin_36_[0] , chanx_right_in[10] , 
        chanx_left_in[10] } ) ,
    .sram ( mux_tree_tapbuf_size3_0_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size3_0_sram_inv ) , 
    .out ( chany_top_out[6] ) , .p0 ( optlc_net_125 ) ) ;
mux_tree_tapbuf_size3_1_1 mux_top_track_14 (
    .in ( { top_left_grid_pin_37_[0] , chanx_right_in[12] , 
        chanx_left_in[12] } ) ,
    .sram ( mux_tree_tapbuf_size3_1_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size3_1_sram_inv ) , 
    .out ( chany_top_out[7] ) , .p0 ( optlc_net_125 ) ) ;
mux_tree_tapbuf_size3_2_1 mux_top_track_16 (
    .in ( { top_left_grid_pin_38_[0] , chanx_right_in[13] , 
        chanx_left_in[13] } ) ,
    .sram ( mux_tree_tapbuf_size3_2_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size3_2_sram_inv ) , 
    .out ( chany_top_out[8] ) , .p0 ( optlc_net_125 ) ) ;
mux_tree_tapbuf_size3_3_1 mux_top_track_18 (
    .in ( { top_left_grid_pin_39_[0] , chanx_right_in[14] , 
        chanx_left_in[14] } ) ,
    .sram ( mux_tree_tapbuf_size3_3_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size3_3_sram_inv ) , 
    .out ( chany_top_out[9] ) , .p0 ( optlc_net_125 ) ) ;
mux_tree_tapbuf_size3_4 mux_top_track_20 (
    .in ( { top_left_grid_pin_40_[0] , chanx_right_in[16] , 
        chanx_left_in[16] } ) ,
    .sram ( mux_tree_tapbuf_size3_4_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size3_4_sram_inv ) ,
    .out ( { ropt_net_134 } ) ,
    .p0 ( optlc_net_124 ) ) ;
mux_tree_tapbuf_size3_5 mux_top_track_22 (
    .in ( { top_left_grid_pin_41_[0] , chanx_right_in[17] , 
        chanx_left_in[17] } ) ,
    .sram ( mux_tree_tapbuf_size3_5_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size3_5_sram_inv ) , 
    .out ( chany_top_out[11] ) , .p0 ( optlc_net_124 ) ) ;
mux_tree_tapbuf_size3_6 mux_top_track_24 (
    .in ( { top_left_grid_pin_34_[0] , chanx_right_in[18] , 
        chanx_left_in[18] } ) ,
    .sram ( mux_tree_tapbuf_size3_6_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size3_6_sram_inv ) , 
    .out ( chany_top_out[12] ) , .p0 ( optlc_net_124 ) ) ;
mux_tree_tapbuf_size3_7 mux_top_track_38 (
    .in ( { top_left_grid_pin_41_[0] , chanx_right_in[0] , chanx_left_in[1] } ) ,
    .sram ( mux_tree_tapbuf_size3_7_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size3_7_sram_inv ) , 
    .out ( chany_top_out[19] ) , .p0 ( optlc_net_125 ) ) ;
mux_tree_tapbuf_size3_mem_0_2 mem_top_track_12 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size4_mem_1_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size3_mem_0_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size3_0_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size3_0_sram_inv ) ) ;
mux_tree_tapbuf_size3_mem_1_1 mem_top_track_14 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size3_mem_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size3_mem_1_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size3_1_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size3_1_sram_inv ) ) ;
mux_tree_tapbuf_size3_mem_2_1 mem_top_track_16 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size3_mem_1_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size3_mem_2_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size3_2_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size3_2_sram_inv ) ) ;
mux_tree_tapbuf_size3_mem_3_1 mem_top_track_18 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size3_mem_2_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size3_mem_3_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size3_3_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size3_3_sram_inv ) ) ;
mux_tree_tapbuf_size3_mem_4 mem_top_track_20 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size3_mem_3_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size3_mem_4_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size3_4_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size3_4_sram_inv ) ) ;
mux_tree_tapbuf_size3_mem_5 mem_top_track_22 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size3_mem_4_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size3_mem_5_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size3_5_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size3_5_sram_inv ) ) ;
mux_tree_tapbuf_size3_mem_6 mem_top_track_24 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size3_mem_5_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size3_mem_6_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size3_6_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size3_6_sram_inv ) ) ;
mux_tree_tapbuf_size3_mem_7 mem_top_track_38 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_4_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size3_mem_7_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size3_7_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size3_7_sram_inv ) ) ;
mux_tree_tapbuf_size2_0_2 mux_top_track_28 (
    .in ( { top_left_grid_pin_36_[0] , chanx_left_in[19] } ) ,
    .sram ( mux_tree_tapbuf_size2_0_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_0_sram_inv ) , 
    .out ( chany_top_out[14] ) , .p0 ( optlc_net_125 ) ) ;
mux_tree_tapbuf_size2_1_2 mux_top_track_30 (
    .in ( { top_left_grid_pin_37_[0] , chanx_left_in[15] } ) ,
    .sram ( mux_tree_tapbuf_size2_1_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_1_sram_inv ) , 
    .out ( chany_top_out[15] ) , .p0 ( optlc_net_125 ) ) ;
mux_tree_tapbuf_size2_2_2 mux_top_track_32 (
    .in ( { top_left_grid_pin_38_[0] , chanx_left_in[11] } ) ,
    .sram ( mux_tree_tapbuf_size2_2_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_2_sram_inv ) ,
    .out ( { ropt_net_130 } ) ,
    .p0 ( optlc_net_125 ) ) ;
mux_tree_tapbuf_size2_3_2 mux_top_track_34 (
    .in ( { top_left_grid_pin_39_[0] , chanx_left_in[7] } ) ,
    .sram ( mux_tree_tapbuf_size2_3_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_3_sram_inv ) , 
    .out ( chany_top_out[17] ) , .p0 ( optlc_net_125 ) ) ;
mux_tree_tapbuf_size2_13 mux_top_track_36 (
    .in ( { top_left_grid_pin_40_[0] , chanx_left_in[3] } ) ,
    .sram ( mux_tree_tapbuf_size2_4_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_4_sram_inv ) , 
    .out ( chany_top_out[18] ) , .p0 ( optlc_net_125 ) ) ;
mux_tree_tapbuf_size2_mem_0_2 mem_top_track_28 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size3_mem_6_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_0_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_0_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_0_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem_1_2 mem_top_track_30 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_1_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_1_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_1_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem_2_2 mem_top_track_32 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_1_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_2_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_2_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_2_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem_3_2 mem_top_track_34 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_2_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_3_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_3_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_3_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem_13 mem_top_track_36 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_3_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_4_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_4_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_4_sram_inv ) ) ;
mux_tree_tapbuf_size9_0 mux_right_track_0 (
    .in ( { chany_top_in[6] , chany_top_in[13] , right_top_grid_pin_42_[0] , 
        right_top_grid_pin_44_[0] , right_top_grid_pin_46_[0] , 
        right_top_grid_pin_48_[0] , right_bottom_grid_pin_1_[0] , 
        chanx_left_in[2] , chanx_left_in[12] } ) ,
    .sram ( mux_tree_tapbuf_size9_0_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size9_0_sram_inv ) , 
    .out ( chanx_right_out[0] ) , .p0 ( optlc_net_127 ) ) ;
mux_tree_tapbuf_size9 mux_right_track_2 (
    .in ( { chany_top_in[0] , chany_top_in[7] , chany_top_in[14] , 
        right_top_grid_pin_43_[0] , right_top_grid_pin_45_[0] , 
        right_top_grid_pin_47_[0] , right_top_grid_pin_49_[0] , 
        chanx_left_in[4] , chanx_left_in[13] } ) ,
    .sram ( mux_tree_tapbuf_size9_1_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size9_1_sram_inv ) , 
    .out ( chanx_right_out[1] ) , .p0 ( optlc_net_125 ) ) ;
mux_tree_tapbuf_size9_mem_0 mem_right_track_0 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size3_mem_7_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size9_mem_0_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size9_0_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size9_0_sram_inv ) ) ;
mux_tree_tapbuf_size9_mem mem_right_track_2 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size9_mem_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size9_mem_1_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size9_1_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size9_1_sram_inv ) ) ;
mux_tree_tapbuf_size14 mux_right_track_4 (
    .in ( { chany_top_in[1] , chany_top_in[8] , chany_top_in[15] , 
        right_top_grid_pin_42_[0] , right_top_grid_pin_43_[0] , 
        right_top_grid_pin_44_[0] , right_top_grid_pin_45_[0] , 
        right_top_grid_pin_46_[0] , right_top_grid_pin_47_[0] , 
        right_top_grid_pin_48_[0] , right_top_grid_pin_49_[0] , 
        right_bottom_grid_pin_1_[0] , chanx_left_in[5] , chanx_left_in[14] } ) ,
    .sram ( mux_tree_tapbuf_size14_0_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size14_0_sram_inv ) , 
    .out ( chanx_right_out[2] ) , .p0 ( optlc_net_127 ) ) ;
mux_tree_tapbuf_size14_0 mux_left_track_5 (
    .in ( { chany_top_in[5] , chany_top_in[12] , chany_top_in[19] , 
        chanx_right_in[5] , chanx_right_in[14] , left_top_grid_pin_42_[0] , 
        left_top_grid_pin_43_[0] , left_top_grid_pin_44_[0] , 
        left_top_grid_pin_45_[0] , left_top_grid_pin_46_[0] , 
        left_top_grid_pin_47_[0] , left_top_grid_pin_48_[0] , 
        left_top_grid_pin_49_[0] , left_bottom_grid_pin_1_[0] } ) ,
    .sram ( mux_tree_tapbuf_size14_1_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size14_1_sram_inv ) , 
    .out ( chanx_left_out[2] ) , .p0 ( optlc_net_126 ) ) ;
mux_tree_tapbuf_size14_mem mem_right_track_4 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size9_mem_1_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size14_mem_0_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size14_0_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size14_0_sram_inv ) ) ;
mux_tree_tapbuf_size14_mem_0 mem_left_track_5 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size8_mem_2_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size14_mem_1_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size14_1_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size14_1_sram_inv ) ) ;
mux_tree_tapbuf_size6_6 mux_right_track_32 (
    .in ( { chany_top_in[5] , chany_top_in[12] , chany_top_in[19] , 
        right_top_grid_pin_45_[0] , right_top_grid_pin_49_[0] , 
        chanx_left_in[10] } ) ,
    .sram ( mux_tree_tapbuf_size6_0_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size6_0_sram_inv ) ,
    .out ( { ropt_net_129 } ) ,
    .p0 ( optlc_net_125 ) ) ;
mux_tree_tapbuf_size6_0_2 mux_left_track_33 (
    .in ( { chany_top_in[1] , chany_top_in[8] , chany_top_in[15] , 
        chanx_right_in[10] , left_top_grid_pin_45_[0] , 
        left_top_grid_pin_49_[0] } ) ,
    .sram ( mux_tree_tapbuf_size6_1_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size6_1_sram_inv ) , 
    .out ( chanx_left_out[16] ) , .p0 ( optlc_net_126 ) ) ;
mux_tree_tapbuf_size6_mem_6 mem_right_track_32 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size7_mem_4_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size6_mem_0_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size6_0_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size6_0_sram_inv ) ) ;
mux_tree_tapbuf_size6_mem_0_2 mem_left_track_33 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size7_mem_6_ccff_tail ) ,
    .ccff_tail ( { ropt_net_131 } ) ,
    .mem_out ( mux_tree_tapbuf_size6_1_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size6_1_sram_inv ) ) ;
mux_tree_tapbuf_size10 mux_left_track_1 (
    .in ( { chany_top_in[0] , chany_top_in[7] , chany_top_in[14] , 
        chanx_right_in[2] , chanx_right_in[12] , left_top_grid_pin_42_[0] , 
        left_top_grid_pin_44_[0] , left_top_grid_pin_46_[0] , 
        left_top_grid_pin_48_[0] , left_bottom_grid_pin_1_[0] } ) ,
    .sram ( mux_tree_tapbuf_size10_0_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size10_0_sram_inv ) , 
    .out ( chanx_left_out[0] ) , .p0 ( optlc_net_126 ) ) ;
mux_tree_tapbuf_size10_mem mem_left_track_1 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size6_mem_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size10_mem_0_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size10_0_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size10_0_sram_inv ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_1__0 ( .A ( top_left_grid_pin_35_[0] ) , 
    .X ( ropt_net_150 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_115 ( .LO ( SYNOPSYS_UNCONNECTED_1 ) , 
    .HI ( optlc_net_124 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_745 ( .A ( ropt_net_155 ) , 
    .X ( chanx_left_out[6] ) ) ;
sky130_fd_sc_hd__conb_1 optlc_117 ( .LO ( SYNOPSYS_UNCONNECTED_2 ) , 
    .HI ( optlc_net_125 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_119 ( .LO ( SYNOPSYS_UNCONNECTED_3 ) , 
    .HI ( optlc_net_126 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_6__5 ( .A ( chanx_right_in[8] ) , 
    .X ( ropt_net_136 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_121 ( .LO ( SYNOPSYS_UNCONNECTED_4 ) , 
    .HI ( optlc_net_127 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_716 ( .A ( chanx_right_in[16] ) , 
    .X ( chanx_left_out[17] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_9__8 ( .A ( chanx_right_in[12] ) , 
    .X ( chanx_left_out[13] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_717 ( .A ( ropt_net_129 ) , 
    .X ( ropt_net_161 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_11__10 ( .A ( chanx_right_in[14] ) , 
    .X ( chanx_left_out[15] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_718 ( .A ( ropt_net_130 ) , 
    .X ( ropt_net_167 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_13__12 ( .A ( chanx_right_in[17] ) , 
    .X ( chanx_left_out[18] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_14__13 ( .A ( chanx_right_in[18] ) , 
    .X ( chanx_left_out[19] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_15__14 ( .A ( chanx_left_in[2] ) , 
    .X ( ropt_net_149 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_16__15 ( .A ( chanx_left_in[4] ) , 
    .X ( ropt_net_145 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_17__16 ( .A ( chanx_left_in[5] ) , 
    .X ( chanx_right_out[6] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_719 ( .A ( ropt_net_131 ) , 
    .X ( ropt_net_157 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_746 ( .A ( ropt_net_156 ) , 
    .X ( chanx_left_out[9] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_20__19 ( .A ( chanx_left_in[9] ) , 
    .X ( ropt_net_141 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_21__20 ( .A ( chanx_left_in[10] ) , 
    .X ( chanx_right_out[11] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_720 ( .A ( ropt_net_132 ) , 
    .X ( chanx_right_out[9] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_721 ( .A ( chanx_right_in[2] ) , 
    .X ( chanx_left_out[3] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_747 ( .A ( ropt_net_157 ) , 
    .X ( ccff_tail[0] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_722 ( .A ( ropt_net_134 ) , 
    .X ( ropt_net_170 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_723 ( .A ( chanx_right_in[6] ) , 
    .X ( ropt_net_172 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_724 ( .A ( ropt_net_136 ) , 
    .X ( ropt_net_156 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_748 ( .A ( ropt_net_158 ) , 
    .X ( chanx_left_out[5] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_749 ( .A ( ropt_net_159 ) , 
    .X ( chanx_right_out[14] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_750 ( .A ( ropt_net_160 ) , 
    .X ( chanx_right_out[15] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_751 ( .A ( ropt_net_161 ) , 
    .X ( chanx_right_out[16] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_74 ( .A ( chanx_right_in[13] ) , 
    .X ( ropt_net_148 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_752 ( .A ( ropt_net_162 ) , 
    .X ( chanx_right_out[7] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_76 ( .A ( chanx_left_in[6] ) , 
    .X ( ropt_net_140 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 BUFT_RR_77 ( .A ( chanx_left_in[8] ) , 
    .X ( ropt_net_132 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_725 ( .A ( chanx_left_in[13] ) , 
    .X ( ropt_net_159 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_RR_79 ( .A ( chanx_left_in[16] ) , 
    .X ( ropt_net_142 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_80 ( .A ( chanx_left_in[17] ) , 
    .X ( ropt_net_147 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_726 ( .A ( chanx_right_in[9] ) , 
    .X ( chanx_left_out[10] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_RR_83 ( .A ( chanx_left_in[12] ) , 
    .X ( ropt_net_146 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_RR_84 ( .A ( chanx_left_in[18] ) , 
    .X ( ropt_net_144 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_727 ( .A ( chanx_left_in[14] ) , 
    .X ( ropt_net_160 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_728 ( .A ( ropt_net_140 ) , 
    .X ( ropt_net_162 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_729 ( .A ( ropt_net_141 ) , 
    .X ( ropt_net_168 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_730 ( .A ( ropt_net_142 ) , 
    .X ( chanx_right_out[17] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_731 ( .A ( chanx_right_in[4] ) , 
    .X ( ropt_net_158 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_P_100 ( .A ( chanx_right_in[10] ) , 
    .X ( ropt_net_171 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_733 ( .A ( ropt_net_144 ) , 
    .X ( chanx_right_out[19] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_753 ( .A ( ropt_net_163 ) , 
    .X ( chanx_right_out[18] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_755 ( .A ( ropt_net_164 ) , 
    .X ( chany_top_out[13] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_735 ( .A ( ropt_net_145 ) , 
    .X ( chanx_right_out[5] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_756 ( .A ( ropt_net_165 ) , 
    .X ( chanx_right_out[3] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_737 ( .A ( ropt_net_146 ) , 
    .X ( chanx_right_out[13] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_738 ( .A ( ropt_net_147 ) , 
    .X ( ropt_net_163 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_739 ( .A ( ropt_net_148 ) , 
    .X ( ropt_net_166 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_741 ( .A ( ropt_net_149 ) , 
    .X ( ropt_net_165 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_743 ( .A ( ropt_net_150 ) , 
    .X ( ropt_net_164 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_744 ( .A ( chanx_right_in[5] ) , 
    .X ( ropt_net_155 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_759 ( .A ( ropt_net_166 ) , 
    .X ( chanx_left_out[14] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_760 ( .A ( ropt_net_167 ) , 
    .X ( chany_top_out[16] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_761 ( .A ( ropt_net_168 ) , 
    .X ( chanx_right_out[10] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_762 ( .A ( ropt_net_169 ) , 
    .X ( chany_top_out[3] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_763 ( .A ( ropt_net_170 ) , 
    .X ( chany_top_out[10] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_764 ( .A ( ropt_net_171 ) , 
    .X ( chanx_left_out[11] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_765 ( .A ( ropt_net_172 ) , 
    .X ( chanx_left_out[7] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_1_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_8__39 ( .A ( mem_out[1] ) , 
    .X ( net_net_71 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_90 ( .A ( net_net_71 ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_3_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_7__38 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_2_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_6__37 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_0_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_5__36 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_5_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_4__35 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_12 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_3__34 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_6_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_2__33 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_4_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_1__32 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_33 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_1_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_33 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
endmodule


module const1_6_3 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_3_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_6_3 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
endmodule


module const1_5_3 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_2_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_5_3 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
endmodule


module const1_4_3 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_0_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_4_3 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
endmodule


module const1_3_3 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_5_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_3_3 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
endmodule


module const1_2_3 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_12 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_2_3 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
endmodule


module const1_1_3 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_6_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_1_3 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
endmodule


module const1_0_3 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_4_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_0_3 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
endmodule


module sb_0__2_ ( prog_clk , chanx_right_in , right_top_grid_pin_1_ , 
    chany_bottom_in , bottom_left_grid_pin_1_ , ccff_head , chanx_right_out , 
    chany_bottom_out , ccff_tail ) ;
input  [0:0] prog_clk ;
input  [0:19] chanx_right_in ;
input  [0:0] right_top_grid_pin_1_ ;
input  [0:19] chany_bottom_in ;
input  [0:0] bottom_left_grid_pin_1_ ;
input  [0:0] ccff_head ;
output [0:19] chanx_right_out ;
output [0:19] chany_bottom_out ;
output [0:0] ccff_tail ;

wire [0:1] mux_tree_tapbuf_size2_0_sram ;
wire [0:1] mux_tree_tapbuf_size2_0_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_1_sram ;
wire [0:1] mux_tree_tapbuf_size2_1_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_2_sram ;
wire [0:1] mux_tree_tapbuf_size2_2_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_3_sram ;
wire [0:1] mux_tree_tapbuf_size2_3_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_4_sram ;
wire [0:1] mux_tree_tapbuf_size2_4_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_5_sram ;
wire [0:1] mux_tree_tapbuf_size2_5_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_6_sram ;
wire [0:1] mux_tree_tapbuf_size2_6_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_7_sram ;
wire [0:1] mux_tree_tapbuf_size2_7_sram_inv ;
wire [0:0] mux_tree_tapbuf_size2_mem_0_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_1_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_2_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_3_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_4_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_5_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_6_ccff_tail ;

mux_tree_tapbuf_size2_4_1 mux_right_track_0 (
    .in ( { right_top_grid_pin_1_[0] , chany_bottom_in[18] } ) ,
    .sram ( mux_tree_tapbuf_size2_0_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_0_sram_inv ) , 
    .out ( chanx_right_out[0] ) , .p0 ( optlc_net_98 ) ) ;
mux_tree_tapbuf_size2_6_1 mux_right_track_4 (
    .in ( { right_top_grid_pin_1_[0] , chany_bottom_in[16] } ) ,
    .sram ( mux_tree_tapbuf_size2_1_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_1_sram_inv ) , 
    .out ( chanx_right_out[2] ) , .p0 ( optlc_net_98 ) ) ;
mux_tree_tapbuf_size2_12 mux_right_track_8 (
    .in ( { right_top_grid_pin_1_[0] , chany_bottom_in[14] } ) ,
    .sram ( mux_tree_tapbuf_size2_2_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_2_sram_inv ) , 
    .out ( chanx_right_out[4] ) , .p0 ( optlc_net_98 ) ) ;
mux_tree_tapbuf_size2_5_1 mux_right_track_24 (
    .in ( { right_top_grid_pin_1_[0] , chany_bottom_in[6] } ) ,
    .sram ( mux_tree_tapbuf_size2_3_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_3_sram_inv ) , 
    .out ( chanx_right_out[12] ) , .p0 ( optlc_net_98 ) ) ;
mux_tree_tapbuf_size2_0_1 mux_bottom_track_1 (
    .in ( { chanx_right_in[18] , bottom_left_grid_pin_1_[0] } ) ,
    .sram ( mux_tree_tapbuf_size2_4_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_4_sram_inv ) , 
    .out ( chany_bottom_out[0] ) , .p0 ( optlc_net_97 ) ) ;
mux_tree_tapbuf_size2_2_1 mux_bottom_track_5 (
    .in ( { chanx_right_in[16] , bottom_left_grid_pin_1_[0] } ) ,
    .sram ( mux_tree_tapbuf_size2_5_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_5_sram_inv ) , 
    .out ( chany_bottom_out[2] ) , .p0 ( optlc_net_97 ) ) ;
mux_tree_tapbuf_size2_3_1 mux_bottom_track_9 (
    .in ( { chanx_right_in[14] , bottom_left_grid_pin_1_[0] } ) ,
    .sram ( mux_tree_tapbuf_size2_6_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_6_sram_inv ) , 
    .out ( chany_bottom_out[4] ) , .p0 ( optlc_net_97 ) ) ;
mux_tree_tapbuf_size2_1_1 mux_bottom_track_25 (
    .in ( { chanx_right_in[6] , bottom_left_grid_pin_1_[0] } ) ,
    .sram ( mux_tree_tapbuf_size2_7_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_7_sram_inv ) , 
    .out ( chany_bottom_out[12] ) , .p0 ( optlc_net_97 ) ) ;
mux_tree_tapbuf_size2_mem_4_1 mem_right_track_0 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( ccff_head ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_0_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_0_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_0_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem_6_1 mem_right_track_4 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_1_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_1_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_1_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem_12 mem_right_track_8 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_1_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_2_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_2_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_2_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem_5_1 mem_right_track_24 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_2_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_3_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_3_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_3_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem_0_1 mem_bottom_track_1 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_3_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_4_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_4_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_4_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem_2_1 mem_bottom_track_5 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_4_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_5_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_5_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_5_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem_3_1 mem_bottom_track_9 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_5_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_6_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_6_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_6_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem_1_1 mem_bottom_track_25 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_6_ccff_tail ) ,
    .ccff_tail ( { ropt_net_103 } ) ,
    .mem_out ( mux_tree_tapbuf_size2_7_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_7_sram_inv ) ) ;
sky130_fd_sc_hd__conb_1 optlc_99 ( .LO ( SYNOPSYS_UNCONNECTED_1 ) , 
    .HI ( optlc_net_97 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_101 ( .LO ( SYNOPSYS_UNCONNECTED_2 ) , 
    .HI ( optlc_net_98 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_722 ( .A ( ropt_net_130 ) , 
    .X ( chany_bottom_out[13] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_723 ( .A ( ropt_net_131 ) , 
    .X ( chany_bottom_out[5] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_724 ( .A ( ropt_net_132 ) , 
    .X ( chany_bottom_out[3] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_725 ( .A ( ropt_net_133 ) , 
    .X ( chany_bottom_out[19] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_726 ( .A ( ropt_net_134 ) , 
    .X ( ccff_tail[0] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_690 ( .A ( chanx_right_in[15] ) , 
    .X ( ropt_net_132 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_691 ( .A ( chanx_right_in[19] ) , 
    .X ( ropt_net_133 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_727 ( .A ( ropt_net_135 ) , 
    .X ( chany_bottom_out[9] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_692 ( 
    .A ( chany_bottom_in[13] ) , .X ( ropt_net_154 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_728 ( .A ( ropt_net_136 ) , 
    .X ( chanx_right_out[10] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_693 ( .A ( ropt_net_102 ) , 
    .X ( ropt_net_130 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_694 ( .A ( ropt_net_103 ) , 
    .X ( ropt_net_134 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_729 ( .A ( ropt_net_137 ) , 
    .X ( chanx_right_out[1] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_695 ( .A ( chanx_right_in[4] ) , 
    .X ( ropt_net_155 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_696 ( .A ( chanx_right_in[10] ) , 
    .X ( ropt_net_150 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_697 ( .A ( chanx_right_in[12] ) , 
    .X ( ropt_net_151 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_698 ( .A ( chanx_right_in[3] ) , 
    .X ( chany_bottom_out[15] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_699 ( .A ( chanx_right_in[17] ) , 
    .X ( chany_bottom_out[1] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_700 ( .A ( chanx_right_in[7] ) , 
    .X ( chany_bottom_out[11] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_701 ( .A ( chany_bottom_in[4] ) , 
    .X ( ropt_net_153 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_702 ( 
    .A ( chany_bottom_in[11] ) , .X ( ropt_net_152 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_703 ( .A ( chany_bottom_in[5] ) , 
    .X ( chanx_right_out[13] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_704 ( .A ( ropt_net_113 ) , 
    .X ( ropt_net_140 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_705 ( .A ( ropt_net_114 ) , 
    .X ( ropt_net_136 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_706 ( .A ( chanx_right_in[9] ) , 
    .X ( ropt_net_135 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_707 ( .A ( ropt_net_116 ) , 
    .X ( chanx_right_out[8] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_708 ( .A ( ropt_net_117 ) , 
    .X ( ropt_net_137 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_709 ( .A ( ropt_net_118 ) , 
    .X ( chanx_right_out[17] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_710 ( .A ( ropt_net_119 ) , 
    .X ( chanx_right_out[16] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_712 ( .A ( ropt_net_120 ) , 
    .X ( ropt_net_143 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_713 ( .A ( ropt_net_121 ) , 
    .X ( ropt_net_131 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_714 ( .A ( ropt_net_122 ) , 
    .X ( ropt_net_142 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_42 ( .A ( chanx_right_in[2] ) , 
    .X ( BUF_net_42 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_730 ( .A ( ropt_net_138 ) , 
    .X ( chany_bottom_out[16] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_731 ( .A ( ropt_net_139 ) , 
    .X ( chanx_right_out[19] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_732 ( .A ( ropt_net_140 ) , 
    .X ( chanx_right_out[18] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_733 ( .A ( ropt_net_141 ) , 
    .X ( chany_bottom_out[17] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_47 ( .A ( chanx_right_in[8] ) , 
    .X ( ropt_net_125 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_734 ( .A ( ropt_net_142 ) , 
    .X ( chanx_right_out[6] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_715 ( .A ( ropt_net_123 ) , 
    .X ( ropt_net_144 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_735 ( .A ( ropt_net_143 ) , 
    .X ( chanx_right_out[3] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_716 ( .A ( ropt_net_124 ) , 
    .X ( ropt_net_145 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_736 ( .A ( ropt_net_144 ) , 
    .X ( chanx_right_out[11] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_737 ( .A ( ropt_net_145 ) , 
    .X ( chany_bottom_out[18] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_738 ( .A ( ropt_net_146 ) , 
    .X ( chanx_right_out[15] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_55 ( .A ( chany_bottom_in[0] ) , 
    .X ( ropt_net_113 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_RR_56 ( .A ( chany_bottom_in[1] ) , 
    .X ( ropt_net_118 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_RR_57 ( .A ( chany_bottom_in[2] ) , 
    .X ( ropt_net_119 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_58 ( .A ( chany_bottom_in[3] ) , 
    .X ( ropt_net_127 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_739 ( .A ( ropt_net_147 ) , 
    .X ( chanx_right_out[9] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_740 ( .A ( ropt_net_148 ) , 
    .X ( chany_bottom_out[10] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_61 ( .A ( chany_bottom_in[7] ) , 
    .X ( ropt_net_123 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_62 ( .A ( chany_bottom_in[8] ) , 
    .X ( ropt_net_114 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_63 ( .A ( chany_bottom_in[9] ) , 
    .X ( ropt_net_128 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_RR_64 ( .A ( chany_bottom_in[10] ) , 
    .X ( ropt_net_116 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_741 ( .A ( ropt_net_149 ) , 
    .X ( chany_bottom_out[7] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_717 ( .A ( ropt_net_125 ) , 
    .X ( ropt_net_148 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_67 ( .A ( chany_bottom_in[15] ) , 
    .X ( ropt_net_120 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_68 ( .A ( chany_bottom_in[17] ) , 
    .X ( ropt_net_117 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_718 ( .A ( ropt_net_126 ) , 
    .X ( ropt_net_139 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_719 ( .A ( ropt_net_127 ) , 
    .X ( ropt_net_146 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_720 ( .A ( ropt_net_128 ) , 
    .X ( ropt_net_147 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_721 ( .A ( ropt_net_129 ) , 
    .X ( ropt_net_141 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_742 ( .A ( ropt_net_150 ) , 
    .X ( chany_bottom_out[8] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_744 ( .A ( ropt_net_151 ) , 
    .X ( chany_bottom_out[6] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_745 ( .A ( ropt_net_152 ) , 
    .X ( chanx_right_out[7] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_746 ( .A ( ropt_net_153 ) , 
    .X ( chanx_right_out[14] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_748 ( .A ( ropt_net_154 ) , 
    .X ( chanx_right_out[5] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 BUFT_P_80 ( .A ( BUF_net_42 ) , 
    .X ( ropt_net_138 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_751 ( .A ( ropt_net_155 ) , 
    .X ( chany_bottom_out[14] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_P_83 ( .A ( chanx_right_in[5] ) , 
    .X ( ropt_net_102 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_P_86 ( .A ( chanx_right_in[11] ) , 
    .X ( ropt_net_149 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_P_88 ( .A ( chanx_right_in[13] ) , 
    .X ( ropt_net_121 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_P_91 ( .A ( chanx_right_in[0] ) , 
    .X ( ropt_net_124 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_P_92 ( .A ( chanx_right_in[1] ) , 
    .X ( ropt_net_129 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_P_95 ( .A ( chany_bottom_in[12] ) , 
    .X ( ropt_net_122 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_P_96 ( .A ( chany_bottom_in[19] ) , 
    .X ( ropt_net_126 ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_11 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_28__58 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_32 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_11 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_32 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
endmodule


module mux_tree_tapbuf_size3_mem_0_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd1_1 FTB_27__57 ( .A ( mem_out[1] ) , 
    .X ( net_net_101 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_101 ( .A ( net_net_101 ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size3_mem_4 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_26__56 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size3_mem_3 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_25__55 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size3_mem_2 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_24__54 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size3_mem_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_23__53 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_26_1 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size3_0_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:2] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;

const1_26_1 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( p0 ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
endmodule


module const1_25_1 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size3_4 ( in , sram , sram_inv , out , p0 ) ;
input  [0:2] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;

const1_25_1 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( p0 ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
endmodule


module const1_24_1 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size3_3 ( in , sram , sram_inv , out , p0 ) ;
input  [0:2] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;

const1_24_1 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( p0 ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
endmodule


module const1_23_1 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size3_2 ( in , sram , sram_inv , out , p0 ) ;
input  [0:2] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;

const1_23_1 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( p0 ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
endmodule


module const1_22_1 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size3_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:2] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;

const1_22_1 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( p0 ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
endmodule


module mux_tree_tapbuf_size7_mem ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_22__52 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size7_mem_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_21__51 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size7_mem_0 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_20__50 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_21_1 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size7 ( in , sram , sram_inv , out , p0 ) ;
input  [0:6] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;

const1_21_1 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_3_ ( .A0 ( p0 ) , .A1 ( in[6] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
endmodule


module const1_20_1 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size7_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:6] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;

const1_20_1 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_3_ ( .A0 ( p0 ) , .A1 ( in[6] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
endmodule


module const1_19_1 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size7_0 ( in , sram , sram_inv , out , p0 ) ;
input  [0:6] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;

const1_19_1 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_3_ ( .A0 ( p0 ) , .A1 ( in[6] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
endmodule


module mux_tree_tapbuf_size4_mem_3 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_19__49 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size4_mem_2 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_18__48 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size4_mem_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_17__47 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size4_mem_0 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_16__46 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size4_mem_4 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_15__45 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size4_mem ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_14__44 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size4_mem_5 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_13__43 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_18_1 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size4_3 ( in , sram , sram_inv , out , p0 ) ;
input  [0:3] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;

const1_18_1 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( in[2] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , .A1 ( in[3] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
endmodule


module const1_17_1 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size4_2 ( in , sram , sram_inv , out , p0 ) ;
input  [0:3] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;

const1_17_1 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( in[2] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , .A1 ( in[3] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
endmodule


module const1_16_2 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size4_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:3] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;

const1_16_2 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( in[2] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , .A1 ( in[3] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
endmodule


module const1_15_2 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size4_0 ( in , sram , sram_inv , out , p0 ) ;
input  [0:3] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;

const1_15_2 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( in[2] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , .A1 ( in[3] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
endmodule


module const1_14_2 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size4_4 ( in , sram , sram_inv , out , p0 ) ;
input  [0:3] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;

const1_14_2 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( in[2] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , .A1 ( in[3] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
endmodule


module const1_13_2 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size4 ( in , sram , sram_inv , out , p0 ) ;
input  [0:3] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;

const1_13_2 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( in[2] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , .A1 ( in[3] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
endmodule


module const1_12_2 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size4_5 ( in , sram , sram_inv , out , p0 ) ;
input  [0:3] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;

const1_12_2 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( in[2] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , .A1 ( in[3] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
endmodule


module mux_tree_tapbuf_size5_mem_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_12__42 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size5_mem_0_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_11__41 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size5_mem_2 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_10__40 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size5_mem_3 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_9__39 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size5_mem_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_8__38 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_11_2 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size5_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:4] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;

const1_11_2 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , .A1 ( in[4] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
endmodule


module const1_10_2 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size5_0_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:4] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;

const1_10_2 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , .A1 ( in[4] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
endmodule


module const1_9_2 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size5_2 ( in , sram , sram_inv , out , p0 ) ;
input  [0:4] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;

const1_9_2 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , .A1 ( in[4] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
endmodule


module const1_8_2 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size5_3 ( in , sram , sram_inv , out , p0 ) ;
input  [0:4] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;

const1_8_2 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , .A1 ( in[4] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
endmodule


module const1_7_2 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size5_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:4] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;

const1_7_2 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , .A1 ( in[4] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
endmodule


module mux_tree_tapbuf_size6_mem_2 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_7__37 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size6_mem_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_6__36 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size6_mem_0_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_5__35 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size6_mem_3 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_4__34 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size6_mem_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_3__33 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size6_mem_5 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_2__32 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size6_mem_4 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_1__31 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_6_2 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size6_2 ( in , sram , sram_inv , out , p0 ) ;
input  [0:5] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;

const1_6_2 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
endmodule


module const1_5_2 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size6_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:5] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;

const1_5_2 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
endmodule


module const1_4_2 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size6_0_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:5] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;

const1_4_2 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
endmodule


module const1_3_2 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size6_3 ( in , sram , sram_inv , out , p0 ) ;
input  [0:5] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;

const1_3_2 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
endmodule


module const1_2_2 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size6_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:5] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;

const1_2_2 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
endmodule


module const1_1_2 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size6_5 ( in , sram , sram_inv , out , p0 ) ;
input  [0:5] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;

const1_1_2 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
endmodule


module const1_0_2 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size6_4 ( in , sram , sram_inv , out , p0 ) ;
input  [0:5] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;

const1_0_2 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
endmodule


module sb_0__1_ ( prog_clk , chany_top_in , top_left_grid_pin_1_ , 
    chanx_right_in , right_top_grid_pin_42_ , right_top_grid_pin_43_ , 
    right_top_grid_pin_44_ , right_top_grid_pin_45_ , right_top_grid_pin_46_ , 
    right_top_grid_pin_47_ , right_top_grid_pin_48_ , right_top_grid_pin_49_ , 
    chany_bottom_in , bottom_left_grid_pin_1_ , ccff_head , chany_top_out , 
    chanx_right_out , chany_bottom_out , ccff_tail ) ;
input  [0:0] prog_clk ;
input  [0:19] chany_top_in ;
input  [0:0] top_left_grid_pin_1_ ;
input  [0:19] chanx_right_in ;
input  [0:0] right_top_grid_pin_42_ ;
input  [0:0] right_top_grid_pin_43_ ;
input  [0:0] right_top_grid_pin_44_ ;
input  [0:0] right_top_grid_pin_45_ ;
input  [0:0] right_top_grid_pin_46_ ;
input  [0:0] right_top_grid_pin_47_ ;
input  [0:0] right_top_grid_pin_48_ ;
input  [0:0] right_top_grid_pin_49_ ;
input  [0:19] chany_bottom_in ;
input  [0:0] bottom_left_grid_pin_1_ ;
input  [0:0] ccff_head ;
output [0:19] chany_top_out ;
output [0:19] chanx_right_out ;
output [0:19] chany_bottom_out ;
output [0:0] ccff_tail ;

wire [0:1] mux_tree_tapbuf_size2_0_sram ;
wire [0:1] mux_tree_tapbuf_size2_0_sram_inv ;
wire [0:0] mux_tree_tapbuf_size2_mem_0_ccff_tail ;
wire [0:1] mux_tree_tapbuf_size3_0_sram ;
wire [0:1] mux_tree_tapbuf_size3_0_sram_inv ;
wire [0:1] mux_tree_tapbuf_size3_1_sram ;
wire [0:1] mux_tree_tapbuf_size3_1_sram_inv ;
wire [0:1] mux_tree_tapbuf_size3_2_sram ;
wire [0:1] mux_tree_tapbuf_size3_2_sram_inv ;
wire [0:1] mux_tree_tapbuf_size3_3_sram ;
wire [0:1] mux_tree_tapbuf_size3_3_sram_inv ;
wire [0:1] mux_tree_tapbuf_size3_4_sram ;
wire [0:1] mux_tree_tapbuf_size3_4_sram_inv ;
wire [0:0] mux_tree_tapbuf_size3_mem_0_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size3_mem_1_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size3_mem_2_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size3_mem_3_ccff_tail ;
wire [0:2] mux_tree_tapbuf_size4_0_sram ;
wire [0:2] mux_tree_tapbuf_size4_0_sram_inv ;
wire [0:2] mux_tree_tapbuf_size4_1_sram ;
wire [0:2] mux_tree_tapbuf_size4_1_sram_inv ;
wire [0:2] mux_tree_tapbuf_size4_2_sram ;
wire [0:2] mux_tree_tapbuf_size4_2_sram_inv ;
wire [0:2] mux_tree_tapbuf_size4_3_sram ;
wire [0:2] mux_tree_tapbuf_size4_3_sram_inv ;
wire [0:2] mux_tree_tapbuf_size4_4_sram ;
wire [0:2] mux_tree_tapbuf_size4_4_sram_inv ;
wire [0:2] mux_tree_tapbuf_size4_5_sram ;
wire [0:2] mux_tree_tapbuf_size4_5_sram_inv ;
wire [0:2] mux_tree_tapbuf_size4_6_sram ;
wire [0:2] mux_tree_tapbuf_size4_6_sram_inv ;
wire [0:0] mux_tree_tapbuf_size4_mem_0_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size4_mem_1_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size4_mem_2_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size4_mem_3_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size4_mem_4_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size4_mem_5_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size4_mem_6_ccff_tail ;
wire [0:2] mux_tree_tapbuf_size5_0_sram ;
wire [0:2] mux_tree_tapbuf_size5_0_sram_inv ;
wire [0:2] mux_tree_tapbuf_size5_1_sram ;
wire [0:2] mux_tree_tapbuf_size5_1_sram_inv ;
wire [0:2] mux_tree_tapbuf_size5_2_sram ;
wire [0:2] mux_tree_tapbuf_size5_2_sram_inv ;
wire [0:2] mux_tree_tapbuf_size5_3_sram ;
wire [0:2] mux_tree_tapbuf_size5_3_sram_inv ;
wire [0:2] mux_tree_tapbuf_size5_4_sram ;
wire [0:2] mux_tree_tapbuf_size5_4_sram_inv ;
wire [0:0] mux_tree_tapbuf_size5_mem_0_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size5_mem_1_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size5_mem_2_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size5_mem_3_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size5_mem_4_ccff_tail ;
wire [0:2] mux_tree_tapbuf_size6_0_sram ;
wire [0:2] mux_tree_tapbuf_size6_0_sram_inv ;
wire [0:2] mux_tree_tapbuf_size6_1_sram ;
wire [0:2] mux_tree_tapbuf_size6_1_sram_inv ;
wire [0:2] mux_tree_tapbuf_size6_2_sram ;
wire [0:2] mux_tree_tapbuf_size6_2_sram_inv ;
wire [0:2] mux_tree_tapbuf_size6_3_sram ;
wire [0:2] mux_tree_tapbuf_size6_3_sram_inv ;
wire [0:2] mux_tree_tapbuf_size6_4_sram ;
wire [0:2] mux_tree_tapbuf_size6_4_sram_inv ;
wire [0:2] mux_tree_tapbuf_size6_5_sram ;
wire [0:2] mux_tree_tapbuf_size6_5_sram_inv ;
wire [0:2] mux_tree_tapbuf_size6_6_sram ;
wire [0:2] mux_tree_tapbuf_size6_6_sram_inv ;
wire [0:0] mux_tree_tapbuf_size6_mem_0_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size6_mem_1_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size6_mem_2_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size6_mem_3_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size6_mem_4_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size6_mem_5_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size6_mem_6_ccff_tail ;
wire [0:2] mux_tree_tapbuf_size7_0_sram ;
wire [0:2] mux_tree_tapbuf_size7_0_sram_inv ;
wire [0:2] mux_tree_tapbuf_size7_1_sram ;
wire [0:2] mux_tree_tapbuf_size7_1_sram_inv ;
wire [0:2] mux_tree_tapbuf_size7_2_sram ;
wire [0:2] mux_tree_tapbuf_size7_2_sram_inv ;
wire [0:0] mux_tree_tapbuf_size7_mem_0_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size7_mem_1_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size7_mem_2_ccff_tail ;

mux_tree_tapbuf_size6_4 mux_top_track_0 (
    .in ( { top_left_grid_pin_1_[0] , chanx_right_in[1] , chanx_right_in[8] , 
        chanx_right_in[15] , chany_bottom_in[2] , chany_bottom_in[12] } ) ,
    .sram ( mux_tree_tapbuf_size6_0_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size6_0_sram_inv ) , 
    .out ( chany_top_out[0] ) , .p0 ( optlc_net_122 ) ) ;
mux_tree_tapbuf_size6_5 mux_top_track_4 (
    .in ( { top_left_grid_pin_1_[0] , chanx_right_in[3] , chanx_right_in[10] , 
        chanx_right_in[17] , chany_bottom_in[5] , chany_bottom_in[14] } ) ,
    .sram ( mux_tree_tapbuf_size6_1_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size6_1_sram_inv ) , 
    .out ( chany_top_out[2] ) , .p0 ( optlc_net_122 ) ) ;
mux_tree_tapbuf_size6_1 mux_top_track_8 (
    .in ( { top_left_grid_pin_1_[0] , chanx_right_in[4] , chanx_right_in[11] , 
        chanx_right_in[18] , chany_bottom_in[6] , chany_bottom_in[16] } ) ,
    .sram ( mux_tree_tapbuf_size6_2_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size6_2_sram_inv ) , 
    .out ( chany_top_out[4] ) , .p0 ( optlc_net_123 ) ) ;
mux_tree_tapbuf_size6_3 mux_right_track_0 (
    .in ( { chany_top_in[2] , right_top_grid_pin_42_[0] , 
        right_top_grid_pin_44_[0] , right_top_grid_pin_46_[0] , 
        right_top_grid_pin_48_[0] , chany_bottom_in[2] } ) ,
    .sram ( mux_tree_tapbuf_size6_3_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size6_3_sram_inv ) , 
    .out ( chanx_right_out[0] ) , .p0 ( optlc_net_122 ) ) ;
mux_tree_tapbuf_size6_0_1 mux_bottom_track_1 (
    .in ( { chany_top_in[2] , chany_top_in[12] , chanx_right_in[5] , 
        chanx_right_in[12] , chanx_right_in[19] , bottom_left_grid_pin_1_[0] } ) ,
    .sram ( mux_tree_tapbuf_size6_4_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size6_4_sram_inv ) , 
    .out ( chany_bottom_out[0] ) , .p0 ( optlc_net_123 ) ) ;
mux_tree_tapbuf_size6_1 mux_bottom_track_5 (
    .in ( { chany_top_in[5] , chany_top_in[14] , chanx_right_in[3] , 
        chanx_right_in[10] , chanx_right_in[17] , bottom_left_grid_pin_1_[0] } ) ,
    .sram ( mux_tree_tapbuf_size6_5_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size6_5_sram_inv ) , 
    .out ( chany_bottom_out[2] ) , .p0 ( optlc_net_121 ) ) ;
mux_tree_tapbuf_size6_2 mux_bottom_track_9 (
    .in ( { chany_top_in[6] , chany_top_in[16] , chanx_right_in[2] , 
        chanx_right_in[9] , chanx_right_in[16] , bottom_left_grid_pin_1_[0] } ) ,
    .sram ( mux_tree_tapbuf_size6_6_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size6_6_sram_inv ) , 
    .out ( chany_bottom_out[4] ) , .p0 ( optlc_net_121 ) ) ;
mux_tree_tapbuf_size6_mem_4 mem_top_track_0 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( ccff_head ) , 
    .ccff_tail ( mux_tree_tapbuf_size6_mem_0_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size6_0_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size6_0_sram_inv ) ) ;
mux_tree_tapbuf_size6_mem_5 mem_top_track_4 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size5_mem_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size6_mem_1_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size6_1_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size6_1_sram_inv ) ) ;
mux_tree_tapbuf_size6_mem_1 mem_top_track_8 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size6_mem_1_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size6_mem_2_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size6_2_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size6_2_sram_inv ) ) ;
mux_tree_tapbuf_size6_mem_3 mem_right_track_0 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size4_mem_1_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size6_mem_3_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size6_3_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size6_3_sram_inv ) ) ;
mux_tree_tapbuf_size6_mem_0_1 mem_bottom_track_1 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size6_mem_4_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size6_4_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size6_4_sram_inv ) ) ;
mux_tree_tapbuf_size6_mem_1 mem_bottom_track_5 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size5_mem_2_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size6_mem_5_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size6_5_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size6_5_sram_inv ) ) ;
mux_tree_tapbuf_size6_mem_2 mem_bottom_track_9 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size6_mem_5_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size6_mem_6_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size6_6_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size6_6_sram_inv ) ) ;
mux_tree_tapbuf_size5_1 mux_top_track_2 (
    .in ( { chanx_right_in[2] , chanx_right_in[9] , chanx_right_in[16] , 
        chany_bottom_in[4] , chany_bottom_in[13] } ) ,
    .sram ( mux_tree_tapbuf_size5_0_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size5_0_sram_inv ) , 
    .out ( chany_top_out[1] ) , .p0 ( optlc_net_122 ) ) ;
mux_tree_tapbuf_size5_3 mux_top_track_16 (
    .in ( { chanx_right_in[5] , chanx_right_in[12] , chanx_right_in[19] , 
        chany_bottom_in[8] , chany_bottom_in[17] } ) ,
    .sram ( mux_tree_tapbuf_size5_1_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size5_1_sram_inv ) , 
    .out ( chany_top_out[8] ) , .p0 ( optlc_net_123 ) ) ;
mux_tree_tapbuf_size5_2 mux_bottom_track_3 (
    .in ( { chany_top_in[4] , chany_top_in[13] , chanx_right_in[4] , 
        chanx_right_in[11] , chanx_right_in[18] } ) ,
    .sram ( mux_tree_tapbuf_size5_2_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size5_2_sram_inv ) , 
    .out ( chany_bottom_out[1] ) , .p0 ( optlc_net_123 ) ) ;
mux_tree_tapbuf_size5_0_1 mux_bottom_track_17 (
    .in ( { chany_top_in[8] , chany_top_in[17] , chanx_right_in[1] , 
        chanx_right_in[8] , chanx_right_in[15] } ) ,
    .sram ( mux_tree_tapbuf_size5_3_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size5_3_sram_inv ) , 
    .out ( chany_bottom_out[8] ) , .p0 ( optlc_net_122 ) ) ;
mux_tree_tapbuf_size5_1 mux_bottom_track_25 (
    .in ( { chany_top_in[9] , chany_top_in[18] , chanx_right_in[0] , 
        chanx_right_in[7] , chanx_right_in[14] } ) ,
    .sram ( mux_tree_tapbuf_size5_4_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size5_4_sram_inv ) , 
    .out ( chany_bottom_out[12] ) , .p0 ( optlc_net_122 ) ) ;
mux_tree_tapbuf_size5_mem_1 mem_top_track_2 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size6_mem_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size5_mem_0_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size5_0_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size5_0_sram_inv ) ) ;
mux_tree_tapbuf_size5_mem_3 mem_top_track_16 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size6_mem_2_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size5_mem_1_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size5_1_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size5_1_sram_inv ) ) ;
mux_tree_tapbuf_size5_mem_2 mem_bottom_track_3 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size6_mem_4_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size5_mem_2_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size5_2_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size5_2_sram_inv ) ) ;
mux_tree_tapbuf_size5_mem_0_1 mem_bottom_track_17 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size6_mem_6_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size5_mem_3_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size5_3_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size5_3_sram_inv ) ) ;
mux_tree_tapbuf_size5_mem_1 mem_bottom_track_25 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size5_mem_3_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size5_mem_4_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size5_4_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size5_4_sram_inv ) ) ;
mux_tree_tapbuf_size4_5 mux_top_track_24 (
    .in ( { chanx_right_in[6] , chanx_right_in[13] , chany_bottom_in[9] , 
        chany_bottom_in[18] } ) ,
    .sram ( mux_tree_tapbuf_size4_0_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size4_0_sram_inv ) , 
    .out ( chany_top_out[12] ) , .p0 ( optlc_net_124 ) ) ;
mux_tree_tapbuf_size4 mux_top_track_32 (
    .in ( { chanx_right_in[0] , chanx_right_in[7] , chanx_right_in[14] , 
        chany_bottom_in[10] } ) ,
    .sram ( mux_tree_tapbuf_size4_1_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size4_1_sram_inv ) , 
    .out ( chany_top_out[16] ) , .p0 ( optlc_net_122 ) ) ;
mux_tree_tapbuf_size4_4 mux_right_track_8 (
    .in ( { chany_top_in[7] , chany_top_in[8] , right_top_grid_pin_42_[0] , 
        chany_bottom_in[8] } ) ,
    .sram ( mux_tree_tapbuf_size4_2_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size4_2_sram_inv ) , 
    .out ( chanx_right_out[4] ) , .p0 ( optlc_net_124 ) ) ;
mux_tree_tapbuf_size4_0 mux_right_track_10 (
    .in ( { chany_top_in[9] , chany_top_in[11] , right_top_grid_pin_43_[0] , 
        chany_bottom_in[9] } ) ,
    .sram ( mux_tree_tapbuf_size4_3_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size4_3_sram_inv ) , 
    .out ( chanx_right_out[5] ) , .p0 ( optlc_net_124 ) ) ;
mux_tree_tapbuf_size4_1 mux_right_track_12 (
    .in ( { chany_top_in[10] , chany_top_in[15] , right_top_grid_pin_44_[0] , 
        chany_bottom_in[10] } ) ,
    .sram ( mux_tree_tapbuf_size4_4_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size4_4_sram_inv ) , 
    .out ( chanx_right_out[6] ) , .p0 ( optlc_net_124 ) ) ;
mux_tree_tapbuf_size4_2 mux_right_track_14 (
    .in ( { chany_top_in[12] , chany_top_in[19] , right_top_grid_pin_45_[0] , 
        chany_bottom_in[12] } ) ,
    .sram ( mux_tree_tapbuf_size4_5_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size4_5_sram_inv ) , 
    .out ( chanx_right_out[7] ) , .p0 ( optlc_net_122 ) ) ;
mux_tree_tapbuf_size4_3 mux_right_track_24 (
    .in ( { chany_top_in[18] , right_top_grid_pin_42_[0] , 
        chany_bottom_in[18] , chany_bottom_in[19] } ) ,
    .sram ( mux_tree_tapbuf_size4_6_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size4_6_sram_inv ) , 
    .out ( chanx_right_out[12] ) , .p0 ( optlc_net_123 ) ) ;
mux_tree_tapbuf_size4_mem_5 mem_top_track_24 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size5_mem_1_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size4_mem_0_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size4_0_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size4_0_sram_inv ) ) ;
mux_tree_tapbuf_size4_mem mem_top_track_32 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size4_mem_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size4_mem_1_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size4_1_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size4_1_sram_inv ) ) ;
mux_tree_tapbuf_size4_mem_4 mem_right_track_8 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size7_mem_2_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size4_mem_2_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size4_2_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size4_2_sram_inv ) ) ;
mux_tree_tapbuf_size4_mem_0 mem_right_track_10 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size4_mem_2_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size4_mem_3_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size4_3_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size4_3_sram_inv ) ) ;
mux_tree_tapbuf_size4_mem_1 mem_right_track_12 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size4_mem_3_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size4_mem_4_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size4_4_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size4_4_sram_inv ) ) ;
mux_tree_tapbuf_size4_mem_2 mem_right_track_14 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size4_mem_4_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size4_mem_5_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size4_5_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size4_5_sram_inv ) ) ;
mux_tree_tapbuf_size4_mem_3 mem_right_track_24 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size3_mem_3_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size4_mem_6_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size4_6_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size4_6_sram_inv ) ) ;
mux_tree_tapbuf_size7_0 mux_right_track_2 (
    .in ( { chany_top_in[0] , chany_top_in[4] , right_top_grid_pin_43_[0] , 
        right_top_grid_pin_45_[0] , right_top_grid_pin_47_[0] , 
        right_top_grid_pin_49_[0] , chany_bottom_in[4] } ) ,
    .sram ( mux_tree_tapbuf_size7_0_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size7_0_sram_inv ) , 
    .out ( chanx_right_out[1] ) , .p0 ( optlc_net_122 ) ) ;
mux_tree_tapbuf_size7_1 mux_right_track_4 (
    .in ( { chany_top_in[1] , chany_top_in[5] , right_top_grid_pin_42_[0] , 
        right_top_grid_pin_44_[0] , right_top_grid_pin_46_[0] , 
        right_top_grid_pin_48_[0] , chany_bottom_in[5] } ) ,
    .sram ( mux_tree_tapbuf_size7_1_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size7_1_sram_inv ) , 
    .out ( chanx_right_out[2] ) , .p0 ( optlc_net_124 ) ) ;
mux_tree_tapbuf_size7 mux_right_track_6 (
    .in ( { chany_top_in[3] , chany_top_in[6] , right_top_grid_pin_43_[0] , 
        right_top_grid_pin_45_[0] , right_top_grid_pin_47_[0] , 
        right_top_grid_pin_49_[0] , chany_bottom_in[6] } ) ,
    .sram ( mux_tree_tapbuf_size7_2_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size7_2_sram_inv ) , 
    .out ( chanx_right_out[3] ) , .p0 ( optlc_net_124 ) ) ;
mux_tree_tapbuf_size7_mem_0 mem_right_track_2 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size6_mem_3_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size7_mem_0_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size7_0_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size7_0_sram_inv ) ) ;
mux_tree_tapbuf_size7_mem_1 mem_right_track_4 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size7_mem_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size7_mem_1_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size7_1_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size7_1_sram_inv ) ) ;
mux_tree_tapbuf_size7_mem mem_right_track_6 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size7_mem_1_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size7_mem_2_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size7_2_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size7_2_sram_inv ) ) ;
mux_tree_tapbuf_size3_1 mux_right_track_16 (
    .in ( { chany_top_in[13] , right_top_grid_pin_46_[0] , 
        chany_bottom_in[13] } ) ,
    .sram ( mux_tree_tapbuf_size3_0_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size3_0_sram_inv ) , 
    .out ( chanx_right_out[8] ) , .p0 ( optlc_net_122 ) ) ;
mux_tree_tapbuf_size3_2 mux_right_track_18 (
    .in ( { chany_top_in[14] , right_top_grid_pin_47_[0] , 
        chany_bottom_in[14] } ) ,
    .sram ( mux_tree_tapbuf_size3_1_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size3_1_sram_inv ) , 
    .out ( chanx_right_out[9] ) , .p0 ( optlc_net_122 ) ) ;
mux_tree_tapbuf_size3_3 mux_right_track_20 (
    .in ( { chany_top_in[16] , right_top_grid_pin_48_[0] , 
        chany_bottom_in[16] } ) ,
    .sram ( mux_tree_tapbuf_size3_2_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size3_2_sram_inv ) , 
    .out ( chanx_right_out[10] ) , .p0 ( optlc_net_124 ) ) ;
mux_tree_tapbuf_size3_4 mux_right_track_22 (
    .in ( { chany_top_in[17] , right_top_grid_pin_49_[0] , 
        chany_bottom_in[17] } ) ,
    .sram ( mux_tree_tapbuf_size3_3_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size3_3_sram_inv ) , 
    .out ( chanx_right_out[11] ) , .p0 ( optlc_net_124 ) ) ;
mux_tree_tapbuf_size3_0_1 mux_bottom_track_33 (
    .in ( { chany_top_in[10] , chanx_right_in[6] , chanx_right_in[13] } ) ,
    .sram ( mux_tree_tapbuf_size3_4_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size3_4_sram_inv ) , 
    .out ( chany_bottom_out[16] ) , .p0 ( optlc_net_123 ) ) ;
mux_tree_tapbuf_size3_mem_1 mem_right_track_16 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size4_mem_5_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size3_mem_0_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size3_0_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size3_0_sram_inv ) ) ;
mux_tree_tapbuf_size3_mem_2 mem_right_track_18 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size3_mem_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size3_mem_1_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size3_1_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size3_1_sram_inv ) ) ;
mux_tree_tapbuf_size3_mem_3 mem_right_track_20 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size3_mem_1_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size3_mem_2_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size3_2_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size3_2_sram_inv ) ) ;
mux_tree_tapbuf_size3_mem_4 mem_right_track_22 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size3_mem_2_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size3_mem_3_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size3_3_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size3_3_sram_inv ) ) ;
mux_tree_tapbuf_size3_mem_0_1 mem_bottom_track_33 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size5_mem_4_ccff_tail ) ,
    .ccff_tail ( { ropt_net_127 } ) ,
    .mem_out ( mux_tree_tapbuf_size3_4_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size3_4_sram_inv ) ) ;
mux_tree_tapbuf_size2_11 mux_right_track_26 (
    .in ( { right_top_grid_pin_43_[0] , chany_bottom_in[15] } ) ,
    .sram ( mux_tree_tapbuf_size2_0_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_0_sram_inv ) , 
    .out ( chanx_right_out[13] ) , .p0 ( optlc_net_123 ) ) ;
mux_tree_tapbuf_size2_mem_11 mem_right_track_26 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size4_mem_6_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_0_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_0_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_0_sram_inv ) ) ;
sky130_fd_sc_hd__conb_1 optlc_110 ( .LO ( SYNOPSYS_UNCONNECTED_1 ) , 
    .HI ( optlc_net_121 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_2__1 ( .A ( chany_top_in[4] ) , 
    .X ( ropt_net_142 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_3__2 ( .A ( chany_top_in[5] ) , 
    .X ( ropt_net_149 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_112 ( .LO ( SYNOPSYS_UNCONNECTED_2 ) , 
    .HI ( optlc_net_122 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_114 ( .LO ( SYNOPSYS_UNCONNECTED_3 ) , 
    .HI ( optlc_net_123 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_116 ( .LO ( SYNOPSYS_UNCONNECTED_4 ) , 
    .HI ( optlc_net_124 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_715 ( .A ( chany_bottom_in[9] ) , 
    .X ( ropt_net_153 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_8__7 ( .A ( chany_top_in[12] ) , 
    .X ( ropt_net_147 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_9__8 ( .A ( chany_top_in[13] ) , 
    .X ( ropt_net_133 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_716 ( 
    .A ( chany_bottom_in[16] ) , .X ( ropt_net_164 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_717 ( .A ( ropt_net_127 ) , 
    .X ( ropt_net_152 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_718 ( .A ( chany_bottom_in[0] ) , 
    .X ( ropt_net_163 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_719 ( .A ( ropt_net_129 ) , 
    .X ( ropt_net_154 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_720 ( .A ( chany_bottom_in[7] ) , 
    .X ( ropt_net_161 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_721 ( 
    .A ( chany_bottom_in[17] ) , .X ( chany_top_out[18] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_722 ( .A ( chany_top_in[16] ) , 
    .X ( chany_bottom_out[17] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_723 ( .A ( ropt_net_133 ) , 
    .X ( ropt_net_150 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_18__17 ( .A ( chany_bottom_in[4] ) , 
    .X ( ropt_net_144 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_19__18 ( .A ( chany_bottom_in[5] ) , 
    .X ( chany_top_out[6] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_724 ( .A ( ropt_net_134 ) , 
    .X ( ropt_net_151 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_725 ( .A ( ropt_net_135 ) , 
    .X ( ropt_net_155 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_726 ( .A ( chany_bottom_in[6] ) , 
    .X ( chany_top_out[7] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_727 ( .A ( chany_bottom_in[1] ) , 
    .X ( ropt_net_162 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_24__23 ( .A ( chany_bottom_in[10] ) , 
    .X ( ropt_net_145 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_728 ( .A ( ropt_net_138 ) , 
    .X ( ropt_net_158 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_26__25 ( .A ( chany_bottom_in[12] ) , 
    .X ( chany_top_out[13] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_729 ( .A ( ropt_net_139 ) , 
    .X ( chany_bottom_out[15] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_730 ( .A ( ropt_net_140 ) , 
    .X ( ropt_net_157 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_731 ( .A ( ropt_net_141 ) , 
    .X ( chany_bottom_out[11] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_732 ( .A ( ropt_net_142 ) , 
    .X ( chany_bottom_out[5] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_733 ( .A ( ropt_net_143 ) , 
    .X ( ropt_net_156 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_65 ( .A ( chany_top_in[6] ) , 
    .X ( ropt_net_148 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_66 ( .A ( chany_top_in[8] ) , 
    .X ( ropt_net_134 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_67 ( .A ( chany_top_in[9] ) , 
    .X ( ropt_net_129 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_741 ( .A ( ropt_net_150 ) , 
    .X ( chany_bottom_out[14] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_69 ( .A ( chany_top_in[17] ) , 
    .X ( BUF_net_69 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_743 ( .A ( ropt_net_151 ) , 
    .X ( chany_bottom_out[9] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_744 ( .A ( ropt_net_152 ) , 
    .X ( ccff_tail[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_72 ( .A ( chany_bottom_in[2] ) , 
    .X ( ropt_net_135 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_73 ( .A ( chany_bottom_in[3] ) , 
    .X ( ropt_net_138 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_745 ( .A ( ropt_net_153 ) , 
    .X ( chany_top_out[10] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_746 ( .A ( ropt_net_154 ) , 
    .X ( chany_bottom_out[10] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_747 ( .A ( ropt_net_155 ) , 
    .X ( chany_top_out[3] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_734 ( .A ( ropt_net_144 ) , 
    .X ( chany_top_out[5] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_78 ( .A ( chany_bottom_in[13] ) , 
    .X ( ropt_net_140 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_RR_79 ( .A ( chany_bottom_in[14] ) , 
    .X ( ropt_net_160 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_749 ( .A ( ropt_net_156 ) , 
    .X ( chanx_right_out[14] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_755 ( .A ( ropt_net_157 ) , 
    .X ( chany_top_out[14] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_RR_82 ( .A ( chany_bottom_in[18] ) , 
    .X ( chany_top_out[19] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_735 ( .A ( ropt_net_145 ) , 
    .X ( chany_top_out[11] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_736 ( .A ( ropt_net_146 ) , 
    .X ( chany_bottom_out[19] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_737 ( .A ( ropt_net_147 ) , 
    .X ( chany_bottom_out[13] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_738 ( .A ( ropt_net_148 ) , 
    .X ( ropt_net_159 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 BUFT_RR_87 ( .A ( BUF_net_69 ) , 
    .X ( chany_bottom_out[18] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_739 ( .A ( ropt_net_149 ) , 
    .X ( chany_bottom_out[6] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_P_96 ( .A ( chany_top_in[2] ) , 
    .X ( chany_bottom_out[3] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_P_97 ( .A ( chany_top_in[10] ) , 
    .X ( ropt_net_141 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_P_98 ( .A ( chany_top_in[14] ) , 
    .X ( ropt_net_139 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_P_99 ( .A ( chany_top_in[18] ) , 
    .X ( ropt_net_146 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_P_100 ( .A ( chany_bottom_in[8] ) , 
    .X ( chany_top_out[9] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_758 ( .A ( ropt_net_158 ) , 
    .X ( chanx_right_out[16] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_759 ( .A ( ropt_net_159 ) , 
    .X ( chany_bottom_out[7] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_762 ( .A ( ropt_net_160 ) , 
    .X ( chany_top_out[15] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_765 ( .A ( ropt_net_161 ) , 
    .X ( chanx_right_out[15] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_766 ( .A ( ropt_net_162 ) , 
    .X ( chanx_right_out[17] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_P_107 ( .A ( chany_bottom_in[11] ) , 
    .X ( ropt_net_143 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_767 ( .A ( ropt_net_163 ) , 
    .X ( chanx_right_out[18] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_768 ( .A ( ropt_net_164 ) , 
    .X ( chany_top_out[17] ) ) ;
endmodule


module mux_tree_tapbuf_size3_mem_0 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_18__39 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size3_mem ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_17__38 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_31 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size3_0 ( in , sram , sram_inv , out , p0 ) ;
input  [0:2] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;

const1_31 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( p0 ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
endmodule


module const1_16_1 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size3 ( in , sram , sram_inv , out , p0 ) ;
input  [0:2] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;

const1_16_1 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( p0 ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
endmodule


module mux_tree_tapbuf_size5_mem ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_16__37 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size5_mem_0 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_15__36 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_15_1 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size5 ( in , sram , sram_inv , out , p0 ) ;
input  [0:4] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;

const1_15_1 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , .A1 ( in[4] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
endmodule


module const1_14_1 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size5_0 ( in , sram , sram_inv , out , p0 ) ;
input  [0:4] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;

const1_14_1 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , .A1 ( in[4] ) , 
    .S ( sram[1] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
endmodule


module mux_tree_tapbuf_size6_mem ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_14__35 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size6_mem_0 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:2] mem_out ;
output [0:2] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_13__34 ( .A ( mem_out[2] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_13_1 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size6 ( in , sram , sram_inv , out , p0 ) ;
input  [0:5] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;

const1_13_1 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
endmodule


module const1_12_1 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size6_0 ( in , sram , sram_inv , out , p0 ) ;
input  [0:5] in ;
input  [0:2] sram ;
input  [0:2] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;

const1_12_1 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_7 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_12__33 ( .A ( mem_out[1] ) , 
    .X ( net_aps_33 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_71 ( .A ( net_aps_33 ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_6 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_11__32 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_5 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_10__31 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_4 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_9__30 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_3 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_8__29 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_2 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_7__28 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_1 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_6__27 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_0 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_5__26 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_9 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_4__25 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_3__24 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_10 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_2__23 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_tapbuf_size2_mem_8 ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_1__22 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_11_1 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_7 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_11_1 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
endmodule


module const1_10_1 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_6 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_10_1 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
endmodule


module const1_9_1 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_5 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_9_1 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
endmodule


module const1_8_1 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_4 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_8_1 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
endmodule


module const1_7_1 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_3 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_7_1 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
endmodule


module const1_6_1 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_2 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_6_1 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
endmodule


module const1_5_1 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_5_1 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
endmodule


module const1_4_1 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_0 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_4_1 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
endmodule


module const1_3_1 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_9 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_3_1 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_P_81 ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
endmodule


module const1_2_1 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;

const1_2_1 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_8 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , .X ( out[0] ) ) ;
endmodule


module const1_1_1 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_10 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_1_1 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
endmodule


module const1_0_1 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_tapbuf_size2_8 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;

const1_0_1 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__buf_4 sky130_fd_sc_hd__buf_4_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , .X ( out[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
endmodule


module sb_0__0_ ( prog_clk , chany_top_in , top_left_grid_pin_1_ , 
    chanx_right_in , right_top_grid_pin_42_ , right_top_grid_pin_43_ , 
    right_top_grid_pin_44_ , right_top_grid_pin_45_ , right_top_grid_pin_46_ , 
    right_top_grid_pin_47_ , right_top_grid_pin_48_ , right_top_grid_pin_49_ , 
    right_bottom_grid_pin_1_ , ccff_head , chany_top_out , chanx_right_out , 
    ccff_tail ) ;
input  [0:0] prog_clk ;
input  [0:19] chany_top_in ;
input  [0:0] top_left_grid_pin_1_ ;
input  [0:19] chanx_right_in ;
input  [0:0] right_top_grid_pin_42_ ;
input  [0:0] right_top_grid_pin_43_ ;
input  [0:0] right_top_grid_pin_44_ ;
input  [0:0] right_top_grid_pin_45_ ;
input  [0:0] right_top_grid_pin_46_ ;
input  [0:0] right_top_grid_pin_47_ ;
input  [0:0] right_top_grid_pin_48_ ;
input  [0:0] right_top_grid_pin_49_ ;
input  [0:0] right_bottom_grid_pin_1_ ;
input  [0:0] ccff_head ;
output [0:19] chany_top_out ;
output [0:19] chanx_right_out ;
output [0:0] ccff_tail ;

wire [0:1] mux_tree_tapbuf_size2_0_sram ;
wire [0:1] mux_tree_tapbuf_size2_0_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_10_sram ;
wire [0:1] mux_tree_tapbuf_size2_10_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_11_sram ;
wire [0:1] mux_tree_tapbuf_size2_11_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_1_sram ;
wire [0:1] mux_tree_tapbuf_size2_1_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_2_sram ;
wire [0:1] mux_tree_tapbuf_size2_2_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_3_sram ;
wire [0:1] mux_tree_tapbuf_size2_3_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_4_sram ;
wire [0:1] mux_tree_tapbuf_size2_4_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_5_sram ;
wire [0:1] mux_tree_tapbuf_size2_5_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_6_sram ;
wire [0:1] mux_tree_tapbuf_size2_6_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_7_sram ;
wire [0:1] mux_tree_tapbuf_size2_7_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_8_sram ;
wire [0:1] mux_tree_tapbuf_size2_8_sram_inv ;
wire [0:1] mux_tree_tapbuf_size2_9_sram ;
wire [0:1] mux_tree_tapbuf_size2_9_sram_inv ;
wire [0:0] mux_tree_tapbuf_size2_mem_0_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_10_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_1_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_2_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_3_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_4_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_5_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_6_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_7_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_8_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size2_mem_9_ccff_tail ;
wire [0:1] mux_tree_tapbuf_size3_0_sram ;
wire [0:1] mux_tree_tapbuf_size3_0_sram_inv ;
wire [0:1] mux_tree_tapbuf_size3_1_sram ;
wire [0:1] mux_tree_tapbuf_size3_1_sram_inv ;
wire [0:0] mux_tree_tapbuf_size3_mem_0_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size3_mem_1_ccff_tail ;
wire [0:2] mux_tree_tapbuf_size5_0_sram ;
wire [0:2] mux_tree_tapbuf_size5_0_sram_inv ;
wire [0:2] mux_tree_tapbuf_size5_1_sram ;
wire [0:2] mux_tree_tapbuf_size5_1_sram_inv ;
wire [0:0] mux_tree_tapbuf_size5_mem_0_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size5_mem_1_ccff_tail ;
wire [0:2] mux_tree_tapbuf_size6_0_sram ;
wire [0:2] mux_tree_tapbuf_size6_0_sram_inv ;
wire [0:2] mux_tree_tapbuf_size6_1_sram ;
wire [0:2] mux_tree_tapbuf_size6_1_sram_inv ;
wire [0:0] mux_tree_tapbuf_size6_mem_0_ccff_tail ;
wire [0:0] mux_tree_tapbuf_size6_mem_1_ccff_tail ;

mux_tree_tapbuf_size2_8 mux_top_track_0 (
    .in ( { top_left_grid_pin_1_[0] , chanx_right_in[1] } ) ,
    .sram ( mux_tree_tapbuf_size2_0_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_0_sram_inv ) , 
    .out ( chany_top_out[0] ) , .p0 ( optlc_net_99 ) ) ;
mux_tree_tapbuf_size2_10 mux_top_track_4 (
    .in ( { top_left_grid_pin_1_[0] , chanx_right_in[3] } ) ,
    .sram ( mux_tree_tapbuf_size2_1_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_1_sram_inv ) , 
    .out ( chany_top_out[2] ) , .p0 ( optlc_net_99 ) ) ;
mux_tree_tapbuf_size2 mux_top_track_8 (
    .in ( { top_left_grid_pin_1_[0] , chanx_right_in[5] } ) ,
    .sram ( mux_tree_tapbuf_size2_2_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_2_sram_inv ) , 
    .out ( chany_top_out[4] ) , .p0 ( optlc_net_100 ) ) ;
mux_tree_tapbuf_size2_9 mux_top_track_24 (
    .in ( { top_left_grid_pin_1_[0] , chanx_right_in[13] } ) ,
    .sram ( mux_tree_tapbuf_size2_3_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_3_sram_inv ) ,
    .out ( { ropt_net_107 } ) ,
    .p0 ( optlc_net_100 ) ) ;
mux_tree_tapbuf_size2_0 mux_right_track_10 (
    .in ( { chany_top_in[4] , right_top_grid_pin_43_[0] } ) ,
    .sram ( mux_tree_tapbuf_size2_4_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_4_sram_inv ) , 
    .out ( chanx_right_out[5] ) , .p0 ( optlc_net_100 ) ) ;
mux_tree_tapbuf_size2_1 mux_right_track_12 (
    .in ( { chany_top_in[5] , right_top_grid_pin_44_[0] } ) ,
    .sram ( mux_tree_tapbuf_size2_5_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_5_sram_inv ) , 
    .out ( chanx_right_out[6] ) , .p0 ( optlc_net_99 ) ) ;
mux_tree_tapbuf_size2_2 mux_right_track_14 (
    .in ( { chany_top_in[6] , right_top_grid_pin_45_[0] } ) ,
    .sram ( mux_tree_tapbuf_size2_6_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_6_sram_inv ) , 
    .out ( chanx_right_out[7] ) , .p0 ( optlc_net_99 ) ) ;
mux_tree_tapbuf_size2_3 mux_right_track_16 (
    .in ( { chany_top_in[7] , right_top_grid_pin_46_[0] } ) ,
    .sram ( mux_tree_tapbuf_size2_7_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_7_sram_inv ) , 
    .out ( chanx_right_out[8] ) , .p0 ( optlc_net_102 ) ) ;
mux_tree_tapbuf_size2_4 mux_right_track_18 (
    .in ( { chany_top_in[8] , right_top_grid_pin_47_[0] } ) ,
    .sram ( mux_tree_tapbuf_size2_8_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_8_sram_inv ) , 
    .out ( chanx_right_out[9] ) , .p0 ( optlc_net_102 ) ) ;
mux_tree_tapbuf_size2_5 mux_right_track_20 (
    .in ( { chany_top_in[9] , right_top_grid_pin_48_[0] } ) ,
    .sram ( mux_tree_tapbuf_size2_9_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_9_sram_inv ) , 
    .out ( chanx_right_out[10] ) , .p0 ( optlc_net_102 ) ) ;
mux_tree_tapbuf_size2_6 mux_right_track_22 (
    .in ( { chany_top_in[10] , right_top_grid_pin_49_[0] } ) ,
    .sram ( mux_tree_tapbuf_size2_10_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_10_sram_inv ) , 
    .out ( chanx_right_out[11] ) , .p0 ( optlc_net_101 ) ) ;
mux_tree_tapbuf_size2_7 mux_right_track_26 (
    .in ( { chany_top_in[12] , right_top_grid_pin_43_[0] } ) ,
    .sram ( mux_tree_tapbuf_size2_11_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size2_11_sram_inv ) , 
    .out ( chanx_right_out[13] ) , .p0 ( optlc_net_101 ) ) ;
mux_tree_tapbuf_size2_mem_8 mem_top_track_0 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( ccff_head ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_0_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_0_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_0_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem_10 mem_top_track_4 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_1_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_1_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_1_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem mem_top_track_8 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_1_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_2_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_2_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_2_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem_9 mem_top_track_24 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_2_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_3_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_3_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_3_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem_0 mem_right_track_10 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size3_mem_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_4_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_4_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_4_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem_1 mem_right_track_12 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_4_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_5_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_5_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_5_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem_2 mem_right_track_14 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_5_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_6_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_6_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_6_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem_3 mem_right_track_16 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_6_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_7_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_7_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_7_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem_4 mem_right_track_18 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_7_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_8_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_8_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_8_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem_5 mem_right_track_20 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_8_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_9_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_9_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_9_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem_6 mem_right_track_22 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_9_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size2_mem_10_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size2_10_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_10_sram_inv ) ) ;
mux_tree_tapbuf_size2_mem_7 mem_right_track_26 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size3_mem_1_ccff_tail ) ,
    .ccff_tail ( { ropt_net_105 } ) ,
    .mem_out ( mux_tree_tapbuf_size2_11_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size2_11_sram_inv ) ) ;
mux_tree_tapbuf_size6_0 mux_right_track_0 (
    .in ( { chany_top_in[19] , right_top_grid_pin_42_[0] , 
        right_top_grid_pin_44_[0] , right_top_grid_pin_46_[0] , 
        right_top_grid_pin_48_[0] , right_bottom_grid_pin_1_[0] } ) ,
    .sram ( mux_tree_tapbuf_size6_0_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size6_0_sram_inv ) , 
    .out ( chanx_right_out[0] ) , .p0 ( optlc_net_99 ) ) ;
mux_tree_tapbuf_size6 mux_right_track_4 (
    .in ( { chany_top_in[1] , right_top_grid_pin_42_[0] , 
        right_top_grid_pin_44_[0] , right_top_grid_pin_46_[0] , 
        right_top_grid_pin_48_[0] , right_bottom_grid_pin_1_[0] } ) ,
    .sram ( mux_tree_tapbuf_size6_1_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size6_1_sram_inv ) , 
    .out ( chanx_right_out[2] ) , .p0 ( optlc_net_102 ) ) ;
mux_tree_tapbuf_size6_mem_0 mem_right_track_0 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_3_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size6_mem_0_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size6_0_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size6_0_sram_inv ) ) ;
mux_tree_tapbuf_size6_mem mem_right_track_4 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size5_mem_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size6_mem_1_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size6_1_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size6_1_sram_inv ) ) ;
mux_tree_tapbuf_size5_0 mux_right_track_2 (
    .in ( { chany_top_in[0] , right_top_grid_pin_43_[0] , 
        right_top_grid_pin_45_[0] , right_top_grid_pin_47_[0] , 
        right_top_grid_pin_49_[0] } ) ,
    .sram ( mux_tree_tapbuf_size5_0_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size5_0_sram_inv ) , 
    .out ( chanx_right_out[1] ) , .p0 ( optlc_net_101 ) ) ;
mux_tree_tapbuf_size5 mux_right_track_6 (
    .in ( { chany_top_in[2] , right_top_grid_pin_43_[0] , 
        right_top_grid_pin_45_[0] , right_top_grid_pin_47_[0] , 
        right_top_grid_pin_49_[0] } ) ,
    .sram ( mux_tree_tapbuf_size5_1_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size5_1_sram_inv ) , 
    .out ( chanx_right_out[3] ) , .p0 ( optlc_net_101 ) ) ;
mux_tree_tapbuf_size5_mem_0 mem_right_track_2 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size6_mem_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size5_mem_0_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size5_0_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size5_0_sram_inv ) ) ;
mux_tree_tapbuf_size5_mem mem_right_track_6 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size6_mem_1_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size5_mem_1_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size5_1_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size5_1_sram_inv ) ) ;
mux_tree_tapbuf_size3 mux_right_track_8 (
    .in ( { chany_top_in[3] , right_top_grid_pin_42_[0] , 
        right_bottom_grid_pin_1_[0] } ) ,
    .sram ( mux_tree_tapbuf_size3_0_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size3_0_sram_inv ) , 
    .out ( chanx_right_out[4] ) , .p0 ( optlc_net_100 ) ) ;
mux_tree_tapbuf_size3_0 mux_right_track_24 (
    .in ( { chany_top_in[11] , right_top_grid_pin_42_[0] , 
        right_bottom_grid_pin_1_[0] } ) ,
    .sram ( mux_tree_tapbuf_size3_1_sram ) , 
    .sram_inv ( mux_tree_tapbuf_size3_1_sram_inv ) , 
    .out ( chanx_right_out[12] ) , .p0 ( optlc_net_100 ) ) ;
mux_tree_tapbuf_size3_mem mem_right_track_8 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size5_mem_1_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size3_mem_0_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size3_0_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size3_0_sram_inv ) ) ;
mux_tree_tapbuf_size3_mem_0 mem_right_track_24 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_tapbuf_size2_mem_10_ccff_tail ) , 
    .ccff_tail ( mux_tree_tapbuf_size3_mem_1_ccff_tail ) , 
    .mem_out ( mux_tree_tapbuf_size3_1_sram ) , 
    .mem_outb ( mux_tree_tapbuf_size3_1_sram_inv ) ) ;
sky130_fd_sc_hd__conb_1 optlc_93 ( .LO ( SYNOPSYS_UNCONNECTED_1 ) , 
    .HI ( optlc_net_99 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_95 ( .LO ( SYNOPSYS_UNCONNECTED_2 ) , 
    .HI ( optlc_net_100 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_97 ( .LO ( SYNOPSYS_UNCONNECTED_3 ) , 
    .HI ( optlc_net_101 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_99 ( .LO ( SYNOPSYS_UNCONNECTED_4 ) , 
    .HI ( optlc_net_102 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_688 ( .A ( ropt_net_104 ) , 
    .X ( chany_top_out[13] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_689 ( .A ( ropt_net_105 ) , 
    .X ( ropt_net_131 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_690 ( .A ( ropt_net_106 ) , 
    .X ( ropt_net_122 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_691 ( .A ( ropt_net_107 ) , 
    .X ( ropt_net_132 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_692 ( .A ( chanx_right_in[11] ) , 
    .X ( ropt_net_133 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_705 ( .A ( ropt_net_121 ) , 
    .X ( chany_top_out[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_11__10 ( .A ( chanx_right_in[7] ) , 
    .X ( aps_rename_2_ ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_693 ( .A ( ropt_net_109 ) , 
    .X ( ropt_net_128 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_694 ( .A ( chanx_right_in[2] ) , 
    .X ( ropt_net_121 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_695 ( .A ( ropt_net_111 ) , 
    .X ( ropt_net_124 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_696 ( .A ( chanx_right_in[16] ) , 
    .X ( chany_top_out[15] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_697 ( .A ( ropt_net_113 ) , 
    .X ( chanx_right_out[19] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_706 ( .A ( ropt_net_122 ) , 
    .X ( chany_top_out[19] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_698 ( .A ( ropt_net_114 ) , 
    .X ( ropt_net_126 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_707 ( .A ( ropt_net_123 ) , 
    .X ( chanx_right_out[17] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_20__19 ( .A ( chanx_right_in[17] ) , 
    .X ( ropt_net_111 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_21__20 ( .A ( chanx_right_in[18] ) , 
    .X ( ropt_net_120 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 FTB_22__21 ( .A ( chanx_right_in[19] ) , 
    .X ( chany_top_out[18] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_RR_44 ( .A ( chany_top_in[14] ) , 
    .X ( ropt_net_119 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_45 ( .A ( chany_top_in[16] ) , 
    .X ( ropt_net_116 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_RR_46 ( .A ( chany_top_in[17] ) , 
    .X ( ropt_net_115 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_RR_47 ( .A ( chany_top_in[18] ) , 
    .X ( ropt_net_113 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_708 ( .A ( ropt_net_124 ) , 
    .X ( chany_top_out[16] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_49 ( .A ( chanx_right_in[4] ) , 
    .X ( BUF_net_49 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_709 ( .A ( ropt_net_125 ) , 
    .X ( chany_top_out[17] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_699 ( .A ( ropt_net_115 ) , 
    .X ( chanx_right_out[18] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_700 ( .A ( ropt_net_116 ) , 
    .X ( ropt_net_123 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_701 ( .A ( ropt_net_117 ) , 
    .X ( ropt_net_129 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_702 ( .A ( ropt_net_118 ) , 
    .X ( chanx_right_out[16] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_710 ( .A ( ropt_net_126 ) , 
    .X ( chany_top_out[14] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_56 ( .A ( chanx_right_in[12] ) , 
    .X ( BUF_net_56 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_711 ( .A ( ropt_net_127 ) , 
    .X ( chany_top_out[3] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_58 ( .A ( chanx_right_in[15] ) , 
    .X ( ropt_net_114 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_703 ( .A ( ropt_net_119 ) , 
    .X ( chanx_right_out[15] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_704 ( .A ( ropt_net_120 ) , 
    .X ( ropt_net_125 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_63 ( .A ( chanx_right_in[6] ) , 
    .X ( ropt_net_109 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_712 ( .A ( ropt_net_128 ) , 
    .X ( chany_top_out[5] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_713 ( .A ( ropt_net_129 ) , 
    .X ( chanx_right_out[14] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_714 ( .A ( ropt_net_130 ) , 
    .X ( chany_top_out[8] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_715 ( .A ( ropt_net_131 ) , 
    .X ( ccff_tail[0] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_716 ( .A ( ropt_net_132 ) , 
    .X ( chany_top_out[12] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 BUFT_RR_69 ( .A ( chanx_right_in[14] ) , 
    .X ( ropt_net_104 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_717 ( .A ( ropt_net_133 ) , 
    .X ( chany_top_out[10] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_P_76 ( .A ( chany_top_in[13] ) , 
    .X ( ropt_net_117 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_P_77 ( .A ( chany_top_in[15] ) , 
    .X ( ropt_net_118 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 BUFT_P_80 ( .A ( aps_rename_2_ ) , 
    .X ( chany_top_out[6] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_P_82 ( .A ( chanx_right_in[0] ) , 
    .X ( ropt_net_106 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 BUFT_P_83 ( .A ( BUF_net_49 ) , 
    .X ( ropt_net_127 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_P_84 ( .A ( chanx_right_in[8] ) , 
    .X ( chany_top_out[7] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_P_85 ( .A ( chanx_right_in[9] ) , 
    .X ( ropt_net_130 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_P_86 ( .A ( chanx_right_in[10] ) , 
    .X ( chany_top_out[9] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 BUFT_P_88 ( .A ( BUF_net_56 ) , 
    .X ( chany_top_out[11] ) ) ;
endmodule


module direct_interc_4 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

assign out[0] = in[0] ;
endmodule


module GPIO_sky130_fd_sc_hd__dfxbp_1_mem_3 ( prog_clk , ccff_head , 
    ccff_tail , mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:0] mem_out ;
output [0:0] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( \_gOb0_mem_outb[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_2__2 ( .A ( mem_out[0] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module GPIO_3 ( A , IE , OE , Y , in , out , mem_out ) ;
output A ;
output IE ;
output OE ;
output Y ;
input  in ;
output out ;
input  mem_out ;

wire aps_rename_1_ ;

assign A = in ;
assign out = Y ;

sky130_fd_sc_hd__inv_1 ie_oe_inv ( .A ( IE ) , .Y ( OE ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_1__1 ( .A ( mem_out ) , 
    .X ( aps_rename_1_ ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 BUFT_RR_3 ( .A ( aps_rename_1_ ) , .X ( IE ) ) ;
endmodule


module logical_tile_io_mode_physical__iopad_3 ( prog_clk , gfpga_pad_GPIO_A , 
    gfpga_pad_GPIO_IE , gfpga_pad_GPIO_OE , gfpga_pad_GPIO_Y , iopad_outpad , 
    ccff_head , iopad_inpad , ccff_tail ) ;
input  [0:0] prog_clk ;
output [0:0] gfpga_pad_GPIO_A ;
output [0:0] gfpga_pad_GPIO_IE ;
output [0:0] gfpga_pad_GPIO_OE ;
inout  [0:0] gfpga_pad_GPIO_Y ;
input  [0:0] iopad_outpad ;
input  [0:0] ccff_head ;
output [0:0] iopad_inpad ;
output [0:0] ccff_tail ;

wire [0:0] GPIO_0_en ;

GPIO_3 GPIO_0_ ( .A ( gfpga_pad_GPIO_A[0] ) , .IE ( gfpga_pad_GPIO_IE[0] ) , 
    .OE ( gfpga_pad_GPIO_OE[0] ) , .Y ( gfpga_pad_GPIO_Y[0] ) , 
    .in ( iopad_outpad[0] ) , .out ( iopad_inpad[0] ) , 
    .mem_out ( GPIO_0_en[0] ) ) ;
GPIO_sky130_fd_sc_hd__dfxbp_1_mem_3 GPIO_sky130_fd_sc_hd__dfxbp_1_mem ( 
    .prog_clk ( prog_clk ) , .ccff_head ( ccff_head ) , 
    .ccff_tail ( ccff_tail ) , .mem_out ( GPIO_0_en ) ,
    .mem_outb ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
endmodule


module logical_tile_io_mode_io__3 ( prog_clk , gfpga_pad_GPIO_A , 
    gfpga_pad_GPIO_IE , gfpga_pad_GPIO_OE , gfpga_pad_GPIO_Y , io_outpad , 
    ccff_head , io_inpad , ccff_tail ) ;
input  [0:0] prog_clk ;
output [0:0] gfpga_pad_GPIO_A ;
output [0:0] gfpga_pad_GPIO_IE ;
output [0:0] gfpga_pad_GPIO_OE ;
inout  [0:0] gfpga_pad_GPIO_Y ;
input  [0:0] io_outpad ;
input  [0:0] ccff_head ;
output [0:0] io_inpad ;
output [0:0] ccff_tail ;

logical_tile_io_mode_physical__iopad_3 logical_tile_io_mode_physical__iopad_0 ( 
    .prog_clk ( prog_clk ) , .gfpga_pad_GPIO_A ( gfpga_pad_GPIO_A ) , 
    .gfpga_pad_GPIO_IE ( gfpga_pad_GPIO_IE ) , 
    .gfpga_pad_GPIO_OE ( gfpga_pad_GPIO_OE ) , 
    .gfpga_pad_GPIO_Y ( gfpga_pad_GPIO_Y ) , .iopad_outpad ( io_outpad ) , 
    .ccff_head ( ccff_head ) , .iopad_inpad ( io_inpad ) , 
    .ccff_tail ( ccff_tail ) ) ;
direct_interc_4 direct_interc_0_ (
    .in ( { SYNOPSYS_UNCONNECTED_1 } ) ,
    .out ( io_inpad ) ) ;
direct_interc_4 direct_interc_1_ (
    .in ( { SYNOPSYS_UNCONNECTED_2 } ) ,
    .out ( io_outpad ) ) ;
endmodule


module grid_io_left ( prog_clk , gfpga_pad_GPIO_A , gfpga_pad_GPIO_IE , 
    gfpga_pad_GPIO_OE , gfpga_pad_GPIO_Y , right_width_0_height_0__pin_0_ , 
    ccff_head , right_width_0_height_0__pin_1_upper , 
    right_width_0_height_0__pin_1_lower , ccff_tail ) ;
input  [0:0] prog_clk ;
output [0:0] gfpga_pad_GPIO_A ;
output [0:0] gfpga_pad_GPIO_IE ;
output [0:0] gfpga_pad_GPIO_OE ;
inout  [0:0] gfpga_pad_GPIO_Y ;
input  [0:0] right_width_0_height_0__pin_0_ ;
input  [0:0] ccff_head ;
output [0:0] right_width_0_height_0__pin_1_upper ;
output [0:0] right_width_0_height_0__pin_1_lower ;
output [0:0] ccff_tail ;

logical_tile_io_mode_io__3 logical_tile_io_mode_io__0 ( 
    .prog_clk ( prog_clk ) , .gfpga_pad_GPIO_A ( gfpga_pad_GPIO_A ) , 
    .gfpga_pad_GPIO_IE ( gfpga_pad_GPIO_IE ) , 
    .gfpga_pad_GPIO_OE ( gfpga_pad_GPIO_OE ) , 
    .gfpga_pad_GPIO_Y ( gfpga_pad_GPIO_Y ) , 
    .io_outpad ( right_width_0_height_0__pin_0_ ) , .ccff_head ( ccff_head ) , 
    .io_inpad ( right_width_0_height_0__pin_1_upper ) ,
    .ccff_tail ( { ropt_net_9 } ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_1__0 ( 
    .A ( right_width_0_height_0__pin_1_upper[0] ) , .X ( aps_rename_2_ ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 BUFT_RR_5 ( .A ( aps_rename_2_ ) , 
    .X ( right_width_0_height_0__pin_1_lower[0] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_569 ( .A ( ropt_net_9 ) , 
    .X ( ropt_net_11 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_570 ( .A ( ropt_net_11 ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module direct_interc_3 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

assign out[0] = in[0] ;
endmodule


module GPIO_sky130_fd_sc_hd__dfxbp_1_mem_2 ( prog_clk , ccff_head , 
    ccff_tail , mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:0] mem_out ;
output [0:0] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( \_gOb0_mem_outb[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_2__2 ( .A ( mem_out[0] ) , 
    .X ( net_net_8 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_RR_13 ( .A ( net_net_8 ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module GPIO_2 ( A , IE , OE , Y , in , out , mem_out ) ;
output A ;
output IE ;
output OE ;
output Y ;
input  in ;
output out ;
input  mem_out ;

wire aps_rename_1_ ;

assign A = in ;
assign out = Y ;

sky130_fd_sc_hd__inv_1 ie_oe_inv ( .A ( aps_rename_1_ ) , .Y ( OE ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_1__1 ( .A ( mem_out ) , 
    .X ( aps_rename_1_ ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_5 ( .A ( aps_rename_1_ ) , .X ( IE ) ) ;
endmodule


module logical_tile_io_mode_physical__iopad_2 ( prog_clk , gfpga_pad_GPIO_A , 
    gfpga_pad_GPIO_IE , gfpga_pad_GPIO_OE , gfpga_pad_GPIO_Y , iopad_outpad , 
    ccff_head , iopad_inpad , ccff_tail ) ;
input  [0:0] prog_clk ;
output [0:0] gfpga_pad_GPIO_A ;
output [0:0] gfpga_pad_GPIO_IE ;
output [0:0] gfpga_pad_GPIO_OE ;
inout  [0:0] gfpga_pad_GPIO_Y ;
input  [0:0] iopad_outpad ;
input  [0:0] ccff_head ;
output [0:0] iopad_inpad ;
output [0:0] ccff_tail ;

wire [0:0] GPIO_0_en ;

GPIO_2 GPIO_0_ ( .A ( gfpga_pad_GPIO_A[0] ) , .IE ( gfpga_pad_GPIO_IE[0] ) , 
    .OE ( gfpga_pad_GPIO_OE[0] ) , .Y ( gfpga_pad_GPIO_Y[0] ) , 
    .in ( iopad_outpad[0] ) , .out ( iopad_inpad[0] ) , 
    .mem_out ( GPIO_0_en[0] ) ) ;
GPIO_sky130_fd_sc_hd__dfxbp_1_mem_2 GPIO_sky130_fd_sc_hd__dfxbp_1_mem ( 
    .prog_clk ( prog_clk ) , .ccff_head ( ccff_head ) , 
    .ccff_tail ( ccff_tail ) , .mem_out ( GPIO_0_en ) ,
    .mem_outb ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
endmodule


module logical_tile_io_mode_io__2 ( prog_clk , gfpga_pad_GPIO_A , 
    gfpga_pad_GPIO_IE , gfpga_pad_GPIO_OE , gfpga_pad_GPIO_Y , io_outpad , 
    ccff_head , io_inpad , ccff_tail ) ;
input  [0:0] prog_clk ;
output [0:0] gfpga_pad_GPIO_A ;
output [0:0] gfpga_pad_GPIO_IE ;
output [0:0] gfpga_pad_GPIO_OE ;
inout  [0:0] gfpga_pad_GPIO_Y ;
input  [0:0] io_outpad ;
input  [0:0] ccff_head ;
output [0:0] io_inpad ;
output [0:0] ccff_tail ;

logical_tile_io_mode_physical__iopad_2 logical_tile_io_mode_physical__iopad_0 ( 
    .prog_clk ( prog_clk ) , .gfpga_pad_GPIO_A ( gfpga_pad_GPIO_A ) , 
    .gfpga_pad_GPIO_IE ( gfpga_pad_GPIO_IE ) , 
    .gfpga_pad_GPIO_OE ( gfpga_pad_GPIO_OE ) , 
    .gfpga_pad_GPIO_Y ( gfpga_pad_GPIO_Y ) , .iopad_outpad ( io_outpad ) , 
    .ccff_head ( ccff_head ) , .iopad_inpad ( io_inpad ) , 
    .ccff_tail ( ccff_tail ) ) ;
direct_interc_3 direct_interc_0_ (
    .in ( { SYNOPSYS_UNCONNECTED_1 } ) ,
    .out ( io_inpad ) ) ;
direct_interc_3 direct_interc_1_ (
    .in ( { SYNOPSYS_UNCONNECTED_2 } ) ,
    .out ( io_outpad ) ) ;
endmodule


module grid_io_bottom ( prog_clk , gfpga_pad_GPIO_A , gfpga_pad_GPIO_IE , 
    gfpga_pad_GPIO_OE , gfpga_pad_GPIO_Y , top_width_0_height_0__pin_0_ , 
    ccff_head , top_width_0_height_0__pin_1_upper , 
    top_width_0_height_0__pin_1_lower , ccff_tail ) ;
input  [0:0] prog_clk ;
output [0:0] gfpga_pad_GPIO_A ;
output [0:0] gfpga_pad_GPIO_IE ;
output [0:0] gfpga_pad_GPIO_OE ;
inout  [0:0] gfpga_pad_GPIO_Y ;
input  [0:0] top_width_0_height_0__pin_0_ ;
input  [0:0] ccff_head ;
output [0:0] top_width_0_height_0__pin_1_upper ;
output [0:0] top_width_0_height_0__pin_1_lower ;
output [0:0] ccff_tail ;

logical_tile_io_mode_io__2 logical_tile_io_mode_io__0 ( 
    .prog_clk ( prog_clk ) , .gfpga_pad_GPIO_A ( gfpga_pad_GPIO_A ) ,
    .gfpga_pad_GPIO_IE ( { ropt_net_16 } ) ,
    .gfpga_pad_GPIO_OE ( gfpga_pad_GPIO_OE ) , 
    .gfpga_pad_GPIO_Y ( gfpga_pad_GPIO_Y ) , 
    .io_outpad ( top_width_0_height_0__pin_0_ ) , .ccff_head ( ccff_head ) , 
    .io_inpad ( top_width_0_height_0__pin_1_upper ) ,
    .ccff_tail ( { ropt_net_17 } ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_1__0 ( 
    .A ( top_width_0_height_0__pin_1_upper[0] ) , .X ( aps_rename_2_ ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_6 ( .A ( aps_rename_2_ ) , 
    .X ( BUF_net_6 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_574 ( .A ( BUF_net_6 ) , 
    .X ( ropt_net_18 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_577 ( .A ( ropt_net_18 ) , 
    .X ( top_width_0_height_0__pin_1_lower[0] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_575 ( .A ( ropt_net_16 ) , 
    .X ( ropt_net_19 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_576 ( .A ( ropt_net_17 ) , 
    .X ( ccff_tail[0] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_578 ( .A ( ropt_net_19 ) , 
    .X ( gfpga_pad_GPIO_IE[0] ) ) ;
endmodule


module direct_interc_2 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

assign out[0] = in[0] ;
endmodule


module GPIO_sky130_fd_sc_hd__dfxbp_1_mem_1 ( prog_clk , ccff_head , 
    ccff_tail , mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:0] mem_out ;
output [0:0] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( \_gOb0_mem_outb[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_2__2 ( .A ( mem_out[0] ) , 
    .X ( net_net_7 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_RR_9 ( .A ( net_net_7 ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module GPIO_1 ( A , IE , OE , Y , in , out , mem_out ) ;
output A ;
output IE ;
output OE ;
output Y ;
input  in ;
output out ;
input  mem_out ;

assign A = in ;
assign out = Y ;

sky130_fd_sc_hd__inv_1 ie_oe_inv ( .A ( IE ) , .Y ( OE ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 FTB_1__1 ( .A ( mem_out ) , .X ( IE ) ) ;
endmodule


module logical_tile_io_mode_physical__iopad_1 ( prog_clk , gfpga_pad_GPIO_A , 
    gfpga_pad_GPIO_IE , gfpga_pad_GPIO_OE , gfpga_pad_GPIO_Y , iopad_outpad , 
    ccff_head , iopad_inpad , ccff_tail ) ;
input  [0:0] prog_clk ;
output [0:0] gfpga_pad_GPIO_A ;
output [0:0] gfpga_pad_GPIO_IE ;
output [0:0] gfpga_pad_GPIO_OE ;
inout  [0:0] gfpga_pad_GPIO_Y ;
input  [0:0] iopad_outpad ;
input  [0:0] ccff_head ;
output [0:0] iopad_inpad ;
output [0:0] ccff_tail ;

wire [0:0] GPIO_0_en ;

GPIO_1 GPIO_0_ ( .A ( gfpga_pad_GPIO_A[0] ) , .IE ( gfpga_pad_GPIO_IE[0] ) , 
    .OE ( gfpga_pad_GPIO_OE[0] ) , .Y ( gfpga_pad_GPIO_Y[0] ) , 
    .in ( iopad_outpad[0] ) , .out ( iopad_inpad[0] ) , 
    .mem_out ( GPIO_0_en[0] ) ) ;
GPIO_sky130_fd_sc_hd__dfxbp_1_mem_1 GPIO_sky130_fd_sc_hd__dfxbp_1_mem ( 
    .prog_clk ( prog_clk ) , .ccff_head ( ccff_head ) , 
    .ccff_tail ( ccff_tail ) , .mem_out ( GPIO_0_en ) ,
    .mem_outb ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
endmodule


module logical_tile_io_mode_io__1 ( prog_clk , gfpga_pad_GPIO_A , 
    gfpga_pad_GPIO_IE , gfpga_pad_GPIO_OE , gfpga_pad_GPIO_Y , io_outpad , 
    ccff_head , io_inpad , ccff_tail ) ;
input  [0:0] prog_clk ;
output [0:0] gfpga_pad_GPIO_A ;
output [0:0] gfpga_pad_GPIO_IE ;
output [0:0] gfpga_pad_GPIO_OE ;
inout  [0:0] gfpga_pad_GPIO_Y ;
input  [0:0] io_outpad ;
input  [0:0] ccff_head ;
output [0:0] io_inpad ;
output [0:0] ccff_tail ;

logical_tile_io_mode_physical__iopad_1 logical_tile_io_mode_physical__iopad_0 ( 
    .prog_clk ( prog_clk ) , .gfpga_pad_GPIO_A ( gfpga_pad_GPIO_A ) , 
    .gfpga_pad_GPIO_IE ( gfpga_pad_GPIO_IE ) , 
    .gfpga_pad_GPIO_OE ( gfpga_pad_GPIO_OE ) , 
    .gfpga_pad_GPIO_Y ( gfpga_pad_GPIO_Y ) , .iopad_outpad ( io_outpad ) , 
    .ccff_head ( ccff_head ) , .iopad_inpad ( io_inpad ) , 
    .ccff_tail ( ccff_tail ) ) ;
direct_interc_2 direct_interc_0_ (
    .in ( { SYNOPSYS_UNCONNECTED_1 } ) ,
    .out ( io_inpad ) ) ;
direct_interc_2 direct_interc_1_ (
    .in ( { SYNOPSYS_UNCONNECTED_2 } ) ,
    .out ( io_outpad ) ) ;
endmodule


module grid_io_right ( prog_clk , gfpga_pad_GPIO_A , gfpga_pad_GPIO_IE , 
    gfpga_pad_GPIO_OE , gfpga_pad_GPIO_Y , left_width_0_height_0__pin_0_ , 
    ccff_head , left_width_0_height_0__pin_1_upper , 
    left_width_0_height_0__pin_1_lower , ccff_tail ) ;
input  [0:0] prog_clk ;
output [0:0] gfpga_pad_GPIO_A ;
output [0:0] gfpga_pad_GPIO_IE ;
output [0:0] gfpga_pad_GPIO_OE ;
inout  [0:0] gfpga_pad_GPIO_Y ;
input  [0:0] left_width_0_height_0__pin_0_ ;
input  [0:0] ccff_head ;
output [0:0] left_width_0_height_0__pin_1_upper ;
output [0:0] left_width_0_height_0__pin_1_lower ;
output [0:0] ccff_tail ;

logical_tile_io_mode_io__1 logical_tile_io_mode_io__0 ( 
    .prog_clk ( prog_clk ) , .gfpga_pad_GPIO_A ( gfpga_pad_GPIO_A ) , 
    .gfpga_pad_GPIO_IE ( gfpga_pad_GPIO_IE ) , 
    .gfpga_pad_GPIO_OE ( gfpga_pad_GPIO_OE ) , 
    .gfpga_pad_GPIO_Y ( gfpga_pad_GPIO_Y ) , 
    .io_outpad ( left_width_0_height_0__pin_0_ ) , .ccff_head ( ccff_head ) , 
    .io_inpad ( left_width_0_height_0__pin_1_upper ) ,
    .ccff_tail ( { ropt_net_11 } ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_1__0 ( 
    .A ( left_width_0_height_0__pin_1_upper[0] ) , .X ( aps_rename_1_ ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_572 ( .A ( ropt_net_12 ) , 
    .X ( left_width_0_height_0__pin_1_lower[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_P_8 ( .A ( aps_rename_1_ ) , 
    .X ( ropt_net_10 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_570 ( .A ( ropt_net_10 ) , 
    .X ( ropt_net_12 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_571 ( .A ( ropt_net_11 ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module direct_interc_1 ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

assign out[0] = in[0] ;
endmodule


module GPIO_sky130_fd_sc_hd__dfxbp_1_mem ( prog_clk , ccff_head , ccff_tail , 
    mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:0] mem_out ;
output [0:0] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( \_gOb0_mem_outb[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_2__2 ( .A ( mem_out[0] ) , 
    .X ( net_net_7 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_13 ( .A ( net_net_7 ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module GPIO ( A , IE , OE , Y , in , out , mem_out ) ;
output A ;
output IE ;
output OE ;
output Y ;
input  in ;
output out ;
input  mem_out ;

wire aps_rename_1_ ;

assign A = in ;
assign out = Y ;

sky130_fd_sc_hd__inv_1 ie_oe_inv ( .A ( aps_rename_1_ ) , .Y ( OE ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_1__1 ( .A ( mem_out ) , 
    .X ( aps_rename_1_ ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 BUFT_P_12 ( .A ( aps_rename_1_ ) , .X ( IE ) ) ;
endmodule


module logical_tile_io_mode_physical__iopad ( prog_clk , gfpga_pad_GPIO_A , 
    gfpga_pad_GPIO_IE , gfpga_pad_GPIO_OE , gfpga_pad_GPIO_Y , iopad_outpad , 
    ccff_head , iopad_inpad , ccff_tail ) ;
input  [0:0] prog_clk ;
output [0:0] gfpga_pad_GPIO_A ;
output [0:0] gfpga_pad_GPIO_IE ;
output [0:0] gfpga_pad_GPIO_OE ;
inout  [0:0] gfpga_pad_GPIO_Y ;
input  [0:0] iopad_outpad ;
input  [0:0] ccff_head ;
output [0:0] iopad_inpad ;
output [0:0] ccff_tail ;

wire [0:0] GPIO_0_en ;

GPIO GPIO_0_ ( .A ( gfpga_pad_GPIO_A[0] ) , .IE ( gfpga_pad_GPIO_IE[0] ) , 
    .OE ( gfpga_pad_GPIO_OE[0] ) , .Y ( gfpga_pad_GPIO_Y[0] ) , 
    .in ( iopad_outpad[0] ) , .out ( iopad_inpad[0] ) , 
    .mem_out ( GPIO_0_en[0] ) ) ;
GPIO_sky130_fd_sc_hd__dfxbp_1_mem GPIO_sky130_fd_sc_hd__dfxbp_1_mem ( 
    .prog_clk ( prog_clk ) , .ccff_head ( ccff_head ) , 
    .ccff_tail ( ccff_tail ) , .mem_out ( GPIO_0_en ) ,
    .mem_outb ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
endmodule


module logical_tile_io_mode_io_ ( prog_clk , gfpga_pad_GPIO_A , 
    gfpga_pad_GPIO_IE , gfpga_pad_GPIO_OE , gfpga_pad_GPIO_Y , io_outpad , 
    ccff_head , io_inpad , ccff_tail ) ;
input  [0:0] prog_clk ;
output [0:0] gfpga_pad_GPIO_A ;
output [0:0] gfpga_pad_GPIO_IE ;
output [0:0] gfpga_pad_GPIO_OE ;
inout  [0:0] gfpga_pad_GPIO_Y ;
input  [0:0] io_outpad ;
input  [0:0] ccff_head ;
output [0:0] io_inpad ;
output [0:0] ccff_tail ;

logical_tile_io_mode_physical__iopad logical_tile_io_mode_physical__iopad_0 ( 
    .prog_clk ( prog_clk ) , .gfpga_pad_GPIO_A ( gfpga_pad_GPIO_A ) , 
    .gfpga_pad_GPIO_IE ( gfpga_pad_GPIO_IE ) , 
    .gfpga_pad_GPIO_OE ( gfpga_pad_GPIO_OE ) , 
    .gfpga_pad_GPIO_Y ( gfpga_pad_GPIO_Y ) , .iopad_outpad ( io_outpad ) , 
    .ccff_head ( ccff_head ) , .iopad_inpad ( io_inpad ) , 
    .ccff_tail ( ccff_tail ) ) ;
direct_interc_1 direct_interc_0_ (
    .in ( { SYNOPSYS_UNCONNECTED_1 } ) ,
    .out ( io_inpad ) ) ;
direct_interc_1 direct_interc_1_ (
    .in ( { SYNOPSYS_UNCONNECTED_2 } ) ,
    .out ( io_outpad ) ) ;
endmodule


module grid_io_top ( prog_clk , gfpga_pad_GPIO_A , gfpga_pad_GPIO_IE , 
    gfpga_pad_GPIO_OE , gfpga_pad_GPIO_Y , bottom_width_0_height_0__pin_0_ , 
    ccff_head , bottom_width_0_height_0__pin_1_upper , 
    bottom_width_0_height_0__pin_1_lower , ccff_tail ) ;
input  [0:0] prog_clk ;
output [0:0] gfpga_pad_GPIO_A ;
output [0:0] gfpga_pad_GPIO_IE ;
output [0:0] gfpga_pad_GPIO_OE ;
inout  [0:0] gfpga_pad_GPIO_Y ;
input  [0:0] bottom_width_0_height_0__pin_0_ ;
input  [0:0] ccff_head ;
output [0:0] bottom_width_0_height_0__pin_1_upper ;
output [0:0] bottom_width_0_height_0__pin_1_lower ;
output [0:0] ccff_tail ;

logical_tile_io_mode_io_ logical_tile_io_mode_io__0 ( .prog_clk ( prog_clk ) , 
    .gfpga_pad_GPIO_A ( gfpga_pad_GPIO_A ) ,
    .gfpga_pad_GPIO_IE ( { ropt_net_16 } ) ,
    .gfpga_pad_GPIO_OE ( gfpga_pad_GPIO_OE ) , 
    .gfpga_pad_GPIO_Y ( gfpga_pad_GPIO_Y ) , 
    .io_outpad ( bottom_width_0_height_0__pin_0_ ) , 
    .ccff_head ( ccff_head ) , 
    .io_inpad ( bottom_width_0_height_0__pin_1_upper ) ,
    .ccff_tail ( { ropt_net_15 } ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_1__0 ( 
    .A ( bottom_width_0_height_0__pin_1_upper[0] ) , .X ( aps_rename_2_ ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_5 ( .A ( aps_rename_2_ ) , 
    .X ( BUF_net_5 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_574 ( .A ( BUF_net_5 ) , 
    .X ( bottom_width_0_height_0__pin_1_lower[0] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_576 ( .A ( ropt_net_16 ) , 
    .X ( gfpga_pad_GPIO_IE[0] ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_575 ( .A ( ropt_net_15 ) , 
    .X ( ropt_net_17 ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_577 ( .A ( ropt_net_17 ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_size2_mem_23 ( prog_clk , ccff_head , ccff_tail , mem_out , 
    mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_40__55 ( .A ( mem_out[1] ) , 
    .X ( net_aps_55 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_109 ( .A ( net_aps_55 ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_size2_mem_22 ( prog_clk , ccff_head , ccff_tail , mem_out , 
    mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_39__54 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_size2_mem_21 ( prog_clk , ccff_head , ccff_tail , mem_out , 
    mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_38__53 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_size2_23 ( in , sram , sram_inv , out , p2 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p2 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;

const1 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p2 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , .X ( out[0] ) ) ;
endmodule


module const1_30 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_size2_22 ( in , sram , sram_inv , out , p2 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p2 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;

const1_30 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p2 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , .X ( out[0] ) ) ;
endmodule


module const1_29 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_size2_21 ( in , sram , sram_inv , out , p2 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p2 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;

const1_29 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p2 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , .X ( out[0] ) ) ;
endmodule


module logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff ( 
    Test_en , clk , ff_D , ff_DI , ff_Q , ff_clk , p_abuf2 ) ;
input  [0:0] Test_en ;
input  [0:0] clk ;
input  [0:0] ff_D ;
input  [0:0] ff_DI ;
output [0:0] ff_Q ;
input  [0:0] ff_clk ;
output p_abuf2 ;

sky130_fd_sc_hd__sdfxbp_1 sky130_fd_sc_hd__sdfxbp_1_0_ ( .D ( ff_D[0] ) , 
    .SCD ( ff_DI[0] ) , .SCE ( Test_en[0] ) , .CLK ( clk[0] ) , 
    .Q ( p_abuf2 ) , .Q_N ( SYNOPSYS_UNCONNECTED_1 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 BUFT_P_114 ( .A ( p_abuf2 ) , .X ( ff_Q[0] ) ) ;
endmodule


module logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_14 ( 
    Test_en , clk , ff_D , ff_DI , ff_Q , ff_clk ) ;
input  [0:0] Test_en ;
input  [0:0] clk ;
input  [0:0] ff_D ;
input  [0:0] ff_DI ;
output [0:0] ff_Q ;
input  [0:0] ff_clk ;

sky130_fd_sc_hd__sdfxbp_1 sky130_fd_sc_hd__sdfxbp_1_0_ ( .D ( ff_D[0] ) , 
    .SCD ( ff_DI[0] ) , .SCE ( Test_en[0] ) , .CLK ( clk[0] ) , 
    .Q ( ff_Q[0] ) , .Q_N ( SYNOPSYS_UNCONNECTED_1 ) ) ;
endmodule


module mux_tree_size2_mem ( prog_clk , ccff_head , ccff_tail , mem_out , 
    mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_37__52 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_28 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_size2 ( in , sram , sram_inv , out , p2 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p2 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;

const1_28 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p2 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , .X ( out[0] ) ) ;
endmodule


module frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem ( prog_clk , ccff_head , 
    ccff_tail , mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:16] mem_out ;
output [0:16] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_4_ ( .D ( mem_out[3] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[4] ) , .Q_N ( mem_outb[4] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_5_ ( .D ( mem_out[4] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[5] ) , .Q_N ( mem_outb[5] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_6_ ( .D ( mem_out[5] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[6] ) , .Q_N ( mem_outb[6] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_7_ ( .D ( mem_out[6] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[7] ) , .Q_N ( mem_outb[7] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_8_ ( .D ( mem_out[7] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[8] ) , .Q_N ( mem_outb[8] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_9_ ( .D ( mem_out[8] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[9] ) , .Q_N ( mem_outb[9] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_10_ ( .D ( mem_out[9] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[10] ) , .Q_N ( mem_outb[10] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_11_ ( .D ( mem_out[10] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[11] ) , .Q_N ( mem_outb[11] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_12_ ( .D ( mem_out[11] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[12] ) , .Q_N ( mem_outb[12] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_13_ ( .D ( mem_out[12] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[13] ) , .Q_N ( mem_outb[13] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_14_ ( .D ( mem_out[13] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[14] ) , .Q_N ( mem_outb[14] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_15_ ( .D ( mem_out[14] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[15] ) , .Q_N ( mem_outb[15] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_16_ ( .D ( mem_out[15] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[16] ) , .Q_N ( \_gOb7_mem_outb[16] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_36__51 ( .A ( mem_out[16] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module frac_lut4_mux ( in , sram , sram_inv , lut3_out , lut4_out ) ;
input  [0:15] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:1] lut3_out ;
output [0:0] lut4_out ;

wire [0:0] sky130_fd_sc_hd__buf_2_3_X ;
wire [0:0] sky130_fd_sc_hd__buf_2_4_X ;
wire [0:0] sky130_fd_sc_hd__buf_2_5_X ;
wire [0:0] sky130_fd_sc_hd__buf_2_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_10_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_11_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_12_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_13_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_14_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_12_X[0] ) , .X ( lut3_out[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_1_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_13_X[0] ) , .X ( lut3_out[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_2_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_14_X[0] ) , .X ( lut4_out[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_3_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .X ( sky130_fd_sc_hd__buf_2_3_X[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_4_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , 
    .X ( sky130_fd_sc_hd__buf_2_4_X[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_5_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_10_X[0] ) , 
    .X ( sky130_fd_sc_hd__buf_2_5_X[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_6_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_11_X[0] ) , 
    .X ( sky130_fd_sc_hd__buf_2_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_3_ ( .A0 ( in[7] ) , .A1 ( in[6] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_4_ ( .A0 ( in[9] ) , .A1 ( in[8] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_5_ ( .A0 ( in[11] ) , .A1 ( in[10] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_6_ ( .A0 ( in[13] ) , .A1 ( in[12] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_7_ ( .A0 ( in[15] ) , .A1 ( in[14] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_10_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_11_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( .A0 ( sky130_fd_sc_hd__buf_2_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__buf_2_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_12_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( .A0 ( sky130_fd_sc_hd__buf_2_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__buf_2_5_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_13_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_13_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_12_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_14_X[0] ) ) ;
endmodule


module frac_lut4 ( in , sram , sram_inv , mode , mode_inv , lut3_out , 
    lut4_out ) ;
input  [0:3] in ;
input  [0:15] sram ;
input  [0:15] sram_inv ;
input  [0:0] mode ;
input  [0:0] mode_inv ;
output [0:1] lut3_out ;
output [0:0] lut4_out ;

wire [0:0] sky130_fd_sc_hd__buf_2_0_X ;
wire [0:0] sky130_fd_sc_hd__buf_2_1_X ;
wire [0:0] sky130_fd_sc_hd__buf_2_2_X ;
wire [0:0] sky130_fd_sc_hd__buf_2_3_X ;
wire [0:0] sky130_fd_sc_hd__inv_1_0_Y ;
wire [0:0] sky130_fd_sc_hd__inv_1_1_Y ;
wire [0:0] sky130_fd_sc_hd__inv_1_2_Y ;
wire [0:0] sky130_fd_sc_hd__inv_1_3_Y ;
wire [0:0] sky130_fd_sc_hd__or2_1_0_X ;

sky130_fd_sc_hd__or2_0 sky130_fd_sc_hd__or2_1_0_ ( .A ( mode[0] ) , 
    .B ( in[3] ) , .X ( sky130_fd_sc_hd__or2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__inv_1 sky130_fd_sc_hd__inv_1_0_ ( .A ( in[0] ) , 
    .Y ( sky130_fd_sc_hd__inv_1_0_Y[0] ) ) ;
sky130_fd_sc_hd__inv_1 sky130_fd_sc_hd__inv_1_1_ ( .A ( in[1] ) , 
    .Y ( sky130_fd_sc_hd__inv_1_1_Y[0] ) ) ;
sky130_fd_sc_hd__inv_1 sky130_fd_sc_hd__inv_1_2_ ( .A ( in[2] ) , 
    .Y ( sky130_fd_sc_hd__inv_1_2_Y[0] ) ) ;
sky130_fd_sc_hd__inv_1 sky130_fd_sc_hd__inv_1_3_ ( 
    .A ( sky130_fd_sc_hd__or2_1_0_X[0] ) , 
    .Y ( sky130_fd_sc_hd__inv_1_3_Y[0] ) ) ;
sky130_fd_sc_hd__buf_2 sky130_fd_sc_hd__buf_2_0_ ( .A ( in[0] ) , 
    .X ( sky130_fd_sc_hd__buf_2_0_X[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_1_ ( .A ( in[1] ) , 
    .X ( sky130_fd_sc_hd__buf_2_1_X[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_2_ ( .A ( in[2] ) , 
    .X ( sky130_fd_sc_hd__buf_2_2_X[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_3_ ( 
    .A ( sky130_fd_sc_hd__or2_1_0_X[0] ) , 
    .X ( sky130_fd_sc_hd__buf_2_3_X[0] ) ) ;
frac_lut4_mux frac_lut4_mux_0_ ( .in ( sram ) ,
    .sram ( { sky130_fd_sc_hd__buf_2_0_X[0] , sky130_fd_sc_hd__buf_2_1_X[0] , 
        sky130_fd_sc_hd__buf_2_2_X[0] , sky130_fd_sc_hd__buf_2_3_X[0] } ) ,
    .sram_inv ( { sky130_fd_sc_hd__inv_1_0_Y[0] , 
        sky130_fd_sc_hd__inv_1_1_Y[0] , sky130_fd_sc_hd__inv_1_2_Y[0] , 
        sky130_fd_sc_hd__inv_1_3_Y[0] } ) ,
    .lut3_out ( lut3_out ) , .lut4_out ( lut4_out ) ) ;
endmodule


module logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4 ( 
    prog_clk , frac_lut4_in , ccff_head , frac_lut4_lut3_out , 
    frac_lut4_lut4_out , ccff_tail ) ;
input  [0:0] prog_clk ;
input  [0:3] frac_lut4_in ;
input  [0:0] ccff_head ;
output [0:1] frac_lut4_lut3_out ;
output [0:0] frac_lut4_lut4_out ;
output [0:0] ccff_tail ;

wire [0:0] frac_lut4_0_mode ;
wire [0:15] frac_lut4_0_sram ;
wire [0:15] frac_lut4_0_sram_inv ;

frac_lut4 frac_lut4_0_ ( .in ( frac_lut4_in ) , .sram ( frac_lut4_0_sram ) , 
    .sram_inv ( frac_lut4_0_sram_inv ) , .mode ( frac_lut4_0_mode ) ,
    .mode_inv ( { SYNOPSYS_UNCONNECTED_1 } ) ,
    .lut3_out ( frac_lut4_lut3_out ) , .lut4_out ( frac_lut4_lut4_out ) ) ;
frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem ( 
    .prog_clk ( prog_clk ) , .ccff_head ( ccff_head ) , 
    .ccff_tail ( ccff_tail ) ,
    .mem_out ( { frac_lut4_0_sram[0] , frac_lut4_0_sram[1] , 
        frac_lut4_0_sram[2] , frac_lut4_0_sram[3] , frac_lut4_0_sram[4] , 
        frac_lut4_0_sram[5] , frac_lut4_0_sram[6] , frac_lut4_0_sram[7] , 
        frac_lut4_0_sram[8] , frac_lut4_0_sram[9] , frac_lut4_0_sram[10] , 
        frac_lut4_0_sram[11] , frac_lut4_0_sram[12] , frac_lut4_0_sram[13] , 
        frac_lut4_0_sram[14] , frac_lut4_0_sram[15] , frac_lut4_0_mode[0] } ) ,
    .mem_outb ( { frac_lut4_0_sram_inv[0] , frac_lut4_0_sram_inv[1] , 
        frac_lut4_0_sram_inv[2] , frac_lut4_0_sram_inv[3] , 
        frac_lut4_0_sram_inv[4] , frac_lut4_0_sram_inv[5] , 
        frac_lut4_0_sram_inv[6] , frac_lut4_0_sram_inv[7] , 
        frac_lut4_0_sram_inv[8] , frac_lut4_0_sram_inv[9] , 
        frac_lut4_0_sram_inv[10] , frac_lut4_0_sram_inv[11] , 
        frac_lut4_0_sram_inv[12] , frac_lut4_0_sram_inv[13] , 
        frac_lut4_0_sram_inv[14] , frac_lut4_0_sram_inv[15] , 
        SYNOPSYS_UNCONNECTED_2 } ) ) ;
endmodule


module logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic ( 
    prog_clk , frac_logic_in , ccff_head , frac_logic_out , ccff_tail , p2 ) ;
input  [0:0] prog_clk ;
input  [0:3] frac_logic_in ;
input  [0:0] ccff_head ;
output [0:1] frac_logic_out ;
output [0:0] ccff_tail ;
input  p2 ;

wire [0:0] logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_ccff_tail ;
wire [0:0] logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_frac_lut4_lut3_out ;
wire [0:0] logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_frac_lut4_lut4_out ;
wire [0:1] mux_tree_size2_0_sram ;
wire [0:1] mux_tree_size2_0_sram_inv ;

logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4 logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0 ( 
    .prog_clk ( prog_clk ) , .frac_lut4_in ( frac_logic_in ) , 
    .ccff_head ( ccff_head ) ,
    .frac_lut4_lut3_out ( { 
        logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_frac_lut4_lut3_out[0] , 
        frac_logic_out[1] } ) ,
    
    .frac_lut4_lut4_out ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_frac_lut4_lut4_out ) , 
    .ccff_tail ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_ccff_tail ) ) ;
mux_tree_size2 mux_frac_logic_out_0 (
    .in ( { 
        logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_frac_lut4_lut4_out[0] , 
        logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_frac_lut4_lut3_out[0]
         } ) ,
    .sram ( mux_tree_size2_0_sram ) , 
    .sram_inv ( mux_tree_size2_0_sram_inv ) , .out ( frac_logic_out[0] ) , 
    .p2 ( p2 ) ) ;
mux_tree_size2_mem mem_frac_logic_out_0 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_ccff_tail ) , 
    .ccff_tail ( ccff_tail ) , .mem_out ( mux_tree_size2_0_sram ) , 
    .mem_outb ( mux_tree_size2_0_sram_inv ) ) ;
direct_interc direct_interc_0_ (
    .in ( { SYNOPSYS_UNCONNECTED_1 } ) ,
    .out ( frac_logic_out[1] ) ) ;
direct_interc direct_interc_1_ (
    .in ( { SYNOPSYS_UNCONNECTED_2 } ) ,
    .out ( frac_logic_in[0] ) ) ;
direct_interc direct_interc_2_ (
    .in ( { SYNOPSYS_UNCONNECTED_3 } ) ,
    .out ( frac_logic_in[1] ) ) ;
direct_interc direct_interc_3_ (
    .in ( { SYNOPSYS_UNCONNECTED_4 } ) ,
    .out ( frac_logic_in[2] ) ) ;
direct_interc direct_interc_4_ (
    .in ( { SYNOPSYS_UNCONNECTED_5 } ) ,
    .out ( frac_logic_in[3] ) ) ;
endmodule


module logical_tile_clb_mode_default__fle_mode_physical__fabric ( prog_clk , 
    Test_en , clk , fabric_in , fabric_regin , fabric_scin , fabric_clk , 
    ccff_head , fabric_out , fabric_regout , fabric_scout , ccff_tail , 
    p_abuf1 , p_abuf2 , p2 ) ;
input  [0:0] prog_clk ;
input  [0:0] Test_en ;
input  [0:0] clk ;
input  [0:3] fabric_in ;
input  [0:0] fabric_regin ;
input  [0:0] fabric_scin ;
input  [0:0] fabric_clk ;
input  [0:0] ccff_head ;
output [0:1] fabric_out ;
output [0:0] fabric_regout ;
output [0:0] fabric_scout ;
output [0:0] ccff_tail ;
output p_abuf1 ;
output p_abuf2 ;
input  p2 ;

wire [0:0] logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0_ff_Q ;
wire [0:0] logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_ccff_tail ;
wire [0:1] logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_frac_logic_out ;
wire [0:1] mux_tree_size2_0_sram ;
wire [0:1] mux_tree_size2_0_sram_inv ;
wire [0:1] mux_tree_size2_1_sram ;
wire [0:1] mux_tree_size2_1_sram_inv ;
wire [0:0] mux_tree_size2_2_out ;
wire [0:1] mux_tree_size2_2_sram ;
wire [0:1] mux_tree_size2_2_sram_inv ;
wire [0:0] mux_tree_size2_mem_0_ccff_tail ;
wire [0:0] mux_tree_size2_mem_1_ccff_tail ;

assign p_abuf1 = p_abuf2 ;

logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0 ( 
    .prog_clk ( prog_clk ) , .frac_logic_in ( fabric_in ) , 
    .ccff_head ( ccff_head ) , 
    .frac_logic_out ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_frac_logic_out ) , 
    .ccff_tail ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_ccff_tail ) , 
    .p2 ( p2 ) ) ;
logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_14 logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0 ( 
    .Test_en ( Test_en ) , .clk ( clk ) , .ff_D ( mux_tree_size2_2_out ) , 
    .ff_DI ( fabric_scin ) , 
    .ff_Q ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0_ff_Q ) ,
    .ff_clk ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1 ( 
    .Test_en ( Test_en ) , .clk ( clk ) , 
    .ff_D ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_frac_logic_out[1] ) , 
    .ff_DI ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0_ff_Q ) , 
    .ff_Q ( fabric_regout ) ,
    .ff_clk ( { SYNOPSYS_UNCONNECTED_2 } ) ,
    .p_abuf2 ( p_abuf2 ) ) ;
mux_tree_size2_21 mux_fabric_out_0 (
    .in ( { 
        logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0_ff_Q[0] , 
        logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_frac_logic_out[0]
         } ) ,
    .sram ( mux_tree_size2_0_sram ) , 
    .sram_inv ( mux_tree_size2_0_sram_inv ) , .out ( fabric_out[0] ) , 
    .p2 ( p2 ) ) ;
mux_tree_size2_22 mux_fabric_out_1 (
    .in ( { fabric_regout[0] , 
        logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_frac_logic_out[1]
         } ) ,
    .sram ( mux_tree_size2_1_sram ) , 
    .sram_inv ( mux_tree_size2_1_sram_inv ) , .out ( fabric_out[1] ) , 
    .p2 ( p2 ) ) ;
mux_tree_size2_23 mux_ff_0_D_0 (
    .in ( { 
        logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_frac_logic_out[0] , 
        fabric_regin[0] } ) ,
    .sram ( mux_tree_size2_2_sram ) , 
    .sram_inv ( mux_tree_size2_2_sram_inv ) , .out ( mux_tree_size2_2_out ) , 
    .p2 ( p2 ) ) ;
mux_tree_size2_mem_21 mem_fabric_out_0 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_size2_mem_0_ccff_tail ) , 
    .mem_out ( mux_tree_size2_0_sram ) , 
    .mem_outb ( mux_tree_size2_0_sram_inv ) ) ;
mux_tree_size2_mem_22 mem_fabric_out_1 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_size2_mem_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_size2_mem_1_ccff_tail ) , 
    .mem_out ( mux_tree_size2_1_sram ) , 
    .mem_outb ( mux_tree_size2_1_sram_inv ) ) ;
mux_tree_size2_mem_23 mem_ff_0_D_0 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_size2_mem_1_ccff_tail ) , .ccff_tail ( ccff_tail ) , 
    .mem_out ( mux_tree_size2_2_sram ) , 
    .mem_outb ( mux_tree_size2_2_sram_inv ) ) ;
direct_interc direct_interc_0_ (
    .in ( { SYNOPSYS_UNCONNECTED_3 } ) ,
    .out ( { p_abuf2 } ) ) ;
direct_interc direct_interc_1_ (
    .in ( { SYNOPSYS_UNCONNECTED_4 } ) ,
    .out ( { p_abuf2 } ) ) ;
direct_interc direct_interc_2_ (
    .in ( { SYNOPSYS_UNCONNECTED_5 } ) ,
    .out ( fabric_in[0] ) ) ;
direct_interc direct_interc_3_ (
    .in ( { SYNOPSYS_UNCONNECTED_6 } ) ,
    .out ( fabric_in[1] ) ) ;
direct_interc direct_interc_4_ (
    .in ( { SYNOPSYS_UNCONNECTED_7 } ) ,
    .out ( fabric_in[2] ) ) ;
direct_interc direct_interc_5_ (
    .in ( { SYNOPSYS_UNCONNECTED_8 } ) ,
    .out ( fabric_in[3] ) ) ;
direct_interc direct_interc_6_ (
    .in ( { SYNOPSYS_UNCONNECTED_9 } ) ,
    .out ( fabric_scin ) ) ;
direct_interc direct_interc_7_ (
    .in ( { SYNOPSYS_UNCONNECTED_10 } ) ,
    .out ( fabric_clk ) ) ;
direct_interc direct_interc_8_ (
    .in ( { SYNOPSYS_UNCONNECTED_11 } ) ,
    
    .out ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_frac_logic_out[1] ) ) ;
direct_interc direct_interc_9_ (
    .in ( { SYNOPSYS_UNCONNECTED_12 } ) ,
    
    .out ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0_ff_Q ) ) ;
direct_interc direct_interc_10_ (
    .in ( { SYNOPSYS_UNCONNECTED_13 } ) ,
    .out ( fabric_clk ) ) ;
sky130_fd_sc_hd__dlygate4sd1_1 FTB_1__256 ( .A ( fabric_regout[0] ) , 
    .X ( fabric_scout[0] ) ) ;
endmodule


module logical_tile_clb_mode_default__fle ( prog_clk , Test_en , clk , 
    fle_in , fle_regin , fle_scin , fle_clk , ccff_head , fle_out , 
    fle_regout , fle_scout , ccff_tail , p_abuf0 , p_abuf1 , p2 ) ;
input  [0:0] prog_clk ;
input  [0:0] Test_en ;
input  [0:0] clk ;
input  [0:3] fle_in ;
input  [0:0] fle_regin ;
input  [0:0] fle_scin ;
input  [0:0] fle_clk ;
input  [0:0] ccff_head ;
output [0:1] fle_out ;
output [0:0] fle_regout ;
output [0:0] fle_scout ;
output [0:0] ccff_tail ;
output p_abuf0 ;
output p_abuf1 ;
input  p2 ;

logical_tile_clb_mode_default__fle_mode_physical__fabric logical_tile_clb_mode_default__fle_mode_physical__fabric_0 ( 
    .prog_clk ( prog_clk ) , .Test_en ( Test_en ) , .clk ( clk ) , 
    .fabric_in ( fle_in ) , .fabric_regin ( fle_regin ) , 
    .fabric_scin ( fle_scin ) , .fabric_clk ( fle_clk ) , 
    .ccff_head ( ccff_head ) , .fabric_out ( fle_out ) , 
    .fabric_regout ( fle_regout ) , .fabric_scout ( fle_scout ) , 
    .ccff_tail ( ccff_tail ) , .p_abuf1 ( p_abuf0 ) , .p_abuf2 ( p_abuf1 ) , 
    .p2 ( p2 ) ) ;
direct_interc direct_interc_0_ (
    .in ( { SYNOPSYS_UNCONNECTED_1 } ) ,
    .out ( fle_out[0] ) ) ;
direct_interc direct_interc_1_ (
    .in ( { SYNOPSYS_UNCONNECTED_2 } ) ,
    .out ( fle_out[1] ) ) ;
direct_interc direct_interc_2_ (
    .in ( { SYNOPSYS_UNCONNECTED_3 } ) ,
    .out ( { p_abuf0 } ) ) ;
direct_interc direct_interc_3_ (
    .in ( { SYNOPSYS_UNCONNECTED_4 } ) ,
    .out ( { p_abuf1 } ) ) ;
direct_interc direct_interc_4_ (
    .in ( { SYNOPSYS_UNCONNECTED_5 } ) ,
    .out ( fle_in[0] ) ) ;
direct_interc direct_interc_5_ (
    .in ( { SYNOPSYS_UNCONNECTED_6 } ) ,
    .out ( fle_in[1] ) ) ;
direct_interc direct_interc_6_ (
    .in ( { SYNOPSYS_UNCONNECTED_7 } ) ,
    .out ( fle_in[2] ) ) ;
direct_interc direct_interc_7_ (
    .in ( { SYNOPSYS_UNCONNECTED_8 } ) ,
    .out ( fle_in[3] ) ) ;
direct_interc direct_interc_8_ (
    .in ( { SYNOPSYS_UNCONNECTED_9 } ) ,
    .out ( fle_regin ) ) ;
direct_interc direct_interc_9_ (
    .in ( { SYNOPSYS_UNCONNECTED_10 } ) ,
    .out ( fle_scin ) ) ;
direct_interc direct_interc_10_ (
    .in ( { SYNOPSYS_UNCONNECTED_11 } ) ,
    .out ( fle_clk ) ) ;
endmodule


module mux_tree_size2_mem_20 ( prog_clk , ccff_head , ccff_tail , mem_out , 
    mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_35__50 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_size2_mem_19 ( prog_clk , ccff_head , ccff_tail , mem_out , 
    mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_34__49 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_size2_mem_18 ( prog_clk , ccff_head , ccff_tail , mem_out , 
    mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_33__48 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_27 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_size2_20 ( in , sram , sram_inv , out , p1 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p1 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;

const1_27 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p1 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , .X ( out[0] ) ) ;
endmodule


module const1_26 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_size2_19 ( in , sram , sram_inv , out , p1 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p1 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;

const1_26 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p1 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , .X ( out[0] ) ) ;
endmodule


module const1_25 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_size2_18 ( in , sram , sram_inv , out , p1 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p1 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;

const1_25 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p1 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , .X ( out[0] ) ) ;
endmodule


module logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_13 ( 
    Test_en , clk , ff_D , ff_DI , ff_Q , ff_clk ) ;
input  [0:0] Test_en ;
input  [0:0] clk ;
input  [0:0] ff_D ;
input  [0:0] ff_DI ;
output [0:0] ff_Q ;
input  [0:0] ff_clk ;

sky130_fd_sc_hd__sdfxbp_1 sky130_fd_sc_hd__sdfxbp_1_0_ ( .D ( ff_D[0] ) , 
    .SCD ( ff_DI[0] ) , .SCE ( Test_en[0] ) , .CLK ( clk[0] ) , 
    .Q ( ff_Q[0] ) , .Q_N ( SYNOPSYS_UNCONNECTED_1 ) ) ;
endmodule


module logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_12 ( 
    Test_en , clk , ff_D , ff_DI , ff_Q , ff_clk ) ;
input  [0:0] Test_en ;
input  [0:0] clk ;
input  [0:0] ff_D ;
input  [0:0] ff_DI ;
output [0:0] ff_Q ;
input  [0:0] ff_clk ;

sky130_fd_sc_hd__sdfxbp_1 sky130_fd_sc_hd__sdfxbp_1_0_ ( .D ( ff_D[0] ) , 
    .SCD ( ff_DI[0] ) , .SCE ( Test_en[0] ) , .CLK ( clk[0] ) , 
    .Q ( ff_Q[0] ) , .Q_N ( SYNOPSYS_UNCONNECTED_1 ) ) ;
endmodule


module mux_tree_size2_mem_30 ( prog_clk , ccff_head , ccff_tail , mem_out , 
    mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_32__47 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_24 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_size2_30 ( in , sram , sram_inv , out , p1 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p1 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;

const1_24 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p1 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , .X ( out[0] ) ) ;
endmodule


module frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem_6 ( prog_clk , ccff_head , 
    ccff_tail , mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:16] mem_out ;
output [0:16] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_4_ ( .D ( mem_out[3] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[4] ) , .Q_N ( mem_outb[4] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_5_ ( .D ( mem_out[4] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[5] ) , .Q_N ( mem_outb[5] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_6_ ( .D ( mem_out[5] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[6] ) , .Q_N ( mem_outb[6] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_7_ ( .D ( mem_out[6] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[7] ) , .Q_N ( mem_outb[7] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_8_ ( .D ( mem_out[7] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[8] ) , .Q_N ( mem_outb[8] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_9_ ( .D ( mem_out[8] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[9] ) , .Q_N ( mem_outb[9] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_10_ ( .D ( mem_out[9] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[10] ) , .Q_N ( mem_outb[10] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_11_ ( .D ( mem_out[10] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[11] ) , .Q_N ( mem_outb[11] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_12_ ( .D ( mem_out[11] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[12] ) , .Q_N ( mem_outb[12] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_13_ ( .D ( mem_out[12] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[13] ) , .Q_N ( mem_outb[13] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_14_ ( .D ( mem_out[13] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[14] ) , .Q_N ( mem_outb[14] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_15_ ( .D ( mem_out[14] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[15] ) , .Q_N ( mem_outb[15] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_16_ ( .D ( mem_out[15] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[16] ) , .Q_N ( \_gOb6_mem_outb[16] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_31__46 ( .A ( mem_out[16] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module frac_lut4_mux_6 ( in , sram , sram_inv , lut3_out , lut4_out ) ;
input  [0:15] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:1] lut3_out ;
output [0:0] lut4_out ;

wire [0:0] sky130_fd_sc_hd__buf_2_3_X ;
wire [0:0] sky130_fd_sc_hd__buf_2_4_X ;
wire [0:0] sky130_fd_sc_hd__buf_2_5_X ;
wire [0:0] sky130_fd_sc_hd__buf_2_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_10_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_11_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_12_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_13_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_14_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

sky130_fd_sc_hd__buf_2 sky130_fd_sc_hd__buf_2_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_12_X[0] ) , .X ( lut3_out[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_1_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_13_X[0] ) , .X ( lut3_out[1] ) ) ;
sky130_fd_sc_hd__buf_2 sky130_fd_sc_hd__buf_2_2_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_14_X[0] ) , .X ( lut4_out[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_3_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .X ( sky130_fd_sc_hd__buf_2_3_X[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_4_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , 
    .X ( sky130_fd_sc_hd__buf_2_4_X[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_5_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_10_X[0] ) , 
    .X ( sky130_fd_sc_hd__buf_2_5_X[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_6_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_11_X[0] ) , 
    .X ( sky130_fd_sc_hd__buf_2_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_3_ ( .A0 ( in[7] ) , .A1 ( in[6] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_4_ ( .A0 ( in[9] ) , .A1 ( in[8] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_5_ ( .A0 ( in[11] ) , .A1 ( in[10] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_6_ ( .A0 ( in[13] ) , .A1 ( in[12] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_7_ ( .A0 ( in[15] ) , .A1 ( in[14] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_10_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_11_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( .A0 ( sky130_fd_sc_hd__buf_2_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__buf_2_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_12_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( .A0 ( sky130_fd_sc_hd__buf_2_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__buf_2_5_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_13_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_13_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_12_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_14_X[0] ) ) ;
endmodule


module frac_lut4_6 ( in , sram , sram_inv , mode , mode_inv , lut3_out , 
    lut4_out ) ;
input  [0:3] in ;
input  [0:15] sram ;
input  [0:15] sram_inv ;
input  [0:0] mode ;
input  [0:0] mode_inv ;
output [0:1] lut3_out ;
output [0:0] lut4_out ;

wire [0:0] sky130_fd_sc_hd__buf_2_0_X ;
wire [0:0] sky130_fd_sc_hd__buf_2_1_X ;
wire [0:0] sky130_fd_sc_hd__buf_2_2_X ;
wire [0:0] sky130_fd_sc_hd__buf_2_3_X ;
wire [0:0] sky130_fd_sc_hd__inv_1_0_Y ;
wire [0:0] sky130_fd_sc_hd__inv_1_1_Y ;
wire [0:0] sky130_fd_sc_hd__inv_1_2_Y ;
wire [0:0] sky130_fd_sc_hd__inv_1_3_Y ;
wire [0:0] sky130_fd_sc_hd__or2_1_0_X ;

sky130_fd_sc_hd__or2_0 sky130_fd_sc_hd__or2_1_0_ ( .A ( mode[0] ) , 
    .B ( in[3] ) , .X ( sky130_fd_sc_hd__or2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__inv_1 sky130_fd_sc_hd__inv_1_0_ ( .A ( in[0] ) , 
    .Y ( sky130_fd_sc_hd__inv_1_0_Y[0] ) ) ;
sky130_fd_sc_hd__inv_1 sky130_fd_sc_hd__inv_1_1_ ( .A ( in[1] ) , 
    .Y ( sky130_fd_sc_hd__inv_1_1_Y[0] ) ) ;
sky130_fd_sc_hd__inv_1 sky130_fd_sc_hd__inv_1_2_ ( .A ( in[2] ) , 
    .Y ( sky130_fd_sc_hd__inv_1_2_Y[0] ) ) ;
sky130_fd_sc_hd__inv_1 sky130_fd_sc_hd__inv_1_3_ ( 
    .A ( sky130_fd_sc_hd__or2_1_0_X[0] ) , 
    .Y ( sky130_fd_sc_hd__inv_1_3_Y[0] ) ) ;
sky130_fd_sc_hd__buf_2 sky130_fd_sc_hd__buf_2_0_ ( .A ( in[0] ) , 
    .X ( sky130_fd_sc_hd__buf_2_0_X[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_1_ ( .A ( in[1] ) , 
    .X ( sky130_fd_sc_hd__buf_2_1_X[0] ) ) ;
sky130_fd_sc_hd__buf_2 sky130_fd_sc_hd__buf_2_2_ ( .A ( in[2] ) , 
    .X ( sky130_fd_sc_hd__buf_2_2_X[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_3_ ( 
    .A ( sky130_fd_sc_hd__or2_1_0_X[0] ) , 
    .X ( sky130_fd_sc_hd__buf_2_3_X[0] ) ) ;
frac_lut4_mux_6 frac_lut4_mux_0_ ( .in ( sram ) ,
    .sram ( { sky130_fd_sc_hd__buf_2_0_X[0] , sky130_fd_sc_hd__buf_2_1_X[0] , 
        sky130_fd_sc_hd__buf_2_2_X[0] , sky130_fd_sc_hd__buf_2_3_X[0] } ) ,
    .sram_inv ( { sky130_fd_sc_hd__inv_1_0_Y[0] , 
        sky130_fd_sc_hd__inv_1_1_Y[0] , sky130_fd_sc_hd__inv_1_2_Y[0] , 
        sky130_fd_sc_hd__inv_1_3_Y[0] } ) ,
    .lut3_out ( lut3_out ) , .lut4_out ( lut4_out ) ) ;
endmodule


module logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_6 ( 
    prog_clk , frac_lut4_in , ccff_head , frac_lut4_lut3_out , 
    frac_lut4_lut4_out , ccff_tail ) ;
input  [0:0] prog_clk ;
input  [0:3] frac_lut4_in ;
input  [0:0] ccff_head ;
output [0:1] frac_lut4_lut3_out ;
output [0:0] frac_lut4_lut4_out ;
output [0:0] ccff_tail ;

wire [0:0] frac_lut4_0_mode ;
wire [0:15] frac_lut4_0_sram ;
wire [0:15] frac_lut4_0_sram_inv ;

frac_lut4_6 frac_lut4_0_ ( .in ( frac_lut4_in ) , .sram ( frac_lut4_0_sram ) , 
    .sram_inv ( frac_lut4_0_sram_inv ) , .mode ( frac_lut4_0_mode ) ,
    .mode_inv ( { SYNOPSYS_UNCONNECTED_1 } ) ,
    .lut3_out ( frac_lut4_lut3_out ) , .lut4_out ( frac_lut4_lut4_out ) ) ;
frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem_6 frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem ( 
    .prog_clk ( prog_clk ) , .ccff_head ( ccff_head ) , 
    .ccff_tail ( ccff_tail ) ,
    .mem_out ( { frac_lut4_0_sram[0] , frac_lut4_0_sram[1] , 
        frac_lut4_0_sram[2] , frac_lut4_0_sram[3] , frac_lut4_0_sram[4] , 
        frac_lut4_0_sram[5] , frac_lut4_0_sram[6] , frac_lut4_0_sram[7] , 
        frac_lut4_0_sram[8] , frac_lut4_0_sram[9] , frac_lut4_0_sram[10] , 
        frac_lut4_0_sram[11] , frac_lut4_0_sram[12] , frac_lut4_0_sram[13] , 
        frac_lut4_0_sram[14] , frac_lut4_0_sram[15] , frac_lut4_0_mode[0] } ) ,
    .mem_outb ( { frac_lut4_0_sram_inv[0] , frac_lut4_0_sram_inv[1] , 
        frac_lut4_0_sram_inv[2] , frac_lut4_0_sram_inv[3] , 
        frac_lut4_0_sram_inv[4] , frac_lut4_0_sram_inv[5] , 
        frac_lut4_0_sram_inv[6] , frac_lut4_0_sram_inv[7] , 
        frac_lut4_0_sram_inv[8] , frac_lut4_0_sram_inv[9] , 
        frac_lut4_0_sram_inv[10] , frac_lut4_0_sram_inv[11] , 
        frac_lut4_0_sram_inv[12] , frac_lut4_0_sram_inv[13] , 
        frac_lut4_0_sram_inv[14] , frac_lut4_0_sram_inv[15] , 
        SYNOPSYS_UNCONNECTED_2 } ) ) ;
endmodule


module logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_6 ( 
    prog_clk , frac_logic_in , ccff_head , frac_logic_out , ccff_tail , p1 ) ;
input  [0:0] prog_clk ;
input  [0:3] frac_logic_in ;
input  [0:0] ccff_head ;
output [0:1] frac_logic_out ;
output [0:0] ccff_tail ;
input  p1 ;

wire [0:0] logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_ccff_tail ;
wire [0:0] logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_frac_lut4_lut3_out ;
wire [0:0] logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_frac_lut4_lut4_out ;
wire [0:1] mux_tree_size2_0_sram ;
wire [0:1] mux_tree_size2_0_sram_inv ;

logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_6 logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0 ( 
    .prog_clk ( prog_clk ) , .frac_lut4_in ( frac_logic_in ) , 
    .ccff_head ( ccff_head ) ,
    .frac_lut4_lut3_out ( { 
        logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_frac_lut4_lut3_out[0] , 
        frac_logic_out[1] } ) ,
    
    .frac_lut4_lut4_out ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_frac_lut4_lut4_out ) , 
    .ccff_tail ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_ccff_tail ) ) ;
mux_tree_size2_30 mux_frac_logic_out_0 (
    .in ( { 
        logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_frac_lut4_lut4_out[0] , 
        logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_frac_lut4_lut3_out[0]
         } ) ,
    .sram ( mux_tree_size2_0_sram ) , 
    .sram_inv ( mux_tree_size2_0_sram_inv ) , .out ( frac_logic_out[0] ) , 
    .p1 ( p1 ) ) ;
mux_tree_size2_mem_30 mem_frac_logic_out_0 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_ccff_tail ) , 
    .ccff_tail ( ccff_tail ) , .mem_out ( mux_tree_size2_0_sram ) , 
    .mem_outb ( mux_tree_size2_0_sram_inv ) ) ;
direct_interc direct_interc_0_ (
    .in ( { SYNOPSYS_UNCONNECTED_1 } ) ,
    .out ( frac_logic_out[1] ) ) ;
direct_interc direct_interc_1_ (
    .in ( { SYNOPSYS_UNCONNECTED_2 } ) ,
    .out ( frac_logic_in[0] ) ) ;
direct_interc direct_interc_2_ (
    .in ( { SYNOPSYS_UNCONNECTED_3 } ) ,
    .out ( frac_logic_in[1] ) ) ;
direct_interc direct_interc_3_ (
    .in ( { SYNOPSYS_UNCONNECTED_4 } ) ,
    .out ( frac_logic_in[2] ) ) ;
direct_interc direct_interc_4_ (
    .in ( { SYNOPSYS_UNCONNECTED_5 } ) ,
    .out ( frac_logic_in[3] ) ) ;
endmodule


module logical_tile_clb_mode_default__fle_mode_physical__fabric_6 ( prog_clk , 
    Test_en , clk , fabric_in , fabric_regin , fabric_scin , fabric_clk , 
    ccff_head , fabric_out , fabric_regout , fabric_scout , ccff_tail , p1 ) ;
input  [0:0] prog_clk ;
input  [0:0] Test_en ;
input  [0:0] clk ;
input  [0:3] fabric_in ;
input  [0:0] fabric_regin ;
input  [0:0] fabric_scin ;
input  [0:0] fabric_clk ;
input  [0:0] ccff_head ;
output [0:1] fabric_out ;
output [0:0] fabric_regout ;
output [0:0] fabric_scout ;
output [0:0] ccff_tail ;
input  p1 ;

wire [0:0] logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0_ff_Q ;
wire [0:0] logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_ccff_tail ;
wire [0:1] logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_frac_logic_out ;
wire [0:1] mux_tree_size2_0_sram ;
wire [0:1] mux_tree_size2_0_sram_inv ;
wire [0:1] mux_tree_size2_1_sram ;
wire [0:1] mux_tree_size2_1_sram_inv ;
wire [0:0] mux_tree_size2_2_out ;
wire [0:1] mux_tree_size2_2_sram ;
wire [0:1] mux_tree_size2_2_sram_inv ;
wire [0:0] mux_tree_size2_mem_0_ccff_tail ;
wire [0:0] mux_tree_size2_mem_1_ccff_tail ;

assign fabric_regout[0] = fabric_scout[0] ;

logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_6 logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0 ( 
    .prog_clk ( prog_clk ) , .frac_logic_in ( fabric_in ) , 
    .ccff_head ( ccff_head ) , 
    .frac_logic_out ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_frac_logic_out ) , 
    .ccff_tail ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_ccff_tail ) , 
    .p1 ( p1 ) ) ;
logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_12 logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0 ( 
    .Test_en ( Test_en ) , .clk ( clk ) , .ff_D ( mux_tree_size2_2_out ) , 
    .ff_DI ( fabric_scin ) , 
    .ff_Q ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0_ff_Q ) ,
    .ff_clk ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_13 logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1 ( 
    .Test_en ( Test_en ) , .clk ( clk ) , 
    .ff_D ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_frac_logic_out[1] ) , 
    .ff_DI ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0_ff_Q ) , 
    .ff_Q ( fabric_scout ) ,
    .ff_clk ( { SYNOPSYS_UNCONNECTED_2 } ) ) ;
mux_tree_size2_18 mux_fabric_out_0 (
    .in ( { 
        logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0_ff_Q[0] , 
        logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_frac_logic_out[0]
         } ) ,
    .sram ( mux_tree_size2_0_sram ) , 
    .sram_inv ( mux_tree_size2_0_sram_inv ) , .out ( fabric_out[0] ) , 
    .p1 ( p1 ) ) ;
mux_tree_size2_19 mux_fabric_out_1 (
    .in ( { fabric_scout[0] , 
        logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_frac_logic_out[1]
         } ) ,
    .sram ( mux_tree_size2_1_sram ) , 
    .sram_inv ( mux_tree_size2_1_sram_inv ) , .out ( fabric_out[1] ) , 
    .p1 ( p1 ) ) ;
mux_tree_size2_20 mux_ff_0_D_0 (
    .in ( { 
        logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_frac_logic_out[0] , 
        fabric_regin[0] } ) ,
    .sram ( mux_tree_size2_2_sram ) , 
    .sram_inv ( mux_tree_size2_2_sram_inv ) , .out ( mux_tree_size2_2_out ) , 
    .p1 ( p1 ) ) ;
mux_tree_size2_mem_18 mem_fabric_out_0 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_size2_mem_0_ccff_tail ) , 
    .mem_out ( mux_tree_size2_0_sram ) , 
    .mem_outb ( mux_tree_size2_0_sram_inv ) ) ;
mux_tree_size2_mem_19 mem_fabric_out_1 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_size2_mem_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_size2_mem_1_ccff_tail ) , 
    .mem_out ( mux_tree_size2_1_sram ) , 
    .mem_outb ( mux_tree_size2_1_sram_inv ) ) ;
mux_tree_size2_mem_20 mem_ff_0_D_0 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_size2_mem_1_ccff_tail ) , .ccff_tail ( ccff_tail ) , 
    .mem_out ( mux_tree_size2_2_sram ) , 
    .mem_outb ( mux_tree_size2_2_sram_inv ) ) ;
direct_interc direct_interc_0_ (
    .in ( { SYNOPSYS_UNCONNECTED_3 } ) ,
    .out ( fabric_scout ) ) ;
direct_interc direct_interc_1_ (
    .in ( { SYNOPSYS_UNCONNECTED_4 } ) ,
    .out ( fabric_scout ) ) ;
direct_interc direct_interc_2_ (
    .in ( { SYNOPSYS_UNCONNECTED_5 } ) ,
    .out ( fabric_in[0] ) ) ;
direct_interc direct_interc_3_ (
    .in ( { SYNOPSYS_UNCONNECTED_6 } ) ,
    .out ( fabric_in[1] ) ) ;
direct_interc direct_interc_4_ (
    .in ( { SYNOPSYS_UNCONNECTED_7 } ) ,
    .out ( fabric_in[2] ) ) ;
direct_interc direct_interc_5_ (
    .in ( { SYNOPSYS_UNCONNECTED_8 } ) ,
    .out ( fabric_in[3] ) ) ;
direct_interc direct_interc_6_ (
    .in ( { SYNOPSYS_UNCONNECTED_9 } ) ,
    .out ( fabric_scin ) ) ;
direct_interc direct_interc_7_ (
    .in ( { SYNOPSYS_UNCONNECTED_10 } ) ,
    .out ( fabric_clk ) ) ;
direct_interc direct_interc_8_ (
    .in ( { SYNOPSYS_UNCONNECTED_11 } ) ,
    
    .out ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_frac_logic_out[1] ) ) ;
direct_interc direct_interc_9_ (
    .in ( { SYNOPSYS_UNCONNECTED_12 } ) ,
    
    .out ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0_ff_Q ) ) ;
direct_interc direct_interc_10_ (
    .in ( { SYNOPSYS_UNCONNECTED_13 } ) ,
    .out ( fabric_clk ) ) ;
endmodule


module logical_tile_clb_mode_default__fle_6 ( prog_clk , Test_en , clk , 
    fle_in , fle_regin , fle_scin , fle_clk , ccff_head , fle_out , 
    fle_regout , fle_scout , ccff_tail , p1 ) ;
input  [0:0] prog_clk ;
input  [0:0] Test_en ;
input  [0:0] clk ;
input  [0:3] fle_in ;
input  [0:0] fle_regin ;
input  [0:0] fle_scin ;
input  [0:0] fle_clk ;
input  [0:0] ccff_head ;
output [0:1] fle_out ;
output [0:0] fle_regout ;
output [0:0] fle_scout ;
output [0:0] ccff_tail ;
input  p1 ;

logical_tile_clb_mode_default__fle_mode_physical__fabric_6 logical_tile_clb_mode_default__fle_mode_physical__fabric_0 ( 
    .prog_clk ( prog_clk ) , .Test_en ( Test_en ) , .clk ( clk ) , 
    .fabric_in ( fle_in ) , .fabric_regin ( fle_regin ) , 
    .fabric_scin ( fle_scin ) , .fabric_clk ( fle_clk ) , 
    .ccff_head ( ccff_head ) , .fabric_out ( fle_out ) , 
    .fabric_regout ( fle_regout ) , .fabric_scout ( fle_scout ) , 
    .ccff_tail ( ccff_tail ) , .p1 ( p1 ) ) ;
direct_interc direct_interc_0_ (
    .in ( { SYNOPSYS_UNCONNECTED_1 } ) ,
    .out ( fle_out[0] ) ) ;
direct_interc direct_interc_1_ (
    .in ( { SYNOPSYS_UNCONNECTED_2 } ) ,
    .out ( fle_out[1] ) ) ;
direct_interc direct_interc_2_ (
    .in ( { SYNOPSYS_UNCONNECTED_3 } ) ,
    .out ( fle_regout ) ) ;
direct_interc direct_interc_3_ (
    .in ( { SYNOPSYS_UNCONNECTED_4 } ) ,
    .out ( fle_scout ) ) ;
direct_interc direct_interc_4_ (
    .in ( { SYNOPSYS_UNCONNECTED_5 } ) ,
    .out ( fle_in[0] ) ) ;
direct_interc direct_interc_5_ (
    .in ( { SYNOPSYS_UNCONNECTED_6 } ) ,
    .out ( fle_in[1] ) ) ;
direct_interc direct_interc_6_ (
    .in ( { SYNOPSYS_UNCONNECTED_7 } ) ,
    .out ( fle_in[2] ) ) ;
direct_interc direct_interc_7_ (
    .in ( { SYNOPSYS_UNCONNECTED_8 } ) ,
    .out ( fle_in[3] ) ) ;
direct_interc direct_interc_8_ (
    .in ( { SYNOPSYS_UNCONNECTED_9 } ) ,
    .out ( fle_regin ) ) ;
direct_interc direct_interc_9_ (
    .in ( { SYNOPSYS_UNCONNECTED_10 } ) ,
    .out ( fle_scin ) ) ;
direct_interc direct_interc_10_ (
    .in ( { SYNOPSYS_UNCONNECTED_11 } ) ,
    .out ( fle_clk ) ) ;
endmodule


module mux_tree_size2_mem_17 ( prog_clk , ccff_head , ccff_tail , mem_out , 
    mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_30__45 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_size2_mem_16 ( prog_clk , ccff_head , ccff_tail , mem_out , 
    mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_29__44 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_size2_mem_15 ( prog_clk , ccff_head , ccff_tail , mem_out , 
    mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_28__43 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_23 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_size2_17 ( in , sram , sram_inv , out , p1 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p1 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;

const1_23 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p1 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , .X ( out[0] ) ) ;
endmodule


module const1_22 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_size2_16 ( in , sram , sram_inv , out , p1 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p1 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;

const1_22 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p1 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , .X ( out[0] ) ) ;
endmodule


module const1_21 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_size2_15 ( in , sram , sram_inv , out , p1 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p1 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;

const1_21 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p1 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , .X ( out[0] ) ) ;
endmodule


module logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_11 ( 
    Test_en , clk , ff_D , ff_DI , ff_Q , ff_clk ) ;
input  [0:0] Test_en ;
input  [0:0] clk ;
input  [0:0] ff_D ;
input  [0:0] ff_DI ;
output [0:0] ff_Q ;
input  [0:0] ff_clk ;

sky130_fd_sc_hd__sdfxbp_1 sky130_fd_sc_hd__sdfxbp_1_0_ ( .D ( ff_D[0] ) , 
    .SCD ( ff_DI[0] ) , .SCE ( Test_en[0] ) , .CLK ( clk[0] ) , 
    .Q ( ff_Q[0] ) , .Q_N ( SYNOPSYS_UNCONNECTED_1 ) ) ;
endmodule


module logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_10 ( 
    Test_en , clk , ff_D , ff_DI , ff_Q , ff_clk ) ;
input  [0:0] Test_en ;
input  [0:0] clk ;
input  [0:0] ff_D ;
input  [0:0] ff_DI ;
output [0:0] ff_Q ;
input  [0:0] ff_clk ;

sky130_fd_sc_hd__sdfxbp_1 sky130_fd_sc_hd__sdfxbp_1_0_ ( .D ( ff_D[0] ) , 
    .SCD ( ff_DI[0] ) , .SCE ( Test_en[0] ) , .CLK ( clk[0] ) , 
    .Q ( ff_Q[0] ) , .Q_N ( SYNOPSYS_UNCONNECTED_1 ) ) ;
endmodule


module mux_tree_size2_mem_29 ( prog_clk , ccff_head , ccff_tail , mem_out , 
    mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_27__42 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_20 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_size2_29 ( in , sram , sram_inv , out , p1 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p1 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;

const1_20 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p1 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , .X ( out[0] ) ) ;
endmodule


module frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem_5 ( prog_clk , ccff_head , 
    ccff_tail , mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:16] mem_out ;
output [0:16] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_4_ ( .D ( mem_out[3] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[4] ) , .Q_N ( mem_outb[4] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_5_ ( .D ( mem_out[4] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[5] ) , .Q_N ( mem_outb[5] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_6_ ( .D ( mem_out[5] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[6] ) , .Q_N ( mem_outb[6] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_7_ ( .D ( mem_out[6] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[7] ) , .Q_N ( mem_outb[7] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_8_ ( .D ( mem_out[7] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[8] ) , .Q_N ( mem_outb[8] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_9_ ( .D ( mem_out[8] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[9] ) , .Q_N ( mem_outb[9] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_10_ ( .D ( mem_out[9] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[10] ) , .Q_N ( mem_outb[10] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_11_ ( .D ( mem_out[10] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[11] ) , .Q_N ( mem_outb[11] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_12_ ( .D ( mem_out[11] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[12] ) , .Q_N ( mem_outb[12] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_13_ ( .D ( mem_out[12] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[13] ) , .Q_N ( mem_outb[13] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_14_ ( .D ( mem_out[13] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[14] ) , .Q_N ( mem_outb[14] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_15_ ( .D ( mem_out[14] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[15] ) , .Q_N ( mem_outb[15] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_16_ ( .D ( mem_out[15] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[16] ) , .Q_N ( \_gOb5_mem_outb[16] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_26__41 ( .A ( mem_out[16] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module frac_lut4_mux_5 ( in , sram , sram_inv , lut3_out , lut4_out ) ;
input  [0:15] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:1] lut3_out ;
output [0:0] lut4_out ;

wire [0:0] sky130_fd_sc_hd__buf_2_3_X ;
wire [0:0] sky130_fd_sc_hd__buf_2_4_X ;
wire [0:0] sky130_fd_sc_hd__buf_2_5_X ;
wire [0:0] sky130_fd_sc_hd__buf_2_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_10_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_11_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_12_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_13_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_14_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_12_X[0] ) , .X ( lut3_out[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_1_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_13_X[0] ) , .X ( lut3_out[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_2_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_14_X[0] ) , .X ( lut4_out[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_3_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .X ( sky130_fd_sc_hd__buf_2_3_X[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_4_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , 
    .X ( sky130_fd_sc_hd__buf_2_4_X[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_5_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_10_X[0] ) , 
    .X ( sky130_fd_sc_hd__buf_2_5_X[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_6_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_11_X[0] ) , 
    .X ( sky130_fd_sc_hd__buf_2_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_3_ ( .A0 ( in[7] ) , .A1 ( in[6] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_4_ ( .A0 ( in[9] ) , .A1 ( in[8] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_5_ ( .A0 ( in[11] ) , .A1 ( in[10] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_6_ ( .A0 ( in[13] ) , .A1 ( in[12] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_7_ ( .A0 ( in[15] ) , .A1 ( in[14] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_10_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_11_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( .A0 ( sky130_fd_sc_hd__buf_2_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__buf_2_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_12_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( .A0 ( sky130_fd_sc_hd__buf_2_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__buf_2_5_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_13_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_13_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_12_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_14_X[0] ) ) ;
endmodule


module frac_lut4_5 ( in , sram , sram_inv , mode , mode_inv , lut3_out , 
    lut4_out ) ;
input  [0:3] in ;
input  [0:15] sram ;
input  [0:15] sram_inv ;
input  [0:0] mode ;
input  [0:0] mode_inv ;
output [0:1] lut3_out ;
output [0:0] lut4_out ;

wire [0:0] sky130_fd_sc_hd__buf_2_0_X ;
wire [0:0] sky130_fd_sc_hd__buf_2_1_X ;
wire [0:0] sky130_fd_sc_hd__buf_2_2_X ;
wire [0:0] sky130_fd_sc_hd__buf_2_3_X ;
wire [0:0] sky130_fd_sc_hd__inv_1_0_Y ;
wire [0:0] sky130_fd_sc_hd__inv_1_1_Y ;
wire [0:0] sky130_fd_sc_hd__inv_1_2_Y ;
wire [0:0] sky130_fd_sc_hd__inv_1_3_Y ;
wire [0:0] sky130_fd_sc_hd__or2_1_0_X ;

sky130_fd_sc_hd__or2_0 sky130_fd_sc_hd__or2_1_0_ ( .A ( mode[0] ) , 
    .B ( in[3] ) , .X ( sky130_fd_sc_hd__or2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__inv_1 sky130_fd_sc_hd__inv_1_0_ ( .A ( in[0] ) , 
    .Y ( sky130_fd_sc_hd__inv_1_0_Y[0] ) ) ;
sky130_fd_sc_hd__inv_1 sky130_fd_sc_hd__inv_1_1_ ( .A ( in[1] ) , 
    .Y ( sky130_fd_sc_hd__inv_1_1_Y[0] ) ) ;
sky130_fd_sc_hd__inv_1 sky130_fd_sc_hd__inv_1_2_ ( .A ( in[2] ) , 
    .Y ( sky130_fd_sc_hd__inv_1_2_Y[0] ) ) ;
sky130_fd_sc_hd__inv_1 sky130_fd_sc_hd__inv_1_3_ ( 
    .A ( sky130_fd_sc_hd__or2_1_0_X[0] ) , 
    .Y ( sky130_fd_sc_hd__inv_1_3_Y[0] ) ) ;
sky130_fd_sc_hd__buf_2 sky130_fd_sc_hd__buf_2_0_ ( .A ( in[0] ) , 
    .X ( sky130_fd_sc_hd__buf_2_0_X[0] ) ) ;
sky130_fd_sc_hd__buf_2 sky130_fd_sc_hd__buf_2_1_ ( .A ( in[1] ) , 
    .X ( sky130_fd_sc_hd__buf_2_1_X[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_2_ ( .A ( in[2] ) , 
    .X ( sky130_fd_sc_hd__buf_2_2_X[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_3_ ( 
    .A ( sky130_fd_sc_hd__or2_1_0_X[0] ) , 
    .X ( sky130_fd_sc_hd__buf_2_3_X[0] ) ) ;
frac_lut4_mux_5 frac_lut4_mux_0_ ( .in ( sram ) ,
    .sram ( { sky130_fd_sc_hd__buf_2_0_X[0] , sky130_fd_sc_hd__buf_2_1_X[0] , 
        sky130_fd_sc_hd__buf_2_2_X[0] , sky130_fd_sc_hd__buf_2_3_X[0] } ) ,
    .sram_inv ( { sky130_fd_sc_hd__inv_1_0_Y[0] , 
        sky130_fd_sc_hd__inv_1_1_Y[0] , sky130_fd_sc_hd__inv_1_2_Y[0] , 
        sky130_fd_sc_hd__inv_1_3_Y[0] } ) ,
    .lut3_out ( lut3_out ) , .lut4_out ( lut4_out ) ) ;
endmodule


module logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_5 ( 
    prog_clk , frac_lut4_in , ccff_head , frac_lut4_lut3_out , 
    frac_lut4_lut4_out , ccff_tail ) ;
input  [0:0] prog_clk ;
input  [0:3] frac_lut4_in ;
input  [0:0] ccff_head ;
output [0:1] frac_lut4_lut3_out ;
output [0:0] frac_lut4_lut4_out ;
output [0:0] ccff_tail ;

wire [0:0] frac_lut4_0_mode ;
wire [0:15] frac_lut4_0_sram ;
wire [0:15] frac_lut4_0_sram_inv ;

frac_lut4_5 frac_lut4_0_ ( .in ( frac_lut4_in ) , .sram ( frac_lut4_0_sram ) , 
    .sram_inv ( frac_lut4_0_sram_inv ) , .mode ( frac_lut4_0_mode ) ,
    .mode_inv ( { SYNOPSYS_UNCONNECTED_1 } ) ,
    .lut3_out ( frac_lut4_lut3_out ) , .lut4_out ( frac_lut4_lut4_out ) ) ;
frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem_5 frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem ( 
    .prog_clk ( prog_clk ) , .ccff_head ( ccff_head ) , 
    .ccff_tail ( ccff_tail ) ,
    .mem_out ( { frac_lut4_0_sram[0] , frac_lut4_0_sram[1] , 
        frac_lut4_0_sram[2] , frac_lut4_0_sram[3] , frac_lut4_0_sram[4] , 
        frac_lut4_0_sram[5] , frac_lut4_0_sram[6] , frac_lut4_0_sram[7] , 
        frac_lut4_0_sram[8] , frac_lut4_0_sram[9] , frac_lut4_0_sram[10] , 
        frac_lut4_0_sram[11] , frac_lut4_0_sram[12] , frac_lut4_0_sram[13] , 
        frac_lut4_0_sram[14] , frac_lut4_0_sram[15] , frac_lut4_0_mode[0] } ) ,
    .mem_outb ( { frac_lut4_0_sram_inv[0] , frac_lut4_0_sram_inv[1] , 
        frac_lut4_0_sram_inv[2] , frac_lut4_0_sram_inv[3] , 
        frac_lut4_0_sram_inv[4] , frac_lut4_0_sram_inv[5] , 
        frac_lut4_0_sram_inv[6] , frac_lut4_0_sram_inv[7] , 
        frac_lut4_0_sram_inv[8] , frac_lut4_0_sram_inv[9] , 
        frac_lut4_0_sram_inv[10] , frac_lut4_0_sram_inv[11] , 
        frac_lut4_0_sram_inv[12] , frac_lut4_0_sram_inv[13] , 
        frac_lut4_0_sram_inv[14] , frac_lut4_0_sram_inv[15] , 
        SYNOPSYS_UNCONNECTED_2 } ) ) ;
endmodule


module logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_5 ( 
    prog_clk , frac_logic_in , ccff_head , frac_logic_out , ccff_tail , p1 ) ;
input  [0:0] prog_clk ;
input  [0:3] frac_logic_in ;
input  [0:0] ccff_head ;
output [0:1] frac_logic_out ;
output [0:0] ccff_tail ;
input  p1 ;

wire [0:0] logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_ccff_tail ;
wire [0:0] logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_frac_lut4_lut3_out ;
wire [0:0] logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_frac_lut4_lut4_out ;
wire [0:1] mux_tree_size2_0_sram ;
wire [0:1] mux_tree_size2_0_sram_inv ;

logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_5 logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0 ( 
    .prog_clk ( prog_clk ) , .frac_lut4_in ( frac_logic_in ) , 
    .ccff_head ( ccff_head ) ,
    .frac_lut4_lut3_out ( { 
        logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_frac_lut4_lut3_out[0] , 
        frac_logic_out[1] } ) ,
    
    .frac_lut4_lut4_out ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_frac_lut4_lut4_out ) , 
    .ccff_tail ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_ccff_tail ) ) ;
mux_tree_size2_29 mux_frac_logic_out_0 (
    .in ( { 
        logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_frac_lut4_lut4_out[0] , 
        logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_frac_lut4_lut3_out[0]
         } ) ,
    .sram ( mux_tree_size2_0_sram ) , 
    .sram_inv ( mux_tree_size2_0_sram_inv ) , .out ( frac_logic_out[0] ) , 
    .p1 ( p1 ) ) ;
mux_tree_size2_mem_29 mem_frac_logic_out_0 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_ccff_tail ) , 
    .ccff_tail ( ccff_tail ) , .mem_out ( mux_tree_size2_0_sram ) , 
    .mem_outb ( mux_tree_size2_0_sram_inv ) ) ;
direct_interc direct_interc_0_ (
    .in ( { SYNOPSYS_UNCONNECTED_1 } ) ,
    .out ( frac_logic_out[1] ) ) ;
direct_interc direct_interc_1_ (
    .in ( { SYNOPSYS_UNCONNECTED_2 } ) ,
    .out ( frac_logic_in[0] ) ) ;
direct_interc direct_interc_2_ (
    .in ( { SYNOPSYS_UNCONNECTED_3 } ) ,
    .out ( frac_logic_in[1] ) ) ;
direct_interc direct_interc_3_ (
    .in ( { SYNOPSYS_UNCONNECTED_4 } ) ,
    .out ( frac_logic_in[2] ) ) ;
direct_interc direct_interc_4_ (
    .in ( { SYNOPSYS_UNCONNECTED_5 } ) ,
    .out ( frac_logic_in[3] ) ) ;
endmodule


module logical_tile_clb_mode_default__fle_mode_physical__fabric_5 ( prog_clk , 
    Test_en , clk , fabric_in , fabric_regin , fabric_scin , fabric_clk , 
    ccff_head , fabric_out , fabric_regout , fabric_scout , ccff_tail , p1 ) ;
input  [0:0] prog_clk ;
input  [0:0] Test_en ;
input  [0:0] clk ;
input  [0:3] fabric_in ;
input  [0:0] fabric_regin ;
input  [0:0] fabric_scin ;
input  [0:0] fabric_clk ;
input  [0:0] ccff_head ;
output [0:1] fabric_out ;
output [0:0] fabric_regout ;
output [0:0] fabric_scout ;
output [0:0] ccff_tail ;
input  p1 ;

wire [0:0] logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0_ff_Q ;
wire [0:0] logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_ccff_tail ;
wire [0:1] logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_frac_logic_out ;
wire [0:1] mux_tree_size2_0_sram ;
wire [0:1] mux_tree_size2_0_sram_inv ;
wire [0:1] mux_tree_size2_1_sram ;
wire [0:1] mux_tree_size2_1_sram_inv ;
wire [0:0] mux_tree_size2_2_out ;
wire [0:1] mux_tree_size2_2_sram ;
wire [0:1] mux_tree_size2_2_sram_inv ;
wire [0:0] mux_tree_size2_mem_0_ccff_tail ;
wire [0:0] mux_tree_size2_mem_1_ccff_tail ;

assign fabric_regout[0] = fabric_scout[0] ;

logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_5 logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0 ( 
    .prog_clk ( prog_clk ) , .frac_logic_in ( fabric_in ) , 
    .ccff_head ( ccff_head ) , 
    .frac_logic_out ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_frac_logic_out ) , 
    .ccff_tail ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_ccff_tail ) , 
    .p1 ( p1 ) ) ;
logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_10 logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0 ( 
    .Test_en ( Test_en ) , .clk ( clk ) , .ff_D ( mux_tree_size2_2_out ) , 
    .ff_DI ( fabric_scin ) , 
    .ff_Q ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0_ff_Q ) ,
    .ff_clk ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_11 logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1 ( 
    .Test_en ( Test_en ) , .clk ( clk ) , 
    .ff_D ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_frac_logic_out[1] ) , 
    .ff_DI ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0_ff_Q ) , 
    .ff_Q ( fabric_scout ) ,
    .ff_clk ( { SYNOPSYS_UNCONNECTED_2 } ) ) ;
mux_tree_size2_15 mux_fabric_out_0 (
    .in ( { 
        logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0_ff_Q[0] , 
        logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_frac_logic_out[0]
         } ) ,
    .sram ( mux_tree_size2_0_sram ) , 
    .sram_inv ( mux_tree_size2_0_sram_inv ) , .out ( fabric_out[0] ) , 
    .p1 ( p1 ) ) ;
mux_tree_size2_16 mux_fabric_out_1 (
    .in ( { fabric_scout[0] , 
        logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_frac_logic_out[1]
         } ) ,
    .sram ( mux_tree_size2_1_sram ) , 
    .sram_inv ( mux_tree_size2_1_sram_inv ) , .out ( fabric_out[1] ) , 
    .p1 ( p1 ) ) ;
mux_tree_size2_17 mux_ff_0_D_0 (
    .in ( { 
        logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_frac_logic_out[0] , 
        fabric_regin[0] } ) ,
    .sram ( mux_tree_size2_2_sram ) , 
    .sram_inv ( mux_tree_size2_2_sram_inv ) , .out ( mux_tree_size2_2_out ) , 
    .p1 ( p1 ) ) ;
mux_tree_size2_mem_15 mem_fabric_out_0 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_size2_mem_0_ccff_tail ) , 
    .mem_out ( mux_tree_size2_0_sram ) , 
    .mem_outb ( mux_tree_size2_0_sram_inv ) ) ;
mux_tree_size2_mem_16 mem_fabric_out_1 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_size2_mem_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_size2_mem_1_ccff_tail ) , 
    .mem_out ( mux_tree_size2_1_sram ) , 
    .mem_outb ( mux_tree_size2_1_sram_inv ) ) ;
mux_tree_size2_mem_17 mem_ff_0_D_0 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_size2_mem_1_ccff_tail ) , .ccff_tail ( ccff_tail ) , 
    .mem_out ( mux_tree_size2_2_sram ) , 
    .mem_outb ( mux_tree_size2_2_sram_inv ) ) ;
direct_interc direct_interc_0_ (
    .in ( { SYNOPSYS_UNCONNECTED_3 } ) ,
    .out ( fabric_scout ) ) ;
direct_interc direct_interc_1_ (
    .in ( { SYNOPSYS_UNCONNECTED_4 } ) ,
    .out ( fabric_scout ) ) ;
direct_interc direct_interc_2_ (
    .in ( { SYNOPSYS_UNCONNECTED_5 } ) ,
    .out ( fabric_in[0] ) ) ;
direct_interc direct_interc_3_ (
    .in ( { SYNOPSYS_UNCONNECTED_6 } ) ,
    .out ( fabric_in[1] ) ) ;
direct_interc direct_interc_4_ (
    .in ( { SYNOPSYS_UNCONNECTED_7 } ) ,
    .out ( fabric_in[2] ) ) ;
direct_interc direct_interc_5_ (
    .in ( { SYNOPSYS_UNCONNECTED_8 } ) ,
    .out ( fabric_in[3] ) ) ;
direct_interc direct_interc_6_ (
    .in ( { SYNOPSYS_UNCONNECTED_9 } ) ,
    .out ( fabric_scin ) ) ;
direct_interc direct_interc_7_ (
    .in ( { SYNOPSYS_UNCONNECTED_10 } ) ,
    .out ( fabric_clk ) ) ;
direct_interc direct_interc_8_ (
    .in ( { SYNOPSYS_UNCONNECTED_11 } ) ,
    
    .out ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_frac_logic_out[1] ) ) ;
direct_interc direct_interc_9_ (
    .in ( { SYNOPSYS_UNCONNECTED_12 } ) ,
    
    .out ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0_ff_Q ) ) ;
direct_interc direct_interc_10_ (
    .in ( { SYNOPSYS_UNCONNECTED_13 } ) ,
    .out ( fabric_clk ) ) ;
endmodule


module logical_tile_clb_mode_default__fle_5 ( prog_clk , Test_en , clk , 
    fle_in , fle_regin , fle_scin , fle_clk , ccff_head , fle_out , 
    fle_regout , fle_scout , ccff_tail , p1 ) ;
input  [0:0] prog_clk ;
input  [0:0] Test_en ;
input  [0:0] clk ;
input  [0:3] fle_in ;
input  [0:0] fle_regin ;
input  [0:0] fle_scin ;
input  [0:0] fle_clk ;
input  [0:0] ccff_head ;
output [0:1] fle_out ;
output [0:0] fle_regout ;
output [0:0] fle_scout ;
output [0:0] ccff_tail ;
input  p1 ;

logical_tile_clb_mode_default__fle_mode_physical__fabric_5 logical_tile_clb_mode_default__fle_mode_physical__fabric_0 ( 
    .prog_clk ( prog_clk ) , .Test_en ( Test_en ) , .clk ( clk ) , 
    .fabric_in ( fle_in ) , .fabric_regin ( fle_regin ) , 
    .fabric_scin ( fle_scin ) , .fabric_clk ( fle_clk ) , 
    .ccff_head ( ccff_head ) , .fabric_out ( fle_out ) , 
    .fabric_regout ( fle_regout ) , .fabric_scout ( fle_scout ) , 
    .ccff_tail ( ccff_tail ) , .p1 ( p1 ) ) ;
direct_interc direct_interc_0_ (
    .in ( { SYNOPSYS_UNCONNECTED_1 } ) ,
    .out ( fle_out[0] ) ) ;
direct_interc direct_interc_1_ (
    .in ( { SYNOPSYS_UNCONNECTED_2 } ) ,
    .out ( fle_out[1] ) ) ;
direct_interc direct_interc_2_ (
    .in ( { SYNOPSYS_UNCONNECTED_3 } ) ,
    .out ( fle_regout ) ) ;
direct_interc direct_interc_3_ (
    .in ( { SYNOPSYS_UNCONNECTED_4 } ) ,
    .out ( fle_scout ) ) ;
direct_interc direct_interc_4_ (
    .in ( { SYNOPSYS_UNCONNECTED_5 } ) ,
    .out ( fle_in[0] ) ) ;
direct_interc direct_interc_5_ (
    .in ( { SYNOPSYS_UNCONNECTED_6 } ) ,
    .out ( fle_in[1] ) ) ;
direct_interc direct_interc_6_ (
    .in ( { SYNOPSYS_UNCONNECTED_7 } ) ,
    .out ( fle_in[2] ) ) ;
direct_interc direct_interc_7_ (
    .in ( { SYNOPSYS_UNCONNECTED_8 } ) ,
    .out ( fle_in[3] ) ) ;
direct_interc direct_interc_8_ (
    .in ( { SYNOPSYS_UNCONNECTED_9 } ) ,
    .out ( fle_regin ) ) ;
direct_interc direct_interc_9_ (
    .in ( { SYNOPSYS_UNCONNECTED_10 } ) ,
    .out ( fle_scin ) ) ;
direct_interc direct_interc_10_ (
    .in ( { SYNOPSYS_UNCONNECTED_11 } ) ,
    .out ( fle_clk ) ) ;
endmodule


module mux_tree_size2_mem_14 ( prog_clk , ccff_head , ccff_tail , mem_out , 
    mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_25__40 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_size2_mem_13 ( prog_clk , ccff_head , ccff_tail , mem_out , 
    mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_24__39 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_size2_mem_12 ( prog_clk , ccff_head , ccff_tail , mem_out , 
    mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_23__38 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_19 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_size2_14 ( in , sram , sram_inv , out , p3 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p3 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;

const1_19 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p3 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , .X ( out[0] ) ) ;
endmodule


module const1_18 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_size2_13 ( in , sram , sram_inv , out , p3 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p3 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;

const1_18 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p3 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , .X ( out[0] ) ) ;
endmodule


module const1_17 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_size2_12 ( in , sram , sram_inv , out , p1 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p1 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;

const1_17 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p1 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , .X ( out[0] ) ) ;
endmodule


module logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_9 ( 
    Test_en , clk , ff_D , ff_DI , ff_Q , ff_clk ) ;
input  [0:0] Test_en ;
input  [0:0] clk ;
input  [0:0] ff_D ;
input  [0:0] ff_DI ;
output [0:0] ff_Q ;
input  [0:0] ff_clk ;

sky130_fd_sc_hd__sdfxbp_1 sky130_fd_sc_hd__sdfxbp_1_0_ ( .D ( ff_D[0] ) , 
    .SCD ( ff_DI[0] ) , .SCE ( Test_en[0] ) , .CLK ( clk[0] ) , 
    .Q ( ff_Q[0] ) , .Q_N ( SYNOPSYS_UNCONNECTED_1 ) ) ;
endmodule


module logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_8 ( 
    Test_en , clk , ff_D , ff_DI , ff_Q , ff_clk ) ;
input  [0:0] Test_en ;
input  [0:0] clk ;
input  [0:0] ff_D ;
input  [0:0] ff_DI ;
output [0:0] ff_Q ;
input  [0:0] ff_clk ;

sky130_fd_sc_hd__sdfxbp_1 sky130_fd_sc_hd__sdfxbp_1_0_ ( .D ( ff_D[0] ) , 
    .SCD ( ff_DI[0] ) , .SCE ( Test_en[0] ) , .CLK ( clk[0] ) , 
    .Q ( ff_Q[0] ) , .Q_N ( SYNOPSYS_UNCONNECTED_1 ) ) ;
endmodule


module mux_tree_size2_mem_28 ( prog_clk , ccff_head , ccff_tail , mem_out , 
    mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_22__37 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_16 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_size2_28 ( in , sram , sram_inv , out , p3 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p3 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;

const1_16 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p3 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , .X ( out[0] ) ) ;
endmodule


module frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem_4 ( prog_clk , ccff_head , 
    ccff_tail , mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:16] mem_out ;
output [0:16] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_4_ ( .D ( mem_out[3] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[4] ) , .Q_N ( mem_outb[4] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_5_ ( .D ( mem_out[4] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[5] ) , .Q_N ( mem_outb[5] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_6_ ( .D ( mem_out[5] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[6] ) , .Q_N ( mem_outb[6] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_7_ ( .D ( mem_out[6] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[7] ) , .Q_N ( mem_outb[7] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_8_ ( .D ( mem_out[7] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[8] ) , .Q_N ( mem_outb[8] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_9_ ( .D ( mem_out[8] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[9] ) , .Q_N ( mem_outb[9] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_10_ ( .D ( mem_out[9] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[10] ) , .Q_N ( mem_outb[10] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_11_ ( .D ( mem_out[10] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[11] ) , .Q_N ( mem_outb[11] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_12_ ( .D ( mem_out[11] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[12] ) , .Q_N ( mem_outb[12] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_13_ ( .D ( mem_out[12] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[13] ) , .Q_N ( mem_outb[13] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_14_ ( .D ( mem_out[13] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[14] ) , .Q_N ( mem_outb[14] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_15_ ( .D ( mem_out[14] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[15] ) , .Q_N ( mem_outb[15] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_16_ ( .D ( mem_out[15] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[16] ) , .Q_N ( \_gOb4_mem_outb[16] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_21__36 ( .A ( mem_out[16] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module frac_lut4_mux_4 ( in , sram , sram_inv , lut3_out , lut4_out ) ;
input  [0:15] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:1] lut3_out ;
output [0:0] lut4_out ;

wire [0:0] sky130_fd_sc_hd__buf_2_3_X ;
wire [0:0] sky130_fd_sc_hd__buf_2_4_X ;
wire [0:0] sky130_fd_sc_hd__buf_2_5_X ;
wire [0:0] sky130_fd_sc_hd__buf_2_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_10_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_11_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_12_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_13_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_14_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_12_X[0] ) , .X ( lut3_out[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_1_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_13_X[0] ) , .X ( lut3_out[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_2_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_14_X[0] ) , .X ( lut4_out[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_3_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .X ( sky130_fd_sc_hd__buf_2_3_X[0] ) ) ;
sky130_fd_sc_hd__buf_2 sky130_fd_sc_hd__buf_2_4_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , 
    .X ( sky130_fd_sc_hd__buf_2_4_X[0] ) ) ;
sky130_fd_sc_hd__buf_2 sky130_fd_sc_hd__buf_2_5_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_10_X[0] ) , 
    .X ( sky130_fd_sc_hd__buf_2_5_X[0] ) ) ;
sky130_fd_sc_hd__buf_2 sky130_fd_sc_hd__buf_2_6_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_11_X[0] ) , 
    .X ( sky130_fd_sc_hd__buf_2_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_3_ ( .A0 ( in[7] ) , .A1 ( in[6] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_4_ ( .A0 ( in[9] ) , .A1 ( in[8] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_5_ ( .A0 ( in[11] ) , .A1 ( in[10] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_6_ ( .A0 ( in[13] ) , .A1 ( in[12] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_7_ ( .A0 ( in[15] ) , .A1 ( in[14] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_10_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_11_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( .A0 ( sky130_fd_sc_hd__buf_2_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__buf_2_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_12_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( .A0 ( sky130_fd_sc_hd__buf_2_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__buf_2_5_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_13_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_13_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_12_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_14_X[0] ) ) ;
endmodule


module frac_lut4_4 ( in , sram , sram_inv , mode , mode_inv , lut3_out , 
    lut4_out ) ;
input  [0:3] in ;
input  [0:15] sram ;
input  [0:15] sram_inv ;
input  [0:0] mode ;
input  [0:0] mode_inv ;
output [0:1] lut3_out ;
output [0:0] lut4_out ;

wire [0:0] sky130_fd_sc_hd__buf_2_0_X ;
wire [0:0] sky130_fd_sc_hd__buf_2_1_X ;
wire [0:0] sky130_fd_sc_hd__buf_2_2_X ;
wire [0:0] sky130_fd_sc_hd__buf_2_3_X ;
wire [0:0] sky130_fd_sc_hd__inv_1_0_Y ;
wire [0:0] sky130_fd_sc_hd__inv_1_1_Y ;
wire [0:0] sky130_fd_sc_hd__inv_1_2_Y ;
wire [0:0] sky130_fd_sc_hd__inv_1_3_Y ;
wire [0:0] sky130_fd_sc_hd__or2_1_0_X ;

sky130_fd_sc_hd__or2_0 sky130_fd_sc_hd__or2_1_0_ ( .A ( mode[0] ) , 
    .B ( in[3] ) , .X ( sky130_fd_sc_hd__or2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__inv_1 sky130_fd_sc_hd__inv_1_0_ ( .A ( in[0] ) , 
    .Y ( sky130_fd_sc_hd__inv_1_0_Y[0] ) ) ;
sky130_fd_sc_hd__inv_1 sky130_fd_sc_hd__inv_1_1_ ( .A ( in[1] ) , 
    .Y ( sky130_fd_sc_hd__inv_1_1_Y[0] ) ) ;
sky130_fd_sc_hd__inv_1 sky130_fd_sc_hd__inv_1_2_ ( .A ( in[2] ) , 
    .Y ( sky130_fd_sc_hd__inv_1_2_Y[0] ) ) ;
sky130_fd_sc_hd__inv_1 sky130_fd_sc_hd__inv_1_3_ ( 
    .A ( sky130_fd_sc_hd__or2_1_0_X[0] ) , 
    .Y ( sky130_fd_sc_hd__inv_1_3_Y[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_0_ ( .A ( in[0] ) , 
    .X ( sky130_fd_sc_hd__buf_2_0_X[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_1_ ( .A ( in[1] ) , 
    .X ( sky130_fd_sc_hd__buf_2_1_X[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_2_ ( .A ( in[2] ) , 
    .X ( sky130_fd_sc_hd__buf_2_2_X[0] ) ) ;
sky130_fd_sc_hd__buf_2 sky130_fd_sc_hd__buf_2_3_ ( 
    .A ( sky130_fd_sc_hd__or2_1_0_X[0] ) , 
    .X ( sky130_fd_sc_hd__buf_2_3_X[0] ) ) ;
frac_lut4_mux_4 frac_lut4_mux_0_ ( .in ( sram ) ,
    .sram ( { sky130_fd_sc_hd__buf_2_0_X[0] , sky130_fd_sc_hd__buf_2_1_X[0] , 
        sky130_fd_sc_hd__buf_2_2_X[0] , sky130_fd_sc_hd__buf_2_3_X[0] } ) ,
    .sram_inv ( { sky130_fd_sc_hd__inv_1_0_Y[0] , 
        sky130_fd_sc_hd__inv_1_1_Y[0] , sky130_fd_sc_hd__inv_1_2_Y[0] , 
        sky130_fd_sc_hd__inv_1_3_Y[0] } ) ,
    .lut3_out ( lut3_out ) , .lut4_out ( lut4_out ) ) ;
endmodule


module logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_4 ( 
    prog_clk , frac_lut4_in , ccff_head , frac_lut4_lut3_out , 
    frac_lut4_lut4_out , ccff_tail ) ;
input  [0:0] prog_clk ;
input  [0:3] frac_lut4_in ;
input  [0:0] ccff_head ;
output [0:1] frac_lut4_lut3_out ;
output [0:0] frac_lut4_lut4_out ;
output [0:0] ccff_tail ;

wire [0:0] frac_lut4_0_mode ;
wire [0:15] frac_lut4_0_sram ;
wire [0:15] frac_lut4_0_sram_inv ;

frac_lut4_4 frac_lut4_0_ ( .in ( frac_lut4_in ) , .sram ( frac_lut4_0_sram ) , 
    .sram_inv ( frac_lut4_0_sram_inv ) , .mode ( frac_lut4_0_mode ) ,
    .mode_inv ( { SYNOPSYS_UNCONNECTED_1 } ) ,
    .lut3_out ( frac_lut4_lut3_out ) , .lut4_out ( frac_lut4_lut4_out ) ) ;
frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem_4 frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem ( 
    .prog_clk ( prog_clk ) , .ccff_head ( ccff_head ) , 
    .ccff_tail ( ccff_tail ) ,
    .mem_out ( { frac_lut4_0_sram[0] , frac_lut4_0_sram[1] , 
        frac_lut4_0_sram[2] , frac_lut4_0_sram[3] , frac_lut4_0_sram[4] , 
        frac_lut4_0_sram[5] , frac_lut4_0_sram[6] , frac_lut4_0_sram[7] , 
        frac_lut4_0_sram[8] , frac_lut4_0_sram[9] , frac_lut4_0_sram[10] , 
        frac_lut4_0_sram[11] , frac_lut4_0_sram[12] , frac_lut4_0_sram[13] , 
        frac_lut4_0_sram[14] , frac_lut4_0_sram[15] , frac_lut4_0_mode[0] } ) ,
    .mem_outb ( { frac_lut4_0_sram_inv[0] , frac_lut4_0_sram_inv[1] , 
        frac_lut4_0_sram_inv[2] , frac_lut4_0_sram_inv[3] , 
        frac_lut4_0_sram_inv[4] , frac_lut4_0_sram_inv[5] , 
        frac_lut4_0_sram_inv[6] , frac_lut4_0_sram_inv[7] , 
        frac_lut4_0_sram_inv[8] , frac_lut4_0_sram_inv[9] , 
        frac_lut4_0_sram_inv[10] , frac_lut4_0_sram_inv[11] , 
        frac_lut4_0_sram_inv[12] , frac_lut4_0_sram_inv[13] , 
        frac_lut4_0_sram_inv[14] , frac_lut4_0_sram_inv[15] , 
        SYNOPSYS_UNCONNECTED_2 } ) ) ;
endmodule


module logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_4 ( 
    prog_clk , frac_logic_in , ccff_head , frac_logic_out , ccff_tail , p3 ) ;
input  [0:0] prog_clk ;
input  [0:3] frac_logic_in ;
input  [0:0] ccff_head ;
output [0:1] frac_logic_out ;
output [0:0] ccff_tail ;
input  p3 ;

wire [0:0] logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_ccff_tail ;
wire [0:0] logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_frac_lut4_lut3_out ;
wire [0:0] logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_frac_lut4_lut4_out ;
wire [0:1] mux_tree_size2_0_sram ;
wire [0:1] mux_tree_size2_0_sram_inv ;

logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_4 logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0 ( 
    .prog_clk ( prog_clk ) , .frac_lut4_in ( frac_logic_in ) , 
    .ccff_head ( ccff_head ) ,
    .frac_lut4_lut3_out ( { 
        logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_frac_lut4_lut3_out[0] , 
        frac_logic_out[1] } ) ,
    
    .frac_lut4_lut4_out ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_frac_lut4_lut4_out ) , 
    .ccff_tail ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_ccff_tail ) ) ;
mux_tree_size2_28 mux_frac_logic_out_0 (
    .in ( { 
        logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_frac_lut4_lut4_out[0] , 
        logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_frac_lut4_lut3_out[0]
         } ) ,
    .sram ( mux_tree_size2_0_sram ) , 
    .sram_inv ( mux_tree_size2_0_sram_inv ) , .out ( frac_logic_out[0] ) , 
    .p3 ( p3 ) ) ;
mux_tree_size2_mem_28 mem_frac_logic_out_0 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_ccff_tail ) , 
    .ccff_tail ( ccff_tail ) , .mem_out ( mux_tree_size2_0_sram ) , 
    .mem_outb ( mux_tree_size2_0_sram_inv ) ) ;
direct_interc direct_interc_0_ (
    .in ( { SYNOPSYS_UNCONNECTED_1 } ) ,
    .out ( frac_logic_out[1] ) ) ;
direct_interc direct_interc_1_ (
    .in ( { SYNOPSYS_UNCONNECTED_2 } ) ,
    .out ( frac_logic_in[0] ) ) ;
direct_interc direct_interc_2_ (
    .in ( { SYNOPSYS_UNCONNECTED_3 } ) ,
    .out ( frac_logic_in[1] ) ) ;
direct_interc direct_interc_3_ (
    .in ( { SYNOPSYS_UNCONNECTED_4 } ) ,
    .out ( frac_logic_in[2] ) ) ;
direct_interc direct_interc_4_ (
    .in ( { SYNOPSYS_UNCONNECTED_5 } ) ,
    .out ( frac_logic_in[3] ) ) ;
endmodule


module logical_tile_clb_mode_default__fle_mode_physical__fabric_4 ( prog_clk , 
    Test_en , clk , fabric_in , fabric_regin , fabric_scin , fabric_clk , 
    ccff_head , fabric_out , fabric_regout , fabric_scout , ccff_tail , p1 , 
    p3 ) ;
input  [0:0] prog_clk ;
input  [0:0] Test_en ;
input  [0:0] clk ;
input  [0:3] fabric_in ;
input  [0:0] fabric_regin ;
input  [0:0] fabric_scin ;
input  [0:0] fabric_clk ;
input  [0:0] ccff_head ;
output [0:1] fabric_out ;
output [0:0] fabric_regout ;
output [0:0] fabric_scout ;
output [0:0] ccff_tail ;
input  p1 ;
input  p3 ;

wire [0:0] logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0_ff_Q ;
wire [0:0] logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_ccff_tail ;
wire [0:1] logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_frac_logic_out ;
wire [0:1] mux_tree_size2_0_sram ;
wire [0:1] mux_tree_size2_0_sram_inv ;
wire [0:1] mux_tree_size2_1_sram ;
wire [0:1] mux_tree_size2_1_sram_inv ;
wire [0:0] mux_tree_size2_2_out ;
wire [0:1] mux_tree_size2_2_sram ;
wire [0:1] mux_tree_size2_2_sram_inv ;
wire [0:0] mux_tree_size2_mem_0_ccff_tail ;
wire [0:0] mux_tree_size2_mem_1_ccff_tail ;

assign fabric_regout[0] = fabric_scout[0] ;

logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_4 logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0 ( 
    .prog_clk ( prog_clk ) , .frac_logic_in ( fabric_in ) , 
    .ccff_head ( ccff_head ) , 
    .frac_logic_out ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_frac_logic_out ) , 
    .ccff_tail ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_ccff_tail ) , 
    .p3 ( p3 ) ) ;
logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_8 logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0 ( 
    .Test_en ( Test_en ) , .clk ( clk ) , .ff_D ( mux_tree_size2_2_out ) , 
    .ff_DI ( fabric_scin ) , 
    .ff_Q ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0_ff_Q ) ,
    .ff_clk ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_9 logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1 ( 
    .Test_en ( Test_en ) , .clk ( clk ) , 
    .ff_D ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_frac_logic_out[1] ) , 
    .ff_DI ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0_ff_Q ) , 
    .ff_Q ( fabric_scout ) ,
    .ff_clk ( { SYNOPSYS_UNCONNECTED_2 } ) ) ;
mux_tree_size2_12 mux_fabric_out_0 (
    .in ( { 
        logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0_ff_Q[0] , 
        logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_frac_logic_out[0]
         } ) ,
    .sram ( mux_tree_size2_0_sram ) , 
    .sram_inv ( mux_tree_size2_0_sram_inv ) , .out ( fabric_out[0] ) , 
    .p1 ( p1 ) ) ;
mux_tree_size2_13 mux_fabric_out_1 (
    .in ( { fabric_scout[0] , 
        logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_frac_logic_out[1]
         } ) ,
    .sram ( mux_tree_size2_1_sram ) , 
    .sram_inv ( mux_tree_size2_1_sram_inv ) , .out ( fabric_out[1] ) , 
    .p3 ( p3 ) ) ;
mux_tree_size2_14 mux_ff_0_D_0 (
    .in ( { 
        logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_frac_logic_out[0] , 
        fabric_regin[0] } ) ,
    .sram ( mux_tree_size2_2_sram ) , 
    .sram_inv ( mux_tree_size2_2_sram_inv ) , .out ( mux_tree_size2_2_out ) , 
    .p3 ( p3 ) ) ;
mux_tree_size2_mem_12 mem_fabric_out_0 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_size2_mem_0_ccff_tail ) , 
    .mem_out ( mux_tree_size2_0_sram ) , 
    .mem_outb ( mux_tree_size2_0_sram_inv ) ) ;
mux_tree_size2_mem_13 mem_fabric_out_1 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_size2_mem_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_size2_mem_1_ccff_tail ) , 
    .mem_out ( mux_tree_size2_1_sram ) , 
    .mem_outb ( mux_tree_size2_1_sram_inv ) ) ;
mux_tree_size2_mem_14 mem_ff_0_D_0 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_size2_mem_1_ccff_tail ) , .ccff_tail ( ccff_tail ) , 
    .mem_out ( mux_tree_size2_2_sram ) , 
    .mem_outb ( mux_tree_size2_2_sram_inv ) ) ;
direct_interc direct_interc_0_ (
    .in ( { SYNOPSYS_UNCONNECTED_3 } ) ,
    .out ( fabric_scout ) ) ;
direct_interc direct_interc_1_ (
    .in ( { SYNOPSYS_UNCONNECTED_4 } ) ,
    .out ( fabric_scout ) ) ;
direct_interc direct_interc_2_ (
    .in ( { SYNOPSYS_UNCONNECTED_5 } ) ,
    .out ( fabric_in[0] ) ) ;
direct_interc direct_interc_3_ (
    .in ( { SYNOPSYS_UNCONNECTED_6 } ) ,
    .out ( fabric_in[1] ) ) ;
direct_interc direct_interc_4_ (
    .in ( { SYNOPSYS_UNCONNECTED_7 } ) ,
    .out ( fabric_in[2] ) ) ;
direct_interc direct_interc_5_ (
    .in ( { SYNOPSYS_UNCONNECTED_8 } ) ,
    .out ( fabric_in[3] ) ) ;
direct_interc direct_interc_6_ (
    .in ( { SYNOPSYS_UNCONNECTED_9 } ) ,
    .out ( fabric_scin ) ) ;
direct_interc direct_interc_7_ (
    .in ( { SYNOPSYS_UNCONNECTED_10 } ) ,
    .out ( fabric_clk ) ) ;
direct_interc direct_interc_8_ (
    .in ( { SYNOPSYS_UNCONNECTED_11 } ) ,
    
    .out ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_frac_logic_out[1] ) ) ;
direct_interc direct_interc_9_ (
    .in ( { SYNOPSYS_UNCONNECTED_12 } ) ,
    
    .out ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0_ff_Q ) ) ;
direct_interc direct_interc_10_ (
    .in ( { SYNOPSYS_UNCONNECTED_13 } ) ,
    .out ( fabric_clk ) ) ;
endmodule


module logical_tile_clb_mode_default__fle_4 ( prog_clk , Test_en , clk , 
    fle_in , fle_regin , fle_scin , fle_clk , ccff_head , fle_out , 
    fle_regout , fle_scout , ccff_tail , p1 , p3 ) ;
input  [0:0] prog_clk ;
input  [0:0] Test_en ;
input  [0:0] clk ;
input  [0:3] fle_in ;
input  [0:0] fle_regin ;
input  [0:0] fle_scin ;
input  [0:0] fle_clk ;
input  [0:0] ccff_head ;
output [0:1] fle_out ;
output [0:0] fle_regout ;
output [0:0] fle_scout ;
output [0:0] ccff_tail ;
input  p1 ;
input  p3 ;

logical_tile_clb_mode_default__fle_mode_physical__fabric_4 logical_tile_clb_mode_default__fle_mode_physical__fabric_0 ( 
    .prog_clk ( prog_clk ) , .Test_en ( Test_en ) , .clk ( clk ) , 
    .fabric_in ( fle_in ) , .fabric_regin ( fle_regin ) , 
    .fabric_scin ( fle_scin ) , .fabric_clk ( fle_clk ) , 
    .ccff_head ( ccff_head ) , .fabric_out ( fle_out ) , 
    .fabric_regout ( fle_regout ) , .fabric_scout ( fle_scout ) , 
    .ccff_tail ( ccff_tail ) , .p1 ( p1 ) , .p3 ( p3 ) ) ;
direct_interc direct_interc_0_ (
    .in ( { SYNOPSYS_UNCONNECTED_1 } ) ,
    .out ( fle_out[0] ) ) ;
direct_interc direct_interc_1_ (
    .in ( { SYNOPSYS_UNCONNECTED_2 } ) ,
    .out ( fle_out[1] ) ) ;
direct_interc direct_interc_2_ (
    .in ( { SYNOPSYS_UNCONNECTED_3 } ) ,
    .out ( fle_regout ) ) ;
direct_interc direct_interc_3_ (
    .in ( { SYNOPSYS_UNCONNECTED_4 } ) ,
    .out ( fle_scout ) ) ;
direct_interc direct_interc_4_ (
    .in ( { SYNOPSYS_UNCONNECTED_5 } ) ,
    .out ( fle_in[0] ) ) ;
direct_interc direct_interc_5_ (
    .in ( { SYNOPSYS_UNCONNECTED_6 } ) ,
    .out ( fle_in[1] ) ) ;
direct_interc direct_interc_6_ (
    .in ( { SYNOPSYS_UNCONNECTED_7 } ) ,
    .out ( fle_in[2] ) ) ;
direct_interc direct_interc_7_ (
    .in ( { SYNOPSYS_UNCONNECTED_8 } ) ,
    .out ( fle_in[3] ) ) ;
direct_interc direct_interc_8_ (
    .in ( { SYNOPSYS_UNCONNECTED_9 } ) ,
    .out ( fle_regin ) ) ;
direct_interc direct_interc_9_ (
    .in ( { SYNOPSYS_UNCONNECTED_10 } ) ,
    .out ( fle_scin ) ) ;
direct_interc direct_interc_10_ (
    .in ( { SYNOPSYS_UNCONNECTED_11 } ) ,
    .out ( fle_clk ) ) ;
endmodule


module mux_tree_size2_mem_11 ( prog_clk , ccff_head , ccff_tail , mem_out , 
    mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_20__35 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_size2_mem_10 ( prog_clk , ccff_head , ccff_tail , mem_out , 
    mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_19__34 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_size2_mem_9 ( prog_clk , ccff_head , ccff_tail , mem_out , 
    mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_18__33 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_15 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_size2_11 ( in , sram , sram_inv , out , p3 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p3 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;

const1_15 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p3 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , .X ( out[0] ) ) ;
endmodule


module const1_14 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_size2_10 ( in , sram , sram_inv , out , p3 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p3 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;

const1_14 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p3 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , .X ( out[0] ) ) ;
endmodule


module const1_13 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_size2_9 ( in , sram , sram_inv , out , p3 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p3 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;

const1_13 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p3 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , .X ( out[0] ) ) ;
endmodule


module logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_7 ( 
    Test_en , clk , ff_D , ff_DI , ff_Q , ff_clk ) ;
input  [0:0] Test_en ;
input  [0:0] clk ;
input  [0:0] ff_D ;
input  [0:0] ff_DI ;
output [0:0] ff_Q ;
input  [0:0] ff_clk ;

sky130_fd_sc_hd__sdfxbp_1 sky130_fd_sc_hd__sdfxbp_1_0_ ( .D ( ff_D[0] ) , 
    .SCD ( ff_DI[0] ) , .SCE ( Test_en[0] ) , .CLK ( clk[0] ) , 
    .Q ( ff_Q[0] ) , .Q_N ( SYNOPSYS_UNCONNECTED_1 ) ) ;
endmodule


module logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_6 ( 
    Test_en , clk , ff_D , ff_DI , ff_Q , ff_clk ) ;
input  [0:0] Test_en ;
input  [0:0] clk ;
input  [0:0] ff_D ;
input  [0:0] ff_DI ;
output [0:0] ff_Q ;
input  [0:0] ff_clk ;

sky130_fd_sc_hd__sdfxbp_1 sky130_fd_sc_hd__sdfxbp_1_0_ ( .D ( ff_D[0] ) , 
    .SCD ( ff_DI[0] ) , .SCE ( Test_en[0] ) , .CLK ( clk[0] ) , 
    .Q ( ff_Q[0] ) , .Q_N ( SYNOPSYS_UNCONNECTED_1 ) ) ;
endmodule


module mux_tree_size2_mem_27 ( prog_clk , ccff_head , ccff_tail , mem_out , 
    mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_17__32 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_12 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_size2_27 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;

const1_12 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , .X ( out[0] ) ) ;
endmodule


module frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem_3 ( prog_clk , ccff_head , 
    ccff_tail , mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:16] mem_out ;
output [0:16] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_4_ ( .D ( mem_out[3] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[4] ) , .Q_N ( mem_outb[4] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_5_ ( .D ( mem_out[4] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[5] ) , .Q_N ( mem_outb[5] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_6_ ( .D ( mem_out[5] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[6] ) , .Q_N ( mem_outb[6] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_7_ ( .D ( mem_out[6] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[7] ) , .Q_N ( mem_outb[7] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_8_ ( .D ( mem_out[7] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[8] ) , .Q_N ( mem_outb[8] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_9_ ( .D ( mem_out[8] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[9] ) , .Q_N ( mem_outb[9] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_10_ ( .D ( mem_out[9] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[10] ) , .Q_N ( mem_outb[10] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_11_ ( .D ( mem_out[10] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[11] ) , .Q_N ( mem_outb[11] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_12_ ( .D ( mem_out[11] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[12] ) , .Q_N ( mem_outb[12] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_13_ ( .D ( mem_out[12] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[13] ) , .Q_N ( mem_outb[13] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_14_ ( .D ( mem_out[13] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[14] ) , .Q_N ( mem_outb[14] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_15_ ( .D ( mem_out[14] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[15] ) , .Q_N ( mem_outb[15] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_16_ ( .D ( mem_out[15] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[16] ) , .Q_N ( \_gOb3_mem_outb[16] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_16__31 ( .A ( mem_out[16] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module frac_lut4_mux_3 ( in , sram , sram_inv , lut3_out , lut4_out ) ;
input  [0:15] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:1] lut3_out ;
output [0:0] lut4_out ;

wire [0:0] sky130_fd_sc_hd__buf_2_3_X ;
wire [0:0] sky130_fd_sc_hd__buf_2_4_X ;
wire [0:0] sky130_fd_sc_hd__buf_2_5_X ;
wire [0:0] sky130_fd_sc_hd__buf_2_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_10_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_11_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_12_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_13_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_14_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_12_X[0] ) , .X ( lut3_out[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_1_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_13_X[0] ) , .X ( lut3_out[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_2_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_14_X[0] ) , .X ( lut4_out[0] ) ) ;
sky130_fd_sc_hd__buf_2 sky130_fd_sc_hd__buf_2_3_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .X ( sky130_fd_sc_hd__buf_2_3_X[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_4_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , 
    .X ( sky130_fd_sc_hd__buf_2_4_X[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_5_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_10_X[0] ) , 
    .X ( sky130_fd_sc_hd__buf_2_5_X[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_6_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_11_X[0] ) , 
    .X ( sky130_fd_sc_hd__buf_2_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_3_ ( .A0 ( in[7] ) , .A1 ( in[6] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_4_ ( .A0 ( in[9] ) , .A1 ( in[8] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_5_ ( .A0 ( in[11] ) , .A1 ( in[10] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_6_ ( .A0 ( in[13] ) , .A1 ( in[12] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_7_ ( .A0 ( in[15] ) , .A1 ( in[14] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_10_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_11_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( .A0 ( sky130_fd_sc_hd__buf_2_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__buf_2_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_12_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( .A0 ( sky130_fd_sc_hd__buf_2_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__buf_2_5_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_13_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_13_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_12_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_14_X[0] ) ) ;
endmodule


module frac_lut4_3 ( in , sram , sram_inv , mode , mode_inv , lut3_out , 
    lut4_out ) ;
input  [0:3] in ;
input  [0:15] sram ;
input  [0:15] sram_inv ;
input  [0:0] mode ;
input  [0:0] mode_inv ;
output [0:1] lut3_out ;
output [0:0] lut4_out ;

wire [0:0] sky130_fd_sc_hd__buf_2_0_X ;
wire [0:0] sky130_fd_sc_hd__buf_2_1_X ;
wire [0:0] sky130_fd_sc_hd__buf_2_2_X ;
wire [0:0] sky130_fd_sc_hd__buf_2_3_X ;
wire [0:0] sky130_fd_sc_hd__inv_1_0_Y ;
wire [0:0] sky130_fd_sc_hd__inv_1_1_Y ;
wire [0:0] sky130_fd_sc_hd__inv_1_2_Y ;
wire [0:0] sky130_fd_sc_hd__inv_1_3_Y ;
wire [0:0] sky130_fd_sc_hd__or2_1_0_X ;

sky130_fd_sc_hd__or2_0 sky130_fd_sc_hd__or2_1_0_ ( .A ( mode[0] ) , 
    .B ( in[3] ) , .X ( sky130_fd_sc_hd__or2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__inv_1 sky130_fd_sc_hd__inv_1_0_ ( .A ( in[0] ) , 
    .Y ( sky130_fd_sc_hd__inv_1_0_Y[0] ) ) ;
sky130_fd_sc_hd__inv_1 sky130_fd_sc_hd__inv_1_1_ ( .A ( in[1] ) , 
    .Y ( sky130_fd_sc_hd__inv_1_1_Y[0] ) ) ;
sky130_fd_sc_hd__inv_1 sky130_fd_sc_hd__inv_1_2_ ( .A ( in[2] ) , 
    .Y ( sky130_fd_sc_hd__inv_1_2_Y[0] ) ) ;
sky130_fd_sc_hd__inv_1 sky130_fd_sc_hd__inv_1_3_ ( 
    .A ( sky130_fd_sc_hd__or2_1_0_X[0] ) , 
    .Y ( sky130_fd_sc_hd__inv_1_3_Y[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_0_ ( .A ( in[0] ) , 
    .X ( sky130_fd_sc_hd__buf_2_0_X[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_1_ ( .A ( in[1] ) , 
    .X ( sky130_fd_sc_hd__buf_2_1_X[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_2_ ( .A ( in[2] ) , 
    .X ( sky130_fd_sc_hd__buf_2_2_X[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_3_ ( 
    .A ( sky130_fd_sc_hd__or2_1_0_X[0] ) , 
    .X ( sky130_fd_sc_hd__buf_2_3_X[0] ) ) ;
frac_lut4_mux_3 frac_lut4_mux_0_ ( .in ( sram ) ,
    .sram ( { sky130_fd_sc_hd__buf_2_0_X[0] , sky130_fd_sc_hd__buf_2_1_X[0] , 
        sky130_fd_sc_hd__buf_2_2_X[0] , sky130_fd_sc_hd__buf_2_3_X[0] } ) ,
    .sram_inv ( { sky130_fd_sc_hd__inv_1_0_Y[0] , 
        sky130_fd_sc_hd__inv_1_1_Y[0] , sky130_fd_sc_hd__inv_1_2_Y[0] , 
        sky130_fd_sc_hd__inv_1_3_Y[0] } ) ,
    .lut3_out ( lut3_out ) , .lut4_out ( lut4_out ) ) ;
endmodule


module logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_3 ( 
    prog_clk , frac_lut4_in , ccff_head , frac_lut4_lut3_out , 
    frac_lut4_lut4_out , ccff_tail ) ;
input  [0:0] prog_clk ;
input  [0:3] frac_lut4_in ;
input  [0:0] ccff_head ;
output [0:1] frac_lut4_lut3_out ;
output [0:0] frac_lut4_lut4_out ;
output [0:0] ccff_tail ;

wire [0:0] frac_lut4_0_mode ;
wire [0:15] frac_lut4_0_sram ;
wire [0:15] frac_lut4_0_sram_inv ;

frac_lut4_3 frac_lut4_0_ ( .in ( frac_lut4_in ) , .sram ( frac_lut4_0_sram ) , 
    .sram_inv ( frac_lut4_0_sram_inv ) , .mode ( frac_lut4_0_mode ) ,
    .mode_inv ( { SYNOPSYS_UNCONNECTED_1 } ) ,
    .lut3_out ( frac_lut4_lut3_out ) , .lut4_out ( frac_lut4_lut4_out ) ) ;
frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem_3 frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem ( 
    .prog_clk ( prog_clk ) , .ccff_head ( ccff_head ) , 
    .ccff_tail ( ccff_tail ) ,
    .mem_out ( { frac_lut4_0_sram[0] , frac_lut4_0_sram[1] , 
        frac_lut4_0_sram[2] , frac_lut4_0_sram[3] , frac_lut4_0_sram[4] , 
        frac_lut4_0_sram[5] , frac_lut4_0_sram[6] , frac_lut4_0_sram[7] , 
        frac_lut4_0_sram[8] , frac_lut4_0_sram[9] , frac_lut4_0_sram[10] , 
        frac_lut4_0_sram[11] , frac_lut4_0_sram[12] , frac_lut4_0_sram[13] , 
        frac_lut4_0_sram[14] , frac_lut4_0_sram[15] , frac_lut4_0_mode[0] } ) ,
    .mem_outb ( { frac_lut4_0_sram_inv[0] , frac_lut4_0_sram_inv[1] , 
        frac_lut4_0_sram_inv[2] , frac_lut4_0_sram_inv[3] , 
        frac_lut4_0_sram_inv[4] , frac_lut4_0_sram_inv[5] , 
        frac_lut4_0_sram_inv[6] , frac_lut4_0_sram_inv[7] , 
        frac_lut4_0_sram_inv[8] , frac_lut4_0_sram_inv[9] , 
        frac_lut4_0_sram_inv[10] , frac_lut4_0_sram_inv[11] , 
        frac_lut4_0_sram_inv[12] , frac_lut4_0_sram_inv[13] , 
        frac_lut4_0_sram_inv[14] , frac_lut4_0_sram_inv[15] , 
        SYNOPSYS_UNCONNECTED_2 } ) ) ;
endmodule


module logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_3 ( 
    prog_clk , frac_logic_in , ccff_head , frac_logic_out , ccff_tail , p0 ) ;
input  [0:0] prog_clk ;
input  [0:3] frac_logic_in ;
input  [0:0] ccff_head ;
output [0:1] frac_logic_out ;
output [0:0] ccff_tail ;
input  p0 ;

wire [0:0] logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_ccff_tail ;
wire [0:0] logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_frac_lut4_lut3_out ;
wire [0:0] logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_frac_lut4_lut4_out ;
wire [0:1] mux_tree_size2_0_sram ;
wire [0:1] mux_tree_size2_0_sram_inv ;

logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_3 logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0 ( 
    .prog_clk ( prog_clk ) , .frac_lut4_in ( frac_logic_in ) , 
    .ccff_head ( ccff_head ) ,
    .frac_lut4_lut3_out ( { 
        logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_frac_lut4_lut3_out[0] , 
        frac_logic_out[1] } ) ,
    
    .frac_lut4_lut4_out ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_frac_lut4_lut4_out ) , 
    .ccff_tail ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_ccff_tail ) ) ;
mux_tree_size2_27 mux_frac_logic_out_0 (
    .in ( { 
        logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_frac_lut4_lut4_out[0] , 
        logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_frac_lut4_lut3_out[0]
         } ) ,
    .sram ( mux_tree_size2_0_sram ) , 
    .sram_inv ( mux_tree_size2_0_sram_inv ) , .out ( frac_logic_out[0] ) , 
    .p0 ( p0 ) ) ;
mux_tree_size2_mem_27 mem_frac_logic_out_0 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_ccff_tail ) , 
    .ccff_tail ( ccff_tail ) , .mem_out ( mux_tree_size2_0_sram ) , 
    .mem_outb ( mux_tree_size2_0_sram_inv ) ) ;
direct_interc direct_interc_0_ (
    .in ( { SYNOPSYS_UNCONNECTED_1 } ) ,
    .out ( frac_logic_out[1] ) ) ;
direct_interc direct_interc_1_ (
    .in ( { SYNOPSYS_UNCONNECTED_2 } ) ,
    .out ( frac_logic_in[0] ) ) ;
direct_interc direct_interc_2_ (
    .in ( { SYNOPSYS_UNCONNECTED_3 } ) ,
    .out ( frac_logic_in[1] ) ) ;
direct_interc direct_interc_3_ (
    .in ( { SYNOPSYS_UNCONNECTED_4 } ) ,
    .out ( frac_logic_in[2] ) ) ;
direct_interc direct_interc_4_ (
    .in ( { SYNOPSYS_UNCONNECTED_5 } ) ,
    .out ( frac_logic_in[3] ) ) ;
endmodule


module logical_tile_clb_mode_default__fle_mode_physical__fabric_3 ( prog_clk , 
    Test_en , clk , fabric_in , fabric_regin , fabric_scin , fabric_clk , 
    ccff_head , fabric_out , fabric_regout , fabric_scout , ccff_tail , p0 , 
    p3 ) ;
input  [0:0] prog_clk ;
input  [0:0] Test_en ;
input  [0:0] clk ;
input  [0:3] fabric_in ;
input  [0:0] fabric_regin ;
input  [0:0] fabric_scin ;
input  [0:0] fabric_clk ;
input  [0:0] ccff_head ;
output [0:1] fabric_out ;
output [0:0] fabric_regout ;
output [0:0] fabric_scout ;
output [0:0] ccff_tail ;
input  p0 ;
input  p3 ;

wire [0:0] logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0_ff_Q ;
wire [0:0] logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_ccff_tail ;
wire [0:1] logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_frac_logic_out ;
wire [0:1] mux_tree_size2_0_sram ;
wire [0:1] mux_tree_size2_0_sram_inv ;
wire [0:1] mux_tree_size2_1_sram ;
wire [0:1] mux_tree_size2_1_sram_inv ;
wire [0:0] mux_tree_size2_2_out ;
wire [0:1] mux_tree_size2_2_sram ;
wire [0:1] mux_tree_size2_2_sram_inv ;
wire [0:0] mux_tree_size2_mem_0_ccff_tail ;
wire [0:0] mux_tree_size2_mem_1_ccff_tail ;

assign fabric_regout[0] = fabric_scout[0] ;

logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_3 logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0 ( 
    .prog_clk ( prog_clk ) , .frac_logic_in ( fabric_in ) , 
    .ccff_head ( ccff_head ) , 
    .frac_logic_out ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_frac_logic_out ) , 
    .ccff_tail ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_ccff_tail ) , 
    .p0 ( p0 ) ) ;
logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_6 logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0 ( 
    .Test_en ( Test_en ) , .clk ( clk ) , .ff_D ( mux_tree_size2_2_out ) , 
    .ff_DI ( fabric_scin ) , 
    .ff_Q ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0_ff_Q ) ,
    .ff_clk ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_7 logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1 ( 
    .Test_en ( Test_en ) , .clk ( clk ) , 
    .ff_D ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_frac_logic_out[1] ) , 
    .ff_DI ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0_ff_Q ) , 
    .ff_Q ( fabric_scout ) ,
    .ff_clk ( { SYNOPSYS_UNCONNECTED_2 } ) ) ;
mux_tree_size2_9 mux_fabric_out_0 (
    .in ( { 
        logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0_ff_Q[0] , 
        logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_frac_logic_out[0]
         } ) ,
    .sram ( mux_tree_size2_0_sram ) , 
    .sram_inv ( mux_tree_size2_0_sram_inv ) , .out ( fabric_out[0] ) , 
    .p3 ( p3 ) ) ;
mux_tree_size2_10 mux_fabric_out_1 (
    .in ( { fabric_scout[0] , 
        logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_frac_logic_out[1]
         } ) ,
    .sram ( mux_tree_size2_1_sram ) , 
    .sram_inv ( mux_tree_size2_1_sram_inv ) , .out ( fabric_out[1] ) , 
    .p3 ( p3 ) ) ;
mux_tree_size2_11 mux_ff_0_D_0 (
    .in ( { 
        logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_frac_logic_out[0] , 
        fabric_regin[0] } ) ,
    .sram ( mux_tree_size2_2_sram ) , 
    .sram_inv ( mux_tree_size2_2_sram_inv ) , .out ( mux_tree_size2_2_out ) , 
    .p3 ( p3 ) ) ;
mux_tree_size2_mem_9 mem_fabric_out_0 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_size2_mem_0_ccff_tail ) , 
    .mem_out ( mux_tree_size2_0_sram ) , 
    .mem_outb ( mux_tree_size2_0_sram_inv ) ) ;
mux_tree_size2_mem_10 mem_fabric_out_1 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_size2_mem_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_size2_mem_1_ccff_tail ) , 
    .mem_out ( mux_tree_size2_1_sram ) , 
    .mem_outb ( mux_tree_size2_1_sram_inv ) ) ;
mux_tree_size2_mem_11 mem_ff_0_D_0 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_size2_mem_1_ccff_tail ) , .ccff_tail ( ccff_tail ) , 
    .mem_out ( mux_tree_size2_2_sram ) , 
    .mem_outb ( mux_tree_size2_2_sram_inv ) ) ;
direct_interc direct_interc_0_ (
    .in ( { SYNOPSYS_UNCONNECTED_3 } ) ,
    .out ( fabric_scout ) ) ;
direct_interc direct_interc_1_ (
    .in ( { SYNOPSYS_UNCONNECTED_4 } ) ,
    .out ( fabric_scout ) ) ;
direct_interc direct_interc_2_ (
    .in ( { SYNOPSYS_UNCONNECTED_5 } ) ,
    .out ( fabric_in[0] ) ) ;
direct_interc direct_interc_3_ (
    .in ( { SYNOPSYS_UNCONNECTED_6 } ) ,
    .out ( fabric_in[1] ) ) ;
direct_interc direct_interc_4_ (
    .in ( { SYNOPSYS_UNCONNECTED_7 } ) ,
    .out ( fabric_in[2] ) ) ;
direct_interc direct_interc_5_ (
    .in ( { SYNOPSYS_UNCONNECTED_8 } ) ,
    .out ( fabric_in[3] ) ) ;
direct_interc direct_interc_6_ (
    .in ( { SYNOPSYS_UNCONNECTED_9 } ) ,
    .out ( fabric_scin ) ) ;
direct_interc direct_interc_7_ (
    .in ( { SYNOPSYS_UNCONNECTED_10 } ) ,
    .out ( fabric_clk ) ) ;
direct_interc direct_interc_8_ (
    .in ( { SYNOPSYS_UNCONNECTED_11 } ) ,
    
    .out ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_frac_logic_out[1] ) ) ;
direct_interc direct_interc_9_ (
    .in ( { SYNOPSYS_UNCONNECTED_12 } ) ,
    
    .out ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0_ff_Q ) ) ;
direct_interc direct_interc_10_ (
    .in ( { SYNOPSYS_UNCONNECTED_13 } ) ,
    .out ( fabric_clk ) ) ;
endmodule


module logical_tile_clb_mode_default__fle_3 ( prog_clk , Test_en , clk , 
    fle_in , fle_regin , fle_scin , fle_clk , ccff_head , fle_out , 
    fle_regout , fle_scout , ccff_tail , p0 , p3 ) ;
input  [0:0] prog_clk ;
input  [0:0] Test_en ;
input  [0:0] clk ;
input  [0:3] fle_in ;
input  [0:0] fle_regin ;
input  [0:0] fle_scin ;
input  [0:0] fle_clk ;
input  [0:0] ccff_head ;
output [0:1] fle_out ;
output [0:0] fle_regout ;
output [0:0] fle_scout ;
output [0:0] ccff_tail ;
input  p0 ;
input  p3 ;

logical_tile_clb_mode_default__fle_mode_physical__fabric_3 logical_tile_clb_mode_default__fle_mode_physical__fabric_0 ( 
    .prog_clk ( prog_clk ) , .Test_en ( Test_en ) , .clk ( clk ) , 
    .fabric_in ( fle_in ) , .fabric_regin ( fle_regin ) , 
    .fabric_scin ( fle_scin ) , .fabric_clk ( fle_clk ) , 
    .ccff_head ( ccff_head ) , .fabric_out ( fle_out ) , 
    .fabric_regout ( fle_regout ) , .fabric_scout ( fle_scout ) , 
    .ccff_tail ( ccff_tail ) , .p0 ( p0 ) , .p3 ( p3 ) ) ;
direct_interc direct_interc_0_ (
    .in ( { SYNOPSYS_UNCONNECTED_1 } ) ,
    .out ( fle_out[0] ) ) ;
direct_interc direct_interc_1_ (
    .in ( { SYNOPSYS_UNCONNECTED_2 } ) ,
    .out ( fle_out[1] ) ) ;
direct_interc direct_interc_2_ (
    .in ( { SYNOPSYS_UNCONNECTED_3 } ) ,
    .out ( fle_regout ) ) ;
direct_interc direct_interc_3_ (
    .in ( { SYNOPSYS_UNCONNECTED_4 } ) ,
    .out ( fle_scout ) ) ;
direct_interc direct_interc_4_ (
    .in ( { SYNOPSYS_UNCONNECTED_5 } ) ,
    .out ( fle_in[0] ) ) ;
direct_interc direct_interc_5_ (
    .in ( { SYNOPSYS_UNCONNECTED_6 } ) ,
    .out ( fle_in[1] ) ) ;
direct_interc direct_interc_6_ (
    .in ( { SYNOPSYS_UNCONNECTED_7 } ) ,
    .out ( fle_in[2] ) ) ;
direct_interc direct_interc_7_ (
    .in ( { SYNOPSYS_UNCONNECTED_8 } ) ,
    .out ( fle_in[3] ) ) ;
direct_interc direct_interc_8_ (
    .in ( { SYNOPSYS_UNCONNECTED_9 } ) ,
    .out ( fle_regin ) ) ;
direct_interc direct_interc_9_ (
    .in ( { SYNOPSYS_UNCONNECTED_10 } ) ,
    .out ( fle_scin ) ) ;
direct_interc direct_interc_10_ (
    .in ( { SYNOPSYS_UNCONNECTED_11 } ) ,
    .out ( fle_clk ) ) ;
endmodule


module mux_tree_size2_mem_8 ( prog_clk , ccff_head , ccff_tail , mem_out , 
    mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_15__30 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_size2_mem_7 ( prog_clk , ccff_head , ccff_tail , mem_out , 
    mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_14__29 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_size2_mem_6 ( prog_clk , ccff_head , ccff_tail , mem_out , 
    mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_13__28 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_11 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_size2_8 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;

const1_11 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , .X ( out[0] ) ) ;
endmodule


module const1_10 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_size2_7 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;

const1_10 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , .X ( out[0] ) ) ;
endmodule


module const1_9 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_size2_6 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;

const1_9 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , .X ( out[0] ) ) ;
endmodule


module logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_5 ( 
    Test_en , clk , ff_D , ff_DI , ff_Q , ff_clk ) ;
input  [0:0] Test_en ;
input  [0:0] clk ;
input  [0:0] ff_D ;
input  [0:0] ff_DI ;
output [0:0] ff_Q ;
input  [0:0] ff_clk ;

sky130_fd_sc_hd__sdfxbp_1 sky130_fd_sc_hd__sdfxbp_1_0_ ( .D ( ff_D[0] ) , 
    .SCD ( ff_DI[0] ) , .SCE ( Test_en[0] ) , .CLK ( clk[0] ) , 
    .Q ( ff_Q[0] ) , .Q_N ( SYNOPSYS_UNCONNECTED_1 ) ) ;
endmodule


module logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_4 ( 
    Test_en , clk , ff_D , ff_DI , ff_Q , ff_clk ) ;
input  [0:0] Test_en ;
input  [0:0] clk ;
input  [0:0] ff_D ;
input  [0:0] ff_DI ;
output [0:0] ff_Q ;
input  [0:0] ff_clk ;

sky130_fd_sc_hd__sdfxbp_1 sky130_fd_sc_hd__sdfxbp_1_0_ ( .D ( ff_D[0] ) , 
    .SCD ( ff_DI[0] ) , .SCE ( Test_en[0] ) , .CLK ( clk[0] ) , 
    .Q ( ff_Q[0] ) , .Q_N ( SYNOPSYS_UNCONNECTED_1 ) ) ;
endmodule


module mux_tree_size2_mem_26 ( prog_clk , ccff_head , ccff_tail , mem_out , 
    mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_12__27 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_8 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_size2_26 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;

const1_8 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , .X ( out[0] ) ) ;
endmodule


module frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem_2 ( prog_clk , ccff_head , 
    ccff_tail , mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:16] mem_out ;
output [0:16] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_4_ ( .D ( mem_out[3] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[4] ) , .Q_N ( mem_outb[4] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_5_ ( .D ( mem_out[4] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[5] ) , .Q_N ( mem_outb[5] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_6_ ( .D ( mem_out[5] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[6] ) , .Q_N ( mem_outb[6] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_7_ ( .D ( mem_out[6] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[7] ) , .Q_N ( mem_outb[7] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_8_ ( .D ( mem_out[7] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[8] ) , .Q_N ( mem_outb[8] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_9_ ( .D ( mem_out[8] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[9] ) , .Q_N ( mem_outb[9] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_10_ ( .D ( mem_out[9] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[10] ) , .Q_N ( mem_outb[10] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_11_ ( .D ( mem_out[10] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[11] ) , .Q_N ( mem_outb[11] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_12_ ( .D ( mem_out[11] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[12] ) , .Q_N ( mem_outb[12] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_13_ ( .D ( mem_out[12] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[13] ) , .Q_N ( mem_outb[13] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_14_ ( .D ( mem_out[13] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[14] ) , .Q_N ( mem_outb[14] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_15_ ( .D ( mem_out[14] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[15] ) , .Q_N ( mem_outb[15] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_16_ ( .D ( mem_out[15] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[16] ) , .Q_N ( \_gOb2_mem_outb[16] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_11__26 ( .A ( mem_out[16] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module frac_lut4_mux_2 ( in , sram , sram_inv , lut3_out , lut4_out ) ;
input  [0:15] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:1] lut3_out ;
output [0:0] lut4_out ;

wire [0:0] sky130_fd_sc_hd__buf_2_3_X ;
wire [0:0] sky130_fd_sc_hd__buf_2_4_X ;
wire [0:0] sky130_fd_sc_hd__buf_2_5_X ;
wire [0:0] sky130_fd_sc_hd__buf_2_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_10_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_11_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_12_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_13_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_14_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_12_X[0] ) , .X ( lut3_out[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_1_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_13_X[0] ) , .X ( lut3_out[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_2_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_14_X[0] ) , .X ( lut4_out[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_3_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .X ( sky130_fd_sc_hd__buf_2_3_X[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_4_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , 
    .X ( sky130_fd_sc_hd__buf_2_4_X[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_5_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_10_X[0] ) , 
    .X ( sky130_fd_sc_hd__buf_2_5_X[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_6_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_11_X[0] ) , 
    .X ( sky130_fd_sc_hd__buf_2_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_3_ ( .A0 ( in[7] ) , .A1 ( in[6] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_4_ ( .A0 ( in[9] ) , .A1 ( in[8] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_5_ ( .A0 ( in[11] ) , .A1 ( in[10] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_6_ ( .A0 ( in[13] ) , .A1 ( in[12] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_7_ ( .A0 ( in[15] ) , .A1 ( in[14] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_10_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_11_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( .A0 ( sky130_fd_sc_hd__buf_2_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__buf_2_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_12_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( .A0 ( sky130_fd_sc_hd__buf_2_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__buf_2_5_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_13_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_13_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_12_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_14_X[0] ) ) ;
endmodule


module frac_lut4_2 ( in , sram , sram_inv , mode , mode_inv , lut3_out , 
    lut4_out ) ;
input  [0:3] in ;
input  [0:15] sram ;
input  [0:15] sram_inv ;
input  [0:0] mode ;
input  [0:0] mode_inv ;
output [0:1] lut3_out ;
output [0:0] lut4_out ;

wire [0:0] sky130_fd_sc_hd__buf_2_0_X ;
wire [0:0] sky130_fd_sc_hd__buf_2_1_X ;
wire [0:0] sky130_fd_sc_hd__buf_2_2_X ;
wire [0:0] sky130_fd_sc_hd__buf_2_3_X ;
wire [0:0] sky130_fd_sc_hd__inv_1_0_Y ;
wire [0:0] sky130_fd_sc_hd__inv_1_1_Y ;
wire [0:0] sky130_fd_sc_hd__inv_1_2_Y ;
wire [0:0] sky130_fd_sc_hd__inv_1_3_Y ;
wire [0:0] sky130_fd_sc_hd__or2_1_0_X ;

sky130_fd_sc_hd__or2_0 sky130_fd_sc_hd__or2_1_0_ ( .A ( mode[0] ) , 
    .B ( in[3] ) , .X ( sky130_fd_sc_hd__or2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__inv_1 sky130_fd_sc_hd__inv_1_0_ ( .A ( in[0] ) , 
    .Y ( sky130_fd_sc_hd__inv_1_0_Y[0] ) ) ;
sky130_fd_sc_hd__inv_1 sky130_fd_sc_hd__inv_1_1_ ( .A ( in[1] ) , 
    .Y ( sky130_fd_sc_hd__inv_1_1_Y[0] ) ) ;
sky130_fd_sc_hd__inv_1 sky130_fd_sc_hd__inv_1_2_ ( .A ( in[2] ) , 
    .Y ( sky130_fd_sc_hd__inv_1_2_Y[0] ) ) ;
sky130_fd_sc_hd__inv_1 sky130_fd_sc_hd__inv_1_3_ ( 
    .A ( sky130_fd_sc_hd__or2_1_0_X[0] ) , 
    .Y ( sky130_fd_sc_hd__inv_1_3_Y[0] ) ) ;
sky130_fd_sc_hd__buf_2 sky130_fd_sc_hd__buf_2_0_ ( .A ( in[0] ) , 
    .X ( sky130_fd_sc_hd__buf_2_0_X[0] ) ) ;
sky130_fd_sc_hd__buf_2 sky130_fd_sc_hd__buf_2_1_ ( .A ( in[1] ) , 
    .X ( sky130_fd_sc_hd__buf_2_1_X[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_2_ ( .A ( in[2] ) , 
    .X ( sky130_fd_sc_hd__buf_2_2_X[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_3_ ( 
    .A ( sky130_fd_sc_hd__or2_1_0_X[0] ) , 
    .X ( sky130_fd_sc_hd__buf_2_3_X[0] ) ) ;
frac_lut4_mux_2 frac_lut4_mux_0_ ( .in ( sram ) ,
    .sram ( { sky130_fd_sc_hd__buf_2_0_X[0] , sky130_fd_sc_hd__buf_2_1_X[0] , 
        sky130_fd_sc_hd__buf_2_2_X[0] , sky130_fd_sc_hd__buf_2_3_X[0] } ) ,
    .sram_inv ( { sky130_fd_sc_hd__inv_1_0_Y[0] , 
        sky130_fd_sc_hd__inv_1_1_Y[0] , sky130_fd_sc_hd__inv_1_2_Y[0] , 
        sky130_fd_sc_hd__inv_1_3_Y[0] } ) ,
    .lut3_out ( lut3_out ) , .lut4_out ( lut4_out ) ) ;
endmodule


module logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_2 ( 
    prog_clk , frac_lut4_in , ccff_head , frac_lut4_lut3_out , 
    frac_lut4_lut4_out , ccff_tail ) ;
input  [0:0] prog_clk ;
input  [0:3] frac_lut4_in ;
input  [0:0] ccff_head ;
output [0:1] frac_lut4_lut3_out ;
output [0:0] frac_lut4_lut4_out ;
output [0:0] ccff_tail ;

wire [0:0] frac_lut4_0_mode ;
wire [0:15] frac_lut4_0_sram ;
wire [0:15] frac_lut4_0_sram_inv ;

frac_lut4_2 frac_lut4_0_ ( .in ( frac_lut4_in ) , .sram ( frac_lut4_0_sram ) , 
    .sram_inv ( frac_lut4_0_sram_inv ) , .mode ( frac_lut4_0_mode ) ,
    .mode_inv ( { SYNOPSYS_UNCONNECTED_1 } ) ,
    .lut3_out ( frac_lut4_lut3_out ) , .lut4_out ( frac_lut4_lut4_out ) ) ;
frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem_2 frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem ( 
    .prog_clk ( prog_clk ) , .ccff_head ( ccff_head ) , 
    .ccff_tail ( ccff_tail ) ,
    .mem_out ( { frac_lut4_0_sram[0] , frac_lut4_0_sram[1] , 
        frac_lut4_0_sram[2] , frac_lut4_0_sram[3] , frac_lut4_0_sram[4] , 
        frac_lut4_0_sram[5] , frac_lut4_0_sram[6] , frac_lut4_0_sram[7] , 
        frac_lut4_0_sram[8] , frac_lut4_0_sram[9] , frac_lut4_0_sram[10] , 
        frac_lut4_0_sram[11] , frac_lut4_0_sram[12] , frac_lut4_0_sram[13] , 
        frac_lut4_0_sram[14] , frac_lut4_0_sram[15] , frac_lut4_0_mode[0] } ) ,
    .mem_outb ( { frac_lut4_0_sram_inv[0] , frac_lut4_0_sram_inv[1] , 
        frac_lut4_0_sram_inv[2] , frac_lut4_0_sram_inv[3] , 
        frac_lut4_0_sram_inv[4] , frac_lut4_0_sram_inv[5] , 
        frac_lut4_0_sram_inv[6] , frac_lut4_0_sram_inv[7] , 
        frac_lut4_0_sram_inv[8] , frac_lut4_0_sram_inv[9] , 
        frac_lut4_0_sram_inv[10] , frac_lut4_0_sram_inv[11] , 
        frac_lut4_0_sram_inv[12] , frac_lut4_0_sram_inv[13] , 
        frac_lut4_0_sram_inv[14] , frac_lut4_0_sram_inv[15] , 
        SYNOPSYS_UNCONNECTED_2 } ) ) ;
endmodule


module logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_2 ( 
    prog_clk , frac_logic_in , ccff_head , frac_logic_out , ccff_tail , p0 ) ;
input  [0:0] prog_clk ;
input  [0:3] frac_logic_in ;
input  [0:0] ccff_head ;
output [0:1] frac_logic_out ;
output [0:0] ccff_tail ;
input  p0 ;

wire [0:0] logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_ccff_tail ;
wire [0:0] logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_frac_lut4_lut3_out ;
wire [0:0] logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_frac_lut4_lut4_out ;
wire [0:1] mux_tree_size2_0_sram ;
wire [0:1] mux_tree_size2_0_sram_inv ;

logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_2 logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0 ( 
    .prog_clk ( prog_clk ) , .frac_lut4_in ( frac_logic_in ) , 
    .ccff_head ( ccff_head ) ,
    .frac_lut4_lut3_out ( { 
        logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_frac_lut4_lut3_out[0] , 
        frac_logic_out[1] } ) ,
    
    .frac_lut4_lut4_out ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_frac_lut4_lut4_out ) , 
    .ccff_tail ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_ccff_tail ) ) ;
mux_tree_size2_26 mux_frac_logic_out_0 (
    .in ( { 
        logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_frac_lut4_lut4_out[0] , 
        logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_frac_lut4_lut3_out[0]
         } ) ,
    .sram ( mux_tree_size2_0_sram ) , 
    .sram_inv ( mux_tree_size2_0_sram_inv ) , .out ( frac_logic_out[0] ) , 
    .p0 ( p0 ) ) ;
mux_tree_size2_mem_26 mem_frac_logic_out_0 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_ccff_tail ) , 
    .ccff_tail ( ccff_tail ) , .mem_out ( mux_tree_size2_0_sram ) , 
    .mem_outb ( mux_tree_size2_0_sram_inv ) ) ;
direct_interc direct_interc_0_ (
    .in ( { SYNOPSYS_UNCONNECTED_1 } ) ,
    .out ( frac_logic_out[1] ) ) ;
direct_interc direct_interc_1_ (
    .in ( { SYNOPSYS_UNCONNECTED_2 } ) ,
    .out ( frac_logic_in[0] ) ) ;
direct_interc direct_interc_2_ (
    .in ( { SYNOPSYS_UNCONNECTED_3 } ) ,
    .out ( frac_logic_in[1] ) ) ;
direct_interc direct_interc_3_ (
    .in ( { SYNOPSYS_UNCONNECTED_4 } ) ,
    .out ( frac_logic_in[2] ) ) ;
direct_interc direct_interc_4_ (
    .in ( { SYNOPSYS_UNCONNECTED_5 } ) ,
    .out ( frac_logic_in[3] ) ) ;
endmodule


module logical_tile_clb_mode_default__fle_mode_physical__fabric_2 ( prog_clk , 
    Test_en , clk , fabric_in , fabric_regin , fabric_scin , fabric_clk , 
    ccff_head , fabric_out , fabric_regout , fabric_scout , ccff_tail , p0 ) ;
input  [0:0] prog_clk ;
input  [0:0] Test_en ;
input  [0:0] clk ;
input  [0:3] fabric_in ;
input  [0:0] fabric_regin ;
input  [0:0] fabric_scin ;
input  [0:0] fabric_clk ;
input  [0:0] ccff_head ;
output [0:1] fabric_out ;
output [0:0] fabric_regout ;
output [0:0] fabric_scout ;
output [0:0] ccff_tail ;
input  p0 ;

wire [0:0] logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0_ff_Q ;
wire [0:0] logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_ccff_tail ;
wire [0:1] logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_frac_logic_out ;
wire [0:1] mux_tree_size2_0_sram ;
wire [0:1] mux_tree_size2_0_sram_inv ;
wire [0:1] mux_tree_size2_1_sram ;
wire [0:1] mux_tree_size2_1_sram_inv ;
wire [0:0] mux_tree_size2_2_out ;
wire [0:1] mux_tree_size2_2_sram ;
wire [0:1] mux_tree_size2_2_sram_inv ;
wire [0:0] mux_tree_size2_mem_0_ccff_tail ;
wire [0:0] mux_tree_size2_mem_1_ccff_tail ;

assign fabric_regout[0] = fabric_scout[0] ;

logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_2 logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0 ( 
    .prog_clk ( prog_clk ) , .frac_logic_in ( fabric_in ) , 
    .ccff_head ( ccff_head ) , 
    .frac_logic_out ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_frac_logic_out ) , 
    .ccff_tail ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_ccff_tail ) , 
    .p0 ( p0 ) ) ;
logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_4 logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0 ( 
    .Test_en ( Test_en ) , .clk ( clk ) , .ff_D ( mux_tree_size2_2_out ) , 
    .ff_DI ( fabric_scin ) , 
    .ff_Q ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0_ff_Q ) ,
    .ff_clk ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_5 logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1 ( 
    .Test_en ( Test_en ) , .clk ( clk ) , 
    .ff_D ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_frac_logic_out[1] ) , 
    .ff_DI ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0_ff_Q ) , 
    .ff_Q ( fabric_scout ) ,
    .ff_clk ( { SYNOPSYS_UNCONNECTED_2 } ) ) ;
mux_tree_size2_6 mux_fabric_out_0 (
    .in ( { 
        logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0_ff_Q[0] , 
        logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_frac_logic_out[0]
         } ) ,
    .sram ( mux_tree_size2_0_sram ) , 
    .sram_inv ( mux_tree_size2_0_sram_inv ) , .out ( fabric_out[0] ) , 
    .p0 ( p0 ) ) ;
mux_tree_size2_7 mux_fabric_out_1 (
    .in ( { fabric_scout[0] , 
        logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_frac_logic_out[1]
         } ) ,
    .sram ( mux_tree_size2_1_sram ) , 
    .sram_inv ( mux_tree_size2_1_sram_inv ) , .out ( fabric_out[1] ) , 
    .p0 ( p0 ) ) ;
mux_tree_size2_8 mux_ff_0_D_0 (
    .in ( { 
        logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_frac_logic_out[0] , 
        fabric_regin[0] } ) ,
    .sram ( mux_tree_size2_2_sram ) , 
    .sram_inv ( mux_tree_size2_2_sram_inv ) , .out ( mux_tree_size2_2_out ) , 
    .p0 ( p0 ) ) ;
mux_tree_size2_mem_6 mem_fabric_out_0 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_size2_mem_0_ccff_tail ) , 
    .mem_out ( mux_tree_size2_0_sram ) , 
    .mem_outb ( mux_tree_size2_0_sram_inv ) ) ;
mux_tree_size2_mem_7 mem_fabric_out_1 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_size2_mem_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_size2_mem_1_ccff_tail ) , 
    .mem_out ( mux_tree_size2_1_sram ) , 
    .mem_outb ( mux_tree_size2_1_sram_inv ) ) ;
mux_tree_size2_mem_8 mem_ff_0_D_0 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_size2_mem_1_ccff_tail ) , .ccff_tail ( ccff_tail ) , 
    .mem_out ( mux_tree_size2_2_sram ) , 
    .mem_outb ( mux_tree_size2_2_sram_inv ) ) ;
direct_interc direct_interc_0_ (
    .in ( { SYNOPSYS_UNCONNECTED_3 } ) ,
    .out ( fabric_scout ) ) ;
direct_interc direct_interc_1_ (
    .in ( { SYNOPSYS_UNCONNECTED_4 } ) ,
    .out ( fabric_scout ) ) ;
direct_interc direct_interc_2_ (
    .in ( { SYNOPSYS_UNCONNECTED_5 } ) ,
    .out ( fabric_in[0] ) ) ;
direct_interc direct_interc_3_ (
    .in ( { SYNOPSYS_UNCONNECTED_6 } ) ,
    .out ( fabric_in[1] ) ) ;
direct_interc direct_interc_4_ (
    .in ( { SYNOPSYS_UNCONNECTED_7 } ) ,
    .out ( fabric_in[2] ) ) ;
direct_interc direct_interc_5_ (
    .in ( { SYNOPSYS_UNCONNECTED_8 } ) ,
    .out ( fabric_in[3] ) ) ;
direct_interc direct_interc_6_ (
    .in ( { SYNOPSYS_UNCONNECTED_9 } ) ,
    .out ( fabric_scin ) ) ;
direct_interc direct_interc_7_ (
    .in ( { SYNOPSYS_UNCONNECTED_10 } ) ,
    .out ( fabric_clk ) ) ;
direct_interc direct_interc_8_ (
    .in ( { SYNOPSYS_UNCONNECTED_11 } ) ,
    
    .out ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_frac_logic_out[1] ) ) ;
direct_interc direct_interc_9_ (
    .in ( { SYNOPSYS_UNCONNECTED_12 } ) ,
    
    .out ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0_ff_Q ) ) ;
direct_interc direct_interc_10_ (
    .in ( { SYNOPSYS_UNCONNECTED_13 } ) ,
    .out ( fabric_clk ) ) ;
endmodule


module logical_tile_clb_mode_default__fle_2 ( prog_clk , Test_en , clk , 
    fle_in , fle_regin , fle_scin , fle_clk , ccff_head , fle_out , 
    fle_regout , fle_scout , ccff_tail , p0 ) ;
input  [0:0] prog_clk ;
input  [0:0] Test_en ;
input  [0:0] clk ;
input  [0:3] fle_in ;
input  [0:0] fle_regin ;
input  [0:0] fle_scin ;
input  [0:0] fle_clk ;
input  [0:0] ccff_head ;
output [0:1] fle_out ;
output [0:0] fle_regout ;
output [0:0] fle_scout ;
output [0:0] ccff_tail ;
input  p0 ;

logical_tile_clb_mode_default__fle_mode_physical__fabric_2 logical_tile_clb_mode_default__fle_mode_physical__fabric_0 ( 
    .prog_clk ( prog_clk ) , .Test_en ( Test_en ) , .clk ( clk ) , 
    .fabric_in ( fle_in ) , .fabric_regin ( fle_regin ) , 
    .fabric_scin ( fle_scin ) , .fabric_clk ( fle_clk ) , 
    .ccff_head ( ccff_head ) , .fabric_out ( fle_out ) , 
    .fabric_regout ( fle_regout ) , .fabric_scout ( fle_scout ) , 
    .ccff_tail ( ccff_tail ) , .p0 ( p0 ) ) ;
direct_interc direct_interc_0_ (
    .in ( { SYNOPSYS_UNCONNECTED_1 } ) ,
    .out ( fle_out[0] ) ) ;
direct_interc direct_interc_1_ (
    .in ( { SYNOPSYS_UNCONNECTED_2 } ) ,
    .out ( fle_out[1] ) ) ;
direct_interc direct_interc_2_ (
    .in ( { SYNOPSYS_UNCONNECTED_3 } ) ,
    .out ( fle_regout ) ) ;
direct_interc direct_interc_3_ (
    .in ( { SYNOPSYS_UNCONNECTED_4 } ) ,
    .out ( fle_scout ) ) ;
direct_interc direct_interc_4_ (
    .in ( { SYNOPSYS_UNCONNECTED_5 } ) ,
    .out ( fle_in[0] ) ) ;
direct_interc direct_interc_5_ (
    .in ( { SYNOPSYS_UNCONNECTED_6 } ) ,
    .out ( fle_in[1] ) ) ;
direct_interc direct_interc_6_ (
    .in ( { SYNOPSYS_UNCONNECTED_7 } ) ,
    .out ( fle_in[2] ) ) ;
direct_interc direct_interc_7_ (
    .in ( { SYNOPSYS_UNCONNECTED_8 } ) ,
    .out ( fle_in[3] ) ) ;
direct_interc direct_interc_8_ (
    .in ( { SYNOPSYS_UNCONNECTED_9 } ) ,
    .out ( fle_regin ) ) ;
direct_interc direct_interc_9_ (
    .in ( { SYNOPSYS_UNCONNECTED_10 } ) ,
    .out ( fle_scin ) ) ;
direct_interc direct_interc_10_ (
    .in ( { SYNOPSYS_UNCONNECTED_11 } ) ,
    .out ( fle_clk ) ) ;
endmodule


module mux_tree_size2_mem_5 ( prog_clk , ccff_head , ccff_tail , mem_out , 
    mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_10__25 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_size2_mem_4 ( prog_clk , ccff_head , ccff_tail , mem_out , 
    mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_9__24 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_size2_mem_3 ( prog_clk , ccff_head , ccff_tail , mem_out , 
    mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_8__23 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_7 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_size2_5 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;

const1_7 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , .X ( out[0] ) ) ;
endmodule


module const1_6 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_size2_4 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;

const1_6 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , .X ( out[0] ) ) ;
endmodule


module const1_5 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_size2_3 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;

const1_5 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , .X ( out[0] ) ) ;
endmodule


module logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_3 ( 
    Test_en , clk , ff_D , ff_DI , ff_Q , ff_clk ) ;
input  [0:0] Test_en ;
input  [0:0] clk ;
input  [0:0] ff_D ;
input  [0:0] ff_DI ;
output [0:0] ff_Q ;
input  [0:0] ff_clk ;

sky130_fd_sc_hd__sdfxbp_1 sky130_fd_sc_hd__sdfxbp_1_0_ ( .D ( ff_D[0] ) , 
    .SCD ( ff_DI[0] ) , .SCE ( Test_en[0] ) , .CLK ( clk[0] ) , 
    .Q ( ff_Q[0] ) , .Q_N ( SYNOPSYS_UNCONNECTED_1 ) ) ;
endmodule


module logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_2 ( 
    Test_en , clk , ff_D , ff_DI , ff_Q , ff_clk ) ;
input  [0:0] Test_en ;
input  [0:0] clk ;
input  [0:0] ff_D ;
input  [0:0] ff_DI ;
output [0:0] ff_Q ;
input  [0:0] ff_clk ;

sky130_fd_sc_hd__sdfxbp_1 sky130_fd_sc_hd__sdfxbp_1_0_ ( .D ( ff_D[0] ) , 
    .SCD ( ff_DI[0] ) , .SCE ( Test_en[0] ) , .CLK ( clk[0] ) , 
    .Q ( ff_Q[0] ) , .Q_N ( SYNOPSYS_UNCONNECTED_1 ) ) ;
endmodule


module mux_tree_size2_mem_25 ( prog_clk , ccff_head , ccff_tail , mem_out , 
    mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_7__22 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_4 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_size2_25 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;

const1_4 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , .X ( out[0] ) ) ;
endmodule


module frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem_1 ( prog_clk , ccff_head , 
    ccff_tail , mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:16] mem_out ;
output [0:16] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_4_ ( .D ( mem_out[3] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[4] ) , .Q_N ( mem_outb[4] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_5_ ( .D ( mem_out[4] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[5] ) , .Q_N ( mem_outb[5] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_6_ ( .D ( mem_out[5] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[6] ) , .Q_N ( mem_outb[6] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_7_ ( .D ( mem_out[6] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[7] ) , .Q_N ( mem_outb[7] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_8_ ( .D ( mem_out[7] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[8] ) , .Q_N ( mem_outb[8] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_9_ ( .D ( mem_out[8] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[9] ) , .Q_N ( mem_outb[9] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_10_ ( .D ( mem_out[9] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[10] ) , .Q_N ( mem_outb[10] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_11_ ( .D ( mem_out[10] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[11] ) , .Q_N ( mem_outb[11] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_12_ ( .D ( mem_out[11] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[12] ) , .Q_N ( mem_outb[12] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_13_ ( .D ( mem_out[12] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[13] ) , .Q_N ( mem_outb[13] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_14_ ( .D ( mem_out[13] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[14] ) , .Q_N ( mem_outb[14] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_15_ ( .D ( mem_out[14] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[15] ) , .Q_N ( mem_outb[15] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_16_ ( .D ( mem_out[15] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[16] ) , .Q_N ( \_gOb1_mem_outb[16] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_6__21 ( .A ( mem_out[16] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module frac_lut4_mux_1 ( in , sram , sram_inv , lut3_out , lut4_out ) ;
input  [0:15] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:1] lut3_out ;
output [0:0] lut4_out ;

wire [0:0] sky130_fd_sc_hd__buf_2_3_X ;
wire [0:0] sky130_fd_sc_hd__buf_2_4_X ;
wire [0:0] sky130_fd_sc_hd__buf_2_5_X ;
wire [0:0] sky130_fd_sc_hd__buf_2_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_10_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_11_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_12_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_13_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_14_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_12_X[0] ) , .X ( lut3_out[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_1_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_13_X[0] ) , .X ( lut3_out[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_2_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_14_X[0] ) , .X ( lut4_out[0] ) ) ;
sky130_fd_sc_hd__buf_2 sky130_fd_sc_hd__buf_2_3_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .X ( sky130_fd_sc_hd__buf_2_3_X[0] ) ) ;
sky130_fd_sc_hd__buf_2 sky130_fd_sc_hd__buf_2_4_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , 
    .X ( sky130_fd_sc_hd__buf_2_4_X[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_5_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_10_X[0] ) , 
    .X ( sky130_fd_sc_hd__buf_2_5_X[0] ) ) ;
sky130_fd_sc_hd__buf_2 sky130_fd_sc_hd__buf_2_6_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_11_X[0] ) , 
    .X ( sky130_fd_sc_hd__buf_2_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_3_ ( .A0 ( in[7] ) , .A1 ( in[6] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_4_ ( .A0 ( in[9] ) , .A1 ( in[8] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_5_ ( .A0 ( in[11] ) , .A1 ( in[10] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_6_ ( .A0 ( in[13] ) , .A1 ( in[12] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_7_ ( .A0 ( in[15] ) , .A1 ( in[14] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_10_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_11_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( .A0 ( sky130_fd_sc_hd__buf_2_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__buf_2_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_12_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( .A0 ( sky130_fd_sc_hd__buf_2_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__buf_2_5_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_13_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_13_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_12_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_14_X[0] ) ) ;
endmodule


module frac_lut4_1 ( in , sram , sram_inv , mode , mode_inv , lut3_out , 
    lut4_out ) ;
input  [0:3] in ;
input  [0:15] sram ;
input  [0:15] sram_inv ;
input  [0:0] mode ;
input  [0:0] mode_inv ;
output [0:1] lut3_out ;
output [0:0] lut4_out ;

wire [0:0] sky130_fd_sc_hd__buf_2_0_X ;
wire [0:0] sky130_fd_sc_hd__buf_2_1_X ;
wire [0:0] sky130_fd_sc_hd__buf_2_2_X ;
wire [0:0] sky130_fd_sc_hd__buf_2_3_X ;
wire [0:0] sky130_fd_sc_hd__inv_1_0_Y ;
wire [0:0] sky130_fd_sc_hd__inv_1_1_Y ;
wire [0:0] sky130_fd_sc_hd__inv_1_2_Y ;
wire [0:0] sky130_fd_sc_hd__inv_1_3_Y ;
wire [0:0] sky130_fd_sc_hd__or2_1_0_X ;

sky130_fd_sc_hd__or2_0 sky130_fd_sc_hd__or2_1_0_ ( .A ( mode[0] ) , 
    .B ( in[3] ) , .X ( sky130_fd_sc_hd__or2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__inv_1 sky130_fd_sc_hd__inv_1_0_ ( .A ( in[0] ) , 
    .Y ( sky130_fd_sc_hd__inv_1_0_Y[0] ) ) ;
sky130_fd_sc_hd__inv_1 sky130_fd_sc_hd__inv_1_1_ ( .A ( in[1] ) , 
    .Y ( sky130_fd_sc_hd__inv_1_1_Y[0] ) ) ;
sky130_fd_sc_hd__inv_1 sky130_fd_sc_hd__inv_1_2_ ( .A ( in[2] ) , 
    .Y ( sky130_fd_sc_hd__inv_1_2_Y[0] ) ) ;
sky130_fd_sc_hd__inv_1 sky130_fd_sc_hd__inv_1_3_ ( 
    .A ( sky130_fd_sc_hd__or2_1_0_X[0] ) , 
    .Y ( sky130_fd_sc_hd__inv_1_3_Y[0] ) ) ;
sky130_fd_sc_hd__buf_2 sky130_fd_sc_hd__buf_2_0_ ( .A ( in[0] ) , 
    .X ( sky130_fd_sc_hd__buf_2_0_X[0] ) ) ;
sky130_fd_sc_hd__buf_2 sky130_fd_sc_hd__buf_2_1_ ( .A ( in[1] ) , 
    .X ( sky130_fd_sc_hd__buf_2_1_X[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_2_ ( .A ( in[2] ) , 
    .X ( sky130_fd_sc_hd__buf_2_2_X[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_3_ ( 
    .A ( sky130_fd_sc_hd__or2_1_0_X[0] ) , 
    .X ( sky130_fd_sc_hd__buf_2_3_X[0] ) ) ;
frac_lut4_mux_1 frac_lut4_mux_0_ ( .in ( sram ) ,
    .sram ( { sky130_fd_sc_hd__buf_2_0_X[0] , sky130_fd_sc_hd__buf_2_1_X[0] , 
        sky130_fd_sc_hd__buf_2_2_X[0] , sky130_fd_sc_hd__buf_2_3_X[0] } ) ,
    .sram_inv ( { sky130_fd_sc_hd__inv_1_0_Y[0] , 
        sky130_fd_sc_hd__inv_1_1_Y[0] , sky130_fd_sc_hd__inv_1_2_Y[0] , 
        sky130_fd_sc_hd__inv_1_3_Y[0] } ) ,
    .lut3_out ( lut3_out ) , .lut4_out ( lut4_out ) ) ;
endmodule


module logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_1 ( 
    prog_clk , frac_lut4_in , ccff_head , frac_lut4_lut3_out , 
    frac_lut4_lut4_out , ccff_tail ) ;
input  [0:0] prog_clk ;
input  [0:3] frac_lut4_in ;
input  [0:0] ccff_head ;
output [0:1] frac_lut4_lut3_out ;
output [0:0] frac_lut4_lut4_out ;
output [0:0] ccff_tail ;

wire [0:0] frac_lut4_0_mode ;
wire [0:15] frac_lut4_0_sram ;
wire [0:15] frac_lut4_0_sram_inv ;

frac_lut4_1 frac_lut4_0_ ( .in ( frac_lut4_in ) , .sram ( frac_lut4_0_sram ) , 
    .sram_inv ( frac_lut4_0_sram_inv ) , .mode ( frac_lut4_0_mode ) ,
    .mode_inv ( { SYNOPSYS_UNCONNECTED_1 } ) ,
    .lut3_out ( frac_lut4_lut3_out ) , .lut4_out ( frac_lut4_lut4_out ) ) ;
frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem_1 frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem ( 
    .prog_clk ( prog_clk ) , .ccff_head ( ccff_head ) , 
    .ccff_tail ( ccff_tail ) ,
    .mem_out ( { frac_lut4_0_sram[0] , frac_lut4_0_sram[1] , 
        frac_lut4_0_sram[2] , frac_lut4_0_sram[3] , frac_lut4_0_sram[4] , 
        frac_lut4_0_sram[5] , frac_lut4_0_sram[6] , frac_lut4_0_sram[7] , 
        frac_lut4_0_sram[8] , frac_lut4_0_sram[9] , frac_lut4_0_sram[10] , 
        frac_lut4_0_sram[11] , frac_lut4_0_sram[12] , frac_lut4_0_sram[13] , 
        frac_lut4_0_sram[14] , frac_lut4_0_sram[15] , frac_lut4_0_mode[0] } ) ,
    .mem_outb ( { frac_lut4_0_sram_inv[0] , frac_lut4_0_sram_inv[1] , 
        frac_lut4_0_sram_inv[2] , frac_lut4_0_sram_inv[3] , 
        frac_lut4_0_sram_inv[4] , frac_lut4_0_sram_inv[5] , 
        frac_lut4_0_sram_inv[6] , frac_lut4_0_sram_inv[7] , 
        frac_lut4_0_sram_inv[8] , frac_lut4_0_sram_inv[9] , 
        frac_lut4_0_sram_inv[10] , frac_lut4_0_sram_inv[11] , 
        frac_lut4_0_sram_inv[12] , frac_lut4_0_sram_inv[13] , 
        frac_lut4_0_sram_inv[14] , frac_lut4_0_sram_inv[15] , 
        SYNOPSYS_UNCONNECTED_2 } ) ) ;
endmodule


module logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_1 ( 
    prog_clk , frac_logic_in , ccff_head , frac_logic_out , ccff_tail , p0 ) ;
input  [0:0] prog_clk ;
input  [0:3] frac_logic_in ;
input  [0:0] ccff_head ;
output [0:1] frac_logic_out ;
output [0:0] ccff_tail ;
input  p0 ;

wire [0:0] logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_ccff_tail ;
wire [0:0] logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_frac_lut4_lut3_out ;
wire [0:0] logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_frac_lut4_lut4_out ;
wire [0:1] mux_tree_size2_0_sram ;
wire [0:1] mux_tree_size2_0_sram_inv ;

logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_1 logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0 ( 
    .prog_clk ( prog_clk ) , .frac_lut4_in ( frac_logic_in ) , 
    .ccff_head ( ccff_head ) ,
    .frac_lut4_lut3_out ( { 
        logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_frac_lut4_lut3_out[0] , 
        frac_logic_out[1] } ) ,
    
    .frac_lut4_lut4_out ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_frac_lut4_lut4_out ) , 
    .ccff_tail ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_ccff_tail ) ) ;
mux_tree_size2_25 mux_frac_logic_out_0 (
    .in ( { 
        logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_frac_lut4_lut4_out[0] , 
        logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_frac_lut4_lut3_out[0]
         } ) ,
    .sram ( mux_tree_size2_0_sram ) , 
    .sram_inv ( mux_tree_size2_0_sram_inv ) , .out ( frac_logic_out[0] ) , 
    .p0 ( p0 ) ) ;
mux_tree_size2_mem_25 mem_frac_logic_out_0 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_ccff_tail ) , 
    .ccff_tail ( ccff_tail ) , .mem_out ( mux_tree_size2_0_sram ) , 
    .mem_outb ( mux_tree_size2_0_sram_inv ) ) ;
direct_interc direct_interc_0_ (
    .in ( { SYNOPSYS_UNCONNECTED_1 } ) ,
    .out ( frac_logic_out[1] ) ) ;
direct_interc direct_interc_1_ (
    .in ( { SYNOPSYS_UNCONNECTED_2 } ) ,
    .out ( frac_logic_in[0] ) ) ;
direct_interc direct_interc_2_ (
    .in ( { SYNOPSYS_UNCONNECTED_3 } ) ,
    .out ( frac_logic_in[1] ) ) ;
direct_interc direct_interc_3_ (
    .in ( { SYNOPSYS_UNCONNECTED_4 } ) ,
    .out ( frac_logic_in[2] ) ) ;
direct_interc direct_interc_4_ (
    .in ( { SYNOPSYS_UNCONNECTED_5 } ) ,
    .out ( frac_logic_in[3] ) ) ;
endmodule


module logical_tile_clb_mode_default__fle_mode_physical__fabric_1 ( prog_clk , 
    Test_en , clk , fabric_in , fabric_regin , fabric_scin , fabric_clk , 
    ccff_head , fabric_out , fabric_regout , fabric_scout , ccff_tail , p0 , 
    p1 ) ;
input  [0:0] prog_clk ;
input  [0:0] Test_en ;
input  [0:0] clk ;
input  [0:3] fabric_in ;
input  [0:0] fabric_regin ;
input  [0:0] fabric_scin ;
input  [0:0] fabric_clk ;
input  [0:0] ccff_head ;
output [0:1] fabric_out ;
output [0:0] fabric_regout ;
output [0:0] fabric_scout ;
output [0:0] ccff_tail ;
input  p0 ;
input  p1 ;

wire [0:0] logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0_ff_Q ;
wire [0:0] logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_ccff_tail ;
wire [0:1] logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_frac_logic_out ;
wire [0:1] mux_tree_size2_0_sram ;
wire [0:1] mux_tree_size2_0_sram_inv ;
wire [0:1] mux_tree_size2_1_sram ;
wire [0:1] mux_tree_size2_1_sram_inv ;
wire [0:0] mux_tree_size2_2_out ;
wire [0:1] mux_tree_size2_2_sram ;
wire [0:1] mux_tree_size2_2_sram_inv ;
wire [0:0] mux_tree_size2_mem_0_ccff_tail ;
wire [0:0] mux_tree_size2_mem_1_ccff_tail ;

assign fabric_regout[0] = fabric_scout[0] ;

logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_1 logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0 ( 
    .prog_clk ( prog_clk ) , .frac_logic_in ( fabric_in ) , 
    .ccff_head ( ccff_head ) , 
    .frac_logic_out ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_frac_logic_out ) , 
    .ccff_tail ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_ccff_tail ) , 
    .p0 ( p0 ) ) ;
logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_2 logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0 ( 
    .Test_en ( Test_en ) , .clk ( clk ) , .ff_D ( mux_tree_size2_2_out ) , 
    .ff_DI ( fabric_scin ) , 
    .ff_Q ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0_ff_Q ) ,
    .ff_clk ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_3 logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1 ( 
    .Test_en ( Test_en ) , .clk ( clk ) , 
    .ff_D ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_frac_logic_out[1] ) , 
    .ff_DI ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0_ff_Q ) , 
    .ff_Q ( fabric_scout ) ,
    .ff_clk ( { SYNOPSYS_UNCONNECTED_2 } ) ) ;
mux_tree_size2_3 mux_fabric_out_0 (
    .in ( { 
        logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0_ff_Q[0] , 
        logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_frac_logic_out[0]
         } ) ,
    .sram ( mux_tree_size2_0_sram ) , 
    .sram_inv ( mux_tree_size2_0_sram_inv ) , .out ( fabric_out[0] ) , 
    .p0 ( p0 ) ) ;
mux_tree_size2_4 mux_fabric_out_1 (
    .in ( { fabric_scout[0] , 
        logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_frac_logic_out[1]
         } ) ,
    .sram ( mux_tree_size2_1_sram ) , 
    .sram_inv ( mux_tree_size2_1_sram_inv ) , .out ( fabric_out[1] ) , 
    .p0 ( p0 ) ) ;
mux_tree_size2_5 mux_ff_0_D_0 (
    .in ( { 
        logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_frac_logic_out[0] , 
        fabric_regin[0] } ) ,
    .sram ( mux_tree_size2_2_sram ) , 
    .sram_inv ( mux_tree_size2_2_sram_inv ) , .out ( mux_tree_size2_2_out ) , 
    .p0 ( p1 ) ) ;
mux_tree_size2_mem_3 mem_fabric_out_0 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_size2_mem_0_ccff_tail ) , 
    .mem_out ( mux_tree_size2_0_sram ) , 
    .mem_outb ( mux_tree_size2_0_sram_inv ) ) ;
mux_tree_size2_mem_4 mem_fabric_out_1 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_size2_mem_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_size2_mem_1_ccff_tail ) , 
    .mem_out ( mux_tree_size2_1_sram ) , 
    .mem_outb ( mux_tree_size2_1_sram_inv ) ) ;
mux_tree_size2_mem_5 mem_ff_0_D_0 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_size2_mem_1_ccff_tail ) , .ccff_tail ( ccff_tail ) , 
    .mem_out ( mux_tree_size2_2_sram ) , 
    .mem_outb ( mux_tree_size2_2_sram_inv ) ) ;
direct_interc direct_interc_0_ (
    .in ( { SYNOPSYS_UNCONNECTED_3 } ) ,
    .out ( fabric_scout ) ) ;
direct_interc direct_interc_1_ (
    .in ( { SYNOPSYS_UNCONNECTED_4 } ) ,
    .out ( fabric_scout ) ) ;
direct_interc direct_interc_2_ (
    .in ( { SYNOPSYS_UNCONNECTED_5 } ) ,
    .out ( fabric_in[0] ) ) ;
direct_interc direct_interc_3_ (
    .in ( { SYNOPSYS_UNCONNECTED_6 } ) ,
    .out ( fabric_in[1] ) ) ;
direct_interc direct_interc_4_ (
    .in ( { SYNOPSYS_UNCONNECTED_7 } ) ,
    .out ( fabric_in[2] ) ) ;
direct_interc direct_interc_5_ (
    .in ( { SYNOPSYS_UNCONNECTED_8 } ) ,
    .out ( fabric_in[3] ) ) ;
direct_interc direct_interc_6_ (
    .in ( { SYNOPSYS_UNCONNECTED_9 } ) ,
    .out ( fabric_scin ) ) ;
direct_interc direct_interc_7_ (
    .in ( { SYNOPSYS_UNCONNECTED_10 } ) ,
    .out ( fabric_clk ) ) ;
direct_interc direct_interc_8_ (
    .in ( { SYNOPSYS_UNCONNECTED_11 } ) ,
    
    .out ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_frac_logic_out[1] ) ) ;
direct_interc direct_interc_9_ (
    .in ( { SYNOPSYS_UNCONNECTED_12 } ) ,
    
    .out ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0_ff_Q ) ) ;
direct_interc direct_interc_10_ (
    .in ( { SYNOPSYS_UNCONNECTED_13 } ) ,
    .out ( fabric_clk ) ) ;
endmodule


module logical_tile_clb_mode_default__fle_1 ( prog_clk , Test_en , clk , 
    fle_in , fle_regin , fle_scin , fle_clk , ccff_head , fle_out , 
    fle_regout , fle_scout , ccff_tail , p0 , p1 ) ;
input  [0:0] prog_clk ;
input  [0:0] Test_en ;
input  [0:0] clk ;
input  [0:3] fle_in ;
input  [0:0] fle_regin ;
input  [0:0] fle_scin ;
input  [0:0] fle_clk ;
input  [0:0] ccff_head ;
output [0:1] fle_out ;
output [0:0] fle_regout ;
output [0:0] fle_scout ;
output [0:0] ccff_tail ;
input  p0 ;
input  p1 ;

logical_tile_clb_mode_default__fle_mode_physical__fabric_1 logical_tile_clb_mode_default__fle_mode_physical__fabric_0 ( 
    .prog_clk ( prog_clk ) , .Test_en ( Test_en ) , .clk ( clk ) , 
    .fabric_in ( fle_in ) , .fabric_regin ( fle_regin ) , 
    .fabric_scin ( fle_scin ) , .fabric_clk ( fle_clk ) , 
    .ccff_head ( ccff_head ) , .fabric_out ( fle_out ) , 
    .fabric_regout ( fle_regout ) , .fabric_scout ( fle_scout ) , 
    .ccff_tail ( ccff_tail ) , .p0 ( p0 ) , .p1 ( p1 ) ) ;
direct_interc direct_interc_0_ (
    .in ( { SYNOPSYS_UNCONNECTED_1 } ) ,
    .out ( fle_out[0] ) ) ;
direct_interc direct_interc_1_ (
    .in ( { SYNOPSYS_UNCONNECTED_2 } ) ,
    .out ( fle_out[1] ) ) ;
direct_interc direct_interc_2_ (
    .in ( { SYNOPSYS_UNCONNECTED_3 } ) ,
    .out ( fle_regout ) ) ;
direct_interc direct_interc_3_ (
    .in ( { SYNOPSYS_UNCONNECTED_4 } ) ,
    .out ( fle_scout ) ) ;
direct_interc direct_interc_4_ (
    .in ( { SYNOPSYS_UNCONNECTED_5 } ) ,
    .out ( fle_in[0] ) ) ;
direct_interc direct_interc_5_ (
    .in ( { SYNOPSYS_UNCONNECTED_6 } ) ,
    .out ( fle_in[1] ) ) ;
direct_interc direct_interc_6_ (
    .in ( { SYNOPSYS_UNCONNECTED_7 } ) ,
    .out ( fle_in[2] ) ) ;
direct_interc direct_interc_7_ (
    .in ( { SYNOPSYS_UNCONNECTED_8 } ) ,
    .out ( fle_in[3] ) ) ;
direct_interc direct_interc_8_ (
    .in ( { SYNOPSYS_UNCONNECTED_9 } ) ,
    .out ( fle_regin ) ) ;
direct_interc direct_interc_9_ (
    .in ( { SYNOPSYS_UNCONNECTED_10 } ) ,
    .out ( fle_scin ) ) ;
direct_interc direct_interc_10_ (
    .in ( { SYNOPSYS_UNCONNECTED_11 } ) ,
    .out ( fle_clk ) ) ;
endmodule


module mux_tree_size2_mem_2 ( prog_clk , ccff_head , ccff_tail , mem_out , 
    mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_5__20 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_size2_mem_1 ( prog_clk , ccff_head , ccff_tail , mem_out , 
    mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_4__19 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module mux_tree_size2_mem_0 ( prog_clk , ccff_head , ccff_tail , mem_out , 
    mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_3__18 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_3 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_size2_2 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;

const1_3 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , .X ( out[0] ) ) ;
endmodule


module const1_2 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_size2_1 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;

const1_2 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , .X ( out[0] ) ) ;
endmodule


module const1_1 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_size2_0 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;

const1_1 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , .X ( out[0] ) ) ;
endmodule


module logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1 ( 
    Test_en , clk , ff_D , ff_DI , ff_Q , ff_clk ) ;
input  [0:0] Test_en ;
input  [0:0] clk ;
input  [0:0] ff_D ;
input  [0:0] ff_DI ;
output [0:0] ff_Q ;
input  [0:0] ff_clk ;

sky130_fd_sc_hd__sdfxbp_1 sky130_fd_sc_hd__sdfxbp_1_0_ ( .D ( ff_D[0] ) , 
    .SCD ( ff_DI[0] ) , .SCE ( Test_en[0] ) , .CLK ( clk[0] ) , 
    .Q ( ff_Q[0] ) , .Q_N ( SYNOPSYS_UNCONNECTED_1 ) ) ;
endmodule


module logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0 ( 
    Test_en , clk , ff_D , ff_DI , ff_Q , ff_clk ) ;
input  [0:0] Test_en ;
input  [0:0] clk ;
input  [0:0] ff_D ;
input  [0:0] ff_DI ;
output [0:0] ff_Q ;
input  [0:0] ff_clk ;

sky130_fd_sc_hd__sdfxbp_1 sky130_fd_sc_hd__sdfxbp_1_0_ ( .D ( ff_D[0] ) , 
    .SCD ( ff_DI[0] ) , .SCE ( Test_en[0] ) , .CLK ( clk[0] ) , 
    .Q ( ff_Q[0] ) , .Q_N ( SYNOPSYS_UNCONNECTED_1 ) ) ;
endmodule


module direct_interc ( in , out ) ;
input  [0:0] in ;
output [0:0] out ;

assign out[0] = in[0] ;
endmodule


module mux_tree_size2_mem_24 ( prog_clk , ccff_head , ccff_tail , mem_out , 
    mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:1] mem_out ;
output [0:1] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_2__17 ( .A ( mem_out[1] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module const1_0 ( const1 ) ;
output [0:0] const1 ;
endmodule


module mux_tree_size2_24 ( in , sram , sram_inv , out , p0 ) ;
input  [0:1] in ;
input  [0:1] sram ;
input  [0:1] sram_inv ;
output [0:0] out ;
input  p0 ;

wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;

const1_0 const1_0_ (
    .const1 ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( .A0 ( p0 ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , .X ( out[0] ) ) ;
endmodule


module frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem_0 ( prog_clk , ccff_head , 
    ccff_tail , mem_out , mem_outb ) ;
input  [0:0] prog_clk ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;
output [0:16] mem_out ;
output [0:16] mem_outb ;

sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_0_ ( .D ( ccff_head[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[0] ) , .Q_N ( mem_outb[0] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_1_ ( .D ( mem_out[0] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[1] ) , .Q_N ( mem_outb[1] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_2_ ( .D ( mem_out[1] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[2] ) , .Q_N ( mem_outb[2] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_3_ ( .D ( mem_out[2] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[3] ) , .Q_N ( mem_outb[3] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_4_ ( .D ( mem_out[3] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[4] ) , .Q_N ( mem_outb[4] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_5_ ( .D ( mem_out[4] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[5] ) , .Q_N ( mem_outb[5] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_6_ ( .D ( mem_out[5] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[6] ) , .Q_N ( mem_outb[6] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_7_ ( .D ( mem_out[6] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[7] ) , .Q_N ( mem_outb[7] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_8_ ( .D ( mem_out[7] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[8] ) , .Q_N ( mem_outb[8] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_9_ ( .D ( mem_out[8] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[9] ) , .Q_N ( mem_outb[9] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_10_ ( .D ( mem_out[9] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[10] ) , .Q_N ( mem_outb[10] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_11_ ( .D ( mem_out[10] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[11] ) , .Q_N ( mem_outb[11] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_12_ ( .D ( mem_out[11] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[12] ) , .Q_N ( mem_outb[12] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_13_ ( .D ( mem_out[12] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[13] ) , .Q_N ( mem_outb[13] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_14_ ( .D ( mem_out[13] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[14] ) , .Q_N ( mem_outb[14] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_15_ ( .D ( mem_out[14] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[15] ) , .Q_N ( mem_outb[15] ) ) ;
sky130_fd_sc_hd__dfxbp_1 sky130_fd_sc_hd__dfxbp_1_16_ ( .D ( mem_out[15] ) , 
    .CLK ( prog_clk[0] ) , .Q ( mem_out[16] ) , .Q_N ( \_gOb0_mem_outb[16] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_1__16 ( .A ( mem_out[16] ) , 
    .X ( ccff_tail[0] ) ) ;
endmodule


module frac_lut4_mux_0 ( in , sram , sram_inv , lut3_out , lut4_out ) ;
input  [0:15] in ;
input  [0:3] sram ;
input  [0:3] sram_inv ;
output [0:1] lut3_out ;
output [0:0] lut4_out ;

wire [0:0] sky130_fd_sc_hd__buf_2_3_X ;
wire [0:0] sky130_fd_sc_hd__buf_2_4_X ;
wire [0:0] sky130_fd_sc_hd__buf_2_5_X ;
wire [0:0] sky130_fd_sc_hd__buf_2_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_0_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_10_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_11_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_12_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_13_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_14_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_1_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_2_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_3_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_4_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_5_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_6_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_7_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_8_X ;
wire [0:0] sky130_fd_sc_hd__mux2_1_9_X ;

sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_0_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_12_X[0] ) , .X ( lut3_out[0] ) ) ;
sky130_fd_sc_hd__buf_2 sky130_fd_sc_hd__buf_2_1_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_13_X[0] ) , .X ( lut3_out[1] ) ) ;
sky130_fd_sc_hd__buf_2 sky130_fd_sc_hd__buf_2_2_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_14_X[0] ) , .X ( lut4_out[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_3_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_8_X[0] ) , 
    .X ( sky130_fd_sc_hd__buf_2_3_X[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_4_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_9_X[0] ) , 
    .X ( sky130_fd_sc_hd__buf_2_4_X[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_5_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_10_X[0] ) , 
    .X ( sky130_fd_sc_hd__buf_2_5_X[0] ) ) ;
sky130_fd_sc_hd__buf_2 sky130_fd_sc_hd__buf_2_6_ ( 
    .A ( sky130_fd_sc_hd__mux2_1_11_X[0] ) , 
    .X ( sky130_fd_sc_hd__buf_2_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_0_ ( .A0 ( in[1] ) , .A1 ( in[0] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_1_ ( .A0 ( in[3] ) , .A1 ( in[2] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_1_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_2_ ( .A0 ( in[5] ) , .A1 ( in[4] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_2_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_3_ ( .A0 ( in[7] ) , .A1 ( in[6] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_3_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_4_ ( .A0 ( in[9] ) , .A1 ( in[8] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_4_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_5_ ( .A0 ( in[11] ) , .A1 ( in[10] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_5_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_6_ ( .A0 ( in[13] ) , .A1 ( in[12] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_6_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l1_in_7_ ( .A0 ( in[15] ) , .A1 ( in[14] ) , 
    .S ( sram[0] ) , .X ( sky130_fd_sc_hd__mux2_1_7_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_1_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_0_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_8_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_1_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_3_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_2_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_9_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_2_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_5_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_4_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_10_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l2_in_3_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_7_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_6_X[0] ) , .S ( sram[1] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_11_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_0_ ( .A0 ( sky130_fd_sc_hd__buf_2_4_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__buf_2_3_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_12_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l3_in_1_ ( .A0 ( sky130_fd_sc_hd__buf_2_6_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__buf_2_5_X[0] ) , .S ( sram[2] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_13_X[0] ) ) ;
sky130_fd_sc_hd__mux2_1 mux_l4_in_0_ ( 
    .A0 ( sky130_fd_sc_hd__mux2_1_13_X[0] ) , 
    .A1 ( sky130_fd_sc_hd__mux2_1_12_X[0] ) , .S ( sram[3] ) , 
    .X ( sky130_fd_sc_hd__mux2_1_14_X[0] ) ) ;
endmodule


module frac_lut4_0 ( in , sram , sram_inv , mode , mode_inv , lut3_out , 
    lut4_out ) ;
input  [0:3] in ;
input  [0:15] sram ;
input  [0:15] sram_inv ;
input  [0:0] mode ;
input  [0:0] mode_inv ;
output [0:1] lut3_out ;
output [0:0] lut4_out ;

wire [0:0] sky130_fd_sc_hd__buf_2_0_X ;
wire [0:0] sky130_fd_sc_hd__buf_2_1_X ;
wire [0:0] sky130_fd_sc_hd__buf_2_2_X ;
wire [0:0] sky130_fd_sc_hd__buf_2_3_X ;
wire [0:0] sky130_fd_sc_hd__inv_1_0_Y ;
wire [0:0] sky130_fd_sc_hd__inv_1_1_Y ;
wire [0:0] sky130_fd_sc_hd__inv_1_2_Y ;
wire [0:0] sky130_fd_sc_hd__inv_1_3_Y ;
wire [0:0] sky130_fd_sc_hd__or2_1_0_X ;

sky130_fd_sc_hd__or2_0 sky130_fd_sc_hd__or2_1_0_ ( .A ( mode[0] ) , 
    .B ( in[3] ) , .X ( sky130_fd_sc_hd__or2_1_0_X[0] ) ) ;
sky130_fd_sc_hd__inv_1 sky130_fd_sc_hd__inv_1_0_ ( .A ( in[0] ) , 
    .Y ( sky130_fd_sc_hd__inv_1_0_Y[0] ) ) ;
sky130_fd_sc_hd__inv_1 sky130_fd_sc_hd__inv_1_1_ ( .A ( in[1] ) , 
    .Y ( sky130_fd_sc_hd__inv_1_1_Y[0] ) ) ;
sky130_fd_sc_hd__inv_1 sky130_fd_sc_hd__inv_1_2_ ( .A ( in[2] ) , 
    .Y ( sky130_fd_sc_hd__inv_1_2_Y[0] ) ) ;
sky130_fd_sc_hd__inv_1 sky130_fd_sc_hd__inv_1_3_ ( 
    .A ( sky130_fd_sc_hd__or2_1_0_X[0] ) , 
    .Y ( sky130_fd_sc_hd__inv_1_3_Y[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_0_ ( .A ( in[0] ) , 
    .X ( sky130_fd_sc_hd__buf_2_0_X[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_1_ ( .A ( in[1] ) , 
    .X ( sky130_fd_sc_hd__buf_2_1_X[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 sky130_fd_sc_hd__buf_2_2_ ( .A ( in[2] ) , 
    .X ( sky130_fd_sc_hd__buf_2_2_X[0] ) ) ;
sky130_fd_sc_hd__buf_2 sky130_fd_sc_hd__buf_2_3_ ( 
    .A ( sky130_fd_sc_hd__or2_1_0_X[0] ) , 
    .X ( sky130_fd_sc_hd__buf_2_3_X[0] ) ) ;
frac_lut4_mux_0 frac_lut4_mux_0_ ( .in ( sram ) ,
    .sram ( { sky130_fd_sc_hd__buf_2_0_X[0] , sky130_fd_sc_hd__buf_2_1_X[0] , 
        sky130_fd_sc_hd__buf_2_2_X[0] , sky130_fd_sc_hd__buf_2_3_X[0] } ) ,
    .sram_inv ( { sky130_fd_sc_hd__inv_1_0_Y[0] , 
        sky130_fd_sc_hd__inv_1_1_Y[0] , sky130_fd_sc_hd__inv_1_2_Y[0] , 
        sky130_fd_sc_hd__inv_1_3_Y[0] } ) ,
    .lut3_out ( lut3_out ) , .lut4_out ( lut4_out ) ) ;
endmodule


module logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0 ( 
    prog_clk , frac_lut4_in , ccff_head , frac_lut4_lut3_out , 
    frac_lut4_lut4_out , ccff_tail ) ;
input  [0:0] prog_clk ;
input  [0:3] frac_lut4_in ;
input  [0:0] ccff_head ;
output [0:1] frac_lut4_lut3_out ;
output [0:0] frac_lut4_lut4_out ;
output [0:0] ccff_tail ;

wire [0:0] frac_lut4_0_mode ;
wire [0:15] frac_lut4_0_sram ;
wire [0:15] frac_lut4_0_sram_inv ;

frac_lut4_0 frac_lut4_0_ ( .in ( frac_lut4_in ) , .sram ( frac_lut4_0_sram ) , 
    .sram_inv ( frac_lut4_0_sram_inv ) , .mode ( frac_lut4_0_mode ) ,
    .mode_inv ( { SYNOPSYS_UNCONNECTED_1 } ) ,
    .lut3_out ( frac_lut4_lut3_out ) , .lut4_out ( frac_lut4_lut4_out ) ) ;
frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem_0 frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem ( 
    .prog_clk ( prog_clk ) , .ccff_head ( ccff_head ) , 
    .ccff_tail ( ccff_tail ) ,
    .mem_out ( { frac_lut4_0_sram[0] , frac_lut4_0_sram[1] , 
        frac_lut4_0_sram[2] , frac_lut4_0_sram[3] , frac_lut4_0_sram[4] , 
        frac_lut4_0_sram[5] , frac_lut4_0_sram[6] , frac_lut4_0_sram[7] , 
        frac_lut4_0_sram[8] , frac_lut4_0_sram[9] , frac_lut4_0_sram[10] , 
        frac_lut4_0_sram[11] , frac_lut4_0_sram[12] , frac_lut4_0_sram[13] , 
        frac_lut4_0_sram[14] , frac_lut4_0_sram[15] , frac_lut4_0_mode[0] } ) ,
    .mem_outb ( { frac_lut4_0_sram_inv[0] , frac_lut4_0_sram_inv[1] , 
        frac_lut4_0_sram_inv[2] , frac_lut4_0_sram_inv[3] , 
        frac_lut4_0_sram_inv[4] , frac_lut4_0_sram_inv[5] , 
        frac_lut4_0_sram_inv[6] , frac_lut4_0_sram_inv[7] , 
        frac_lut4_0_sram_inv[8] , frac_lut4_0_sram_inv[9] , 
        frac_lut4_0_sram_inv[10] , frac_lut4_0_sram_inv[11] , 
        frac_lut4_0_sram_inv[12] , frac_lut4_0_sram_inv[13] , 
        frac_lut4_0_sram_inv[14] , frac_lut4_0_sram_inv[15] , 
        SYNOPSYS_UNCONNECTED_2 } ) ) ;
endmodule


module logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0 ( 
    prog_clk , frac_logic_in , ccff_head , frac_logic_out , ccff_tail , p0 ) ;
input  [0:0] prog_clk ;
input  [0:3] frac_logic_in ;
input  [0:0] ccff_head ;
output [0:1] frac_logic_out ;
output [0:0] ccff_tail ;
input  p0 ;

wire [0:0] logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_ccff_tail ;
wire [0:0] logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_frac_lut4_lut3_out ;
wire [0:0] logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_frac_lut4_lut4_out ;
wire [0:1] mux_tree_size2_0_sram ;
wire [0:1] mux_tree_size2_0_sram_inv ;

logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0 logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0 ( 
    .prog_clk ( prog_clk ) , .frac_lut4_in ( frac_logic_in ) , 
    .ccff_head ( ccff_head ) ,
    .frac_lut4_lut3_out ( { 
        logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_frac_lut4_lut3_out[0] , 
        frac_logic_out[1] } ) ,
    
    .frac_lut4_lut4_out ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_frac_lut4_lut4_out ) , 
    .ccff_tail ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_ccff_tail ) ) ;
mux_tree_size2_24 mux_frac_logic_out_0 (
    .in ( { 
        logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_frac_lut4_lut4_out[0] , 
        logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_frac_lut4_lut3_out[0]
         } ) ,
    .sram ( mux_tree_size2_0_sram ) , 
    .sram_inv ( mux_tree_size2_0_sram_inv ) , .out ( frac_logic_out[0] ) , 
    .p0 ( p0 ) ) ;
mux_tree_size2_mem_24 mem_frac_logic_out_0 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0_ccff_tail ) , 
    .ccff_tail ( ccff_tail ) , .mem_out ( mux_tree_size2_0_sram ) , 
    .mem_outb ( mux_tree_size2_0_sram_inv ) ) ;
direct_interc direct_interc_0_ (
    .in ( { SYNOPSYS_UNCONNECTED_1 } ) ,
    .out ( frac_logic_out[1] ) ) ;
direct_interc direct_interc_1_ (
    .in ( { SYNOPSYS_UNCONNECTED_2 } ) ,
    .out ( frac_logic_in[0] ) ) ;
direct_interc direct_interc_2_ (
    .in ( { SYNOPSYS_UNCONNECTED_3 } ) ,
    .out ( frac_logic_in[1] ) ) ;
direct_interc direct_interc_3_ (
    .in ( { SYNOPSYS_UNCONNECTED_4 } ) ,
    .out ( frac_logic_in[2] ) ) ;
direct_interc direct_interc_4_ (
    .in ( { SYNOPSYS_UNCONNECTED_5 } ) ,
    .out ( frac_logic_in[3] ) ) ;
endmodule


module logical_tile_clb_mode_default__fle_mode_physical__fabric_0 ( prog_clk , 
    Test_en , clk , fabric_in , fabric_regin , fabric_scin , fabric_clk , 
    ccff_head , fabric_out , fabric_regout , fabric_scout , ccff_tail , p1 ) ;
input  [0:0] prog_clk ;
input  [0:0] Test_en ;
input  [0:0] clk ;
input  [0:3] fabric_in ;
input  [0:0] fabric_regin ;
input  [0:0] fabric_scin ;
input  [0:0] fabric_clk ;
input  [0:0] ccff_head ;
output [0:1] fabric_out ;
output [0:0] fabric_regout ;
output [0:0] fabric_scout ;
output [0:0] ccff_tail ;
input  p1 ;

wire [0:0] logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0_ff_Q ;
wire [0:0] logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_ccff_tail ;
wire [0:1] logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_frac_logic_out ;
wire [0:1] mux_tree_size2_0_sram ;
wire [0:1] mux_tree_size2_0_sram_inv ;
wire [0:1] mux_tree_size2_1_sram ;
wire [0:1] mux_tree_size2_1_sram_inv ;
wire [0:0] mux_tree_size2_2_out ;
wire [0:1] mux_tree_size2_2_sram ;
wire [0:1] mux_tree_size2_2_sram_inv ;
wire [0:0] mux_tree_size2_mem_0_ccff_tail ;
wire [0:0] mux_tree_size2_mem_1_ccff_tail ;

assign fabric_regout[0] = fabric_scout[0] ;

logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0 logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0 ( 
    .prog_clk ( prog_clk ) , .frac_logic_in ( fabric_in ) , 
    .ccff_head ( ccff_head ) , 
    .frac_logic_out ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_frac_logic_out ) , 
    .ccff_tail ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_ccff_tail ) , 
    .p0 ( p1 ) ) ;
logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0 logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0 ( 
    .Test_en ( Test_en ) , .clk ( clk ) , .ff_D ( mux_tree_size2_2_out ) , 
    .ff_DI ( fabric_scin ) , 
    .ff_Q ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0_ff_Q ) ,
    .ff_clk ( { SYNOPSYS_UNCONNECTED_1 } ) ) ;
logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1 logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1 ( 
    .Test_en ( Test_en ) , .clk ( clk ) , 
    .ff_D ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_frac_logic_out[1] ) , 
    .ff_DI ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0_ff_Q ) , 
    .ff_Q ( fabric_scout ) ,
    .ff_clk ( { SYNOPSYS_UNCONNECTED_2 } ) ) ;
mux_tree_size2_0 mux_fabric_out_0 (
    .in ( { 
        logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0_ff_Q[0] , 
        logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_frac_logic_out[0]
         } ) ,
    .sram ( mux_tree_size2_0_sram ) , 
    .sram_inv ( mux_tree_size2_0_sram_inv ) , .out ( fabric_out[0] ) , 
    .p0 ( p1 ) ) ;
mux_tree_size2_1 mux_fabric_out_1 (
    .in ( { fabric_scout[0] , 
        logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_frac_logic_out[1]
         } ) ,
    .sram ( mux_tree_size2_1_sram ) , 
    .sram_inv ( mux_tree_size2_1_sram_inv ) , .out ( fabric_out[1] ) , 
    .p0 ( p1 ) ) ;
mux_tree_size2_2 mux_ff_0_D_0 (
    .in ( { 
        logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_frac_logic_out[0] , 
        fabric_regin[0] } ) ,
    .sram ( mux_tree_size2_2_sram ) , 
    .sram_inv ( mux_tree_size2_2_sram_inv ) , .out ( mux_tree_size2_2_out ) , 
    .p0 ( p1 ) ) ;
mux_tree_size2_mem_0 mem_fabric_out_0 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_size2_mem_0_ccff_tail ) , 
    .mem_out ( mux_tree_size2_0_sram ) , 
    .mem_outb ( mux_tree_size2_0_sram_inv ) ) ;
mux_tree_size2_mem_1 mem_fabric_out_1 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_size2_mem_0_ccff_tail ) , 
    .ccff_tail ( mux_tree_size2_mem_1_ccff_tail ) , 
    .mem_out ( mux_tree_size2_1_sram ) , 
    .mem_outb ( mux_tree_size2_1_sram_inv ) ) ;
mux_tree_size2_mem_2 mem_ff_0_D_0 ( .prog_clk ( prog_clk ) , 
    .ccff_head ( mux_tree_size2_mem_1_ccff_tail ) , .ccff_tail ( ccff_tail ) , 
    .mem_out ( mux_tree_size2_2_sram ) , 
    .mem_outb ( mux_tree_size2_2_sram_inv ) ) ;
direct_interc direct_interc_0_ (
    .in ( { SYNOPSYS_UNCONNECTED_3 } ) ,
    .out ( fabric_scout ) ) ;
direct_interc direct_interc_1_ (
    .in ( { SYNOPSYS_UNCONNECTED_4 } ) ,
    .out ( fabric_scout ) ) ;
direct_interc direct_interc_2_ (
    .in ( { SYNOPSYS_UNCONNECTED_5 } ) ,
    .out ( fabric_in[0] ) ) ;
direct_interc direct_interc_3_ (
    .in ( { SYNOPSYS_UNCONNECTED_6 } ) ,
    .out ( fabric_in[1] ) ) ;
direct_interc direct_interc_4_ (
    .in ( { SYNOPSYS_UNCONNECTED_7 } ) ,
    .out ( fabric_in[2] ) ) ;
direct_interc direct_interc_5_ (
    .in ( { SYNOPSYS_UNCONNECTED_8 } ) ,
    .out ( fabric_in[3] ) ) ;
direct_interc direct_interc_6_ (
    .in ( { SYNOPSYS_UNCONNECTED_9 } ) ,
    .out ( fabric_scin ) ) ;
direct_interc direct_interc_7_ (
    .in ( { SYNOPSYS_UNCONNECTED_10 } ) ,
    .out ( fabric_clk ) ) ;
direct_interc direct_interc_8_ (
    .in ( { SYNOPSYS_UNCONNECTED_11 } ) ,
    
    .out ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0_frac_logic_out[1] ) ) ;
direct_interc direct_interc_9_ (
    .in ( { SYNOPSYS_UNCONNECTED_12 } ) ,
    
    .out ( logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0_ff_Q ) ) ;
direct_interc direct_interc_10_ (
    .in ( { SYNOPSYS_UNCONNECTED_13 } ) ,
    .out ( fabric_clk ) ) ;
endmodule


module logical_tile_clb_mode_default__fle_0 ( prog_clk , Test_en , clk , 
    fle_in , fle_regin , fle_scin , fle_clk , ccff_head , fle_out , 
    fle_regout , fle_scout , ccff_tail , p1 ) ;
input  [0:0] prog_clk ;
input  [0:0] Test_en ;
input  [0:0] clk ;
input  [0:3] fle_in ;
input  [0:0] fle_regin ;
input  [0:0] fle_scin ;
input  [0:0] fle_clk ;
input  [0:0] ccff_head ;
output [0:1] fle_out ;
output [0:0] fle_regout ;
output [0:0] fle_scout ;
output [0:0] ccff_tail ;
input  p1 ;

logical_tile_clb_mode_default__fle_mode_physical__fabric_0 logical_tile_clb_mode_default__fle_mode_physical__fabric_0 ( 
    .prog_clk ( prog_clk ) , .Test_en ( Test_en ) , .clk ( clk ) , 
    .fabric_in ( fle_in ) , .fabric_regin ( fle_regin ) , 
    .fabric_scin ( fle_scin ) , .fabric_clk ( fle_clk ) , 
    .ccff_head ( ccff_head ) , .fabric_out ( fle_out ) , 
    .fabric_regout ( fle_regout ) , .fabric_scout ( fle_scout ) , 
    .ccff_tail ( ccff_tail ) , .p1 ( p1 ) ) ;
direct_interc direct_interc_0_ (
    .in ( { SYNOPSYS_UNCONNECTED_1 } ) ,
    .out ( fle_out[0] ) ) ;
direct_interc direct_interc_1_ (
    .in ( { SYNOPSYS_UNCONNECTED_2 } ) ,
    .out ( fle_out[1] ) ) ;
direct_interc direct_interc_2_ (
    .in ( { SYNOPSYS_UNCONNECTED_3 } ) ,
    .out ( fle_regout ) ) ;
direct_interc direct_interc_3_ (
    .in ( { SYNOPSYS_UNCONNECTED_4 } ) ,
    .out ( fle_scout ) ) ;
direct_interc direct_interc_4_ (
    .in ( { SYNOPSYS_UNCONNECTED_5 } ) ,
    .out ( fle_in[0] ) ) ;
direct_interc direct_interc_5_ (
    .in ( { SYNOPSYS_UNCONNECTED_6 } ) ,
    .out ( fle_in[1] ) ) ;
direct_interc direct_interc_6_ (
    .in ( { SYNOPSYS_UNCONNECTED_7 } ) ,
    .out ( fle_in[2] ) ) ;
direct_interc direct_interc_7_ (
    .in ( { SYNOPSYS_UNCONNECTED_8 } ) ,
    .out ( fle_in[3] ) ) ;
direct_interc direct_interc_8_ (
    .in ( { SYNOPSYS_UNCONNECTED_9 } ) ,
    .out ( fle_regin ) ) ;
direct_interc direct_interc_9_ (
    .in ( { SYNOPSYS_UNCONNECTED_10 } ) ,
    .out ( fle_scin ) ) ;
direct_interc direct_interc_10_ (
    .in ( { SYNOPSYS_UNCONNECTED_11 } ) ,
    .out ( fle_clk ) ) ;
endmodule


module logical_tile_clb_mode_clb_ ( prog_clk , Test_en , clk , clb_I0 , 
    clb_I1 , clb_I2 , clb_I3 , clb_I4 , clb_I5 , clb_I6 , clb_I7 , clb_regin , 
    clb_scin , clb_clk , ccff_head , clb_O , clb_regout , clb_scout , 
    ccff_tail , p_abuf0 , p_abuf1 , p_abuf2 , p_abuf3 , p_abuf4 , p_abuf5 , 
    p_abuf6 , p_abuf7 , p_abuf8 , p_abuf9 , p_abuf10 , p_abuf11 , p_abuf12 , 
    p_abuf13 , p_abuf14 , p_abuf15 , p0 , p1 , p2 , p3 , p4 ) ;
input  [0:0] prog_clk ;
input  [0:0] Test_en ;
input  [0:0] clk ;
input  [0:3] clb_I0 ;
input  [0:3] clb_I1 ;
input  [0:3] clb_I2 ;
input  [0:3] clb_I3 ;
input  [0:3] clb_I4 ;
input  [0:3] clb_I5 ;
input  [0:3] clb_I6 ;
input  [0:3] clb_I7 ;
input  [0:0] clb_regin ;
input  [0:0] clb_scin ;
input  [0:0] clb_clk ;
input  [0:0] ccff_head ;
output [0:15] clb_O ;
output [0:0] clb_regout ;
output [0:0] clb_scout ;
output [0:0] ccff_tail ;
output p_abuf0 ;
output p_abuf1 ;
output p_abuf2 ;
output p_abuf3 ;
output p_abuf4 ;
output p_abuf5 ;
output p_abuf6 ;
output p_abuf7 ;
output p_abuf8 ;
output p_abuf9 ;
output p_abuf10 ;
output p_abuf11 ;
output p_abuf12 ;
output p_abuf13 ;
output p_abuf14 ;
output p_abuf15 ;
input  p0 ;
input  p1 ;
input  p2 ;
input  p3 ;
input  p4 ;

wire [0:0] logical_tile_clb_mode_default__fle_0_ccff_tail ;
wire [1:1] logical_tile_clb_mode_default__fle_0_fle_out ;
wire [0:0] logical_tile_clb_mode_default__fle_0_fle_regout ;
wire [0:0] logical_tile_clb_mode_default__fle_0_fle_scout ;
wire [0:0] logical_tile_clb_mode_default__fle_1_ccff_tail ;
wire [1:1] logical_tile_clb_mode_default__fle_1_fle_out ;
wire [0:0] logical_tile_clb_mode_default__fle_1_fle_regout ;
wire [0:0] logical_tile_clb_mode_default__fle_1_fle_scout ;
wire [0:0] logical_tile_clb_mode_default__fle_2_ccff_tail ;
wire [0:0] logical_tile_clb_mode_default__fle_2_fle_regout ;
wire [0:0] logical_tile_clb_mode_default__fle_2_fle_scout ;
wire [0:0] logical_tile_clb_mode_default__fle_3_ccff_tail ;
wire [0:1] logical_tile_clb_mode_default__fle_3_fle_out ;
wire [0:0] logical_tile_clb_mode_default__fle_3_fle_regout ;
wire [0:0] logical_tile_clb_mode_default__fle_3_fle_scout ;
wire [0:0] logical_tile_clb_mode_default__fle_4_ccff_tail ;
wire [1:1] logical_tile_clb_mode_default__fle_4_fle_out ;
wire [0:0] logical_tile_clb_mode_default__fle_4_fle_regout ;
wire [0:0] logical_tile_clb_mode_default__fle_4_fle_scout ;
wire [0:0] logical_tile_clb_mode_default__fle_5_ccff_tail ;
wire [0:0] logical_tile_clb_mode_default__fle_5_fle_out ;
wire [0:0] logical_tile_clb_mode_default__fle_5_fle_regout ;
wire [0:0] logical_tile_clb_mode_default__fle_5_fle_scout ;
wire [0:0] logical_tile_clb_mode_default__fle_6_ccff_tail ;
wire [0:0] logical_tile_clb_mode_default__fle_6_fle_out ;
wire [0:0] logical_tile_clb_mode_default__fle_6_fle_regout ;
wire [0:0] logical_tile_clb_mode_default__fle_6_fle_scout ;

logical_tile_clb_mode_default__fle_0 logical_tile_clb_mode_default__fle_0 ( 
    .prog_clk ( prog_clk ) , .Test_en ( Test_en ) , .clk ( clk ) , 
    .fle_in ( clb_I0 ) , .fle_regin ( clb_regin ) , .fle_scin ( clb_scin ) , 
    .fle_clk ( clb_clk ) , .ccff_head ( ccff_head ) ,
    .fle_out ( { clb_O[1] , logical_tile_clb_mode_default__fle_0_fle_out[1] } ) ,
    .fle_regout ( logical_tile_clb_mode_default__fle_0_fle_regout ) , 
    .fle_scout ( logical_tile_clb_mode_default__fle_0_fle_scout ) , 
    .ccff_tail ( logical_tile_clb_mode_default__fle_0_ccff_tail ) , 
    .p1 ( p1 ) ) ;
logical_tile_clb_mode_default__fle_1 logical_tile_clb_mode_default__fle_1 ( 
    .prog_clk ( prog_clk ) , .Test_en ( Test_en ) , .clk ( clk ) , 
    .fle_in ( clb_I1 ) , 
    .fle_regin ( logical_tile_clb_mode_default__fle_0_fle_regout ) , 
    .fle_scin ( logical_tile_clb_mode_default__fle_0_fle_scout ) , 
    .fle_clk ( clb_clk ) , 
    .ccff_head ( logical_tile_clb_mode_default__fle_0_ccff_tail ) ,
    .fle_out ( { clb_O[3] , logical_tile_clb_mode_default__fle_1_fle_out[1] } ) ,
    .fle_regout ( logical_tile_clb_mode_default__fle_1_fle_regout ) , 
    .fle_scout ( logical_tile_clb_mode_default__fle_1_fle_scout ) , 
    .ccff_tail ( logical_tile_clb_mode_default__fle_1_ccff_tail ) , 
    .p0 ( p0 ) , .p1 ( p1 ) ) ;
logical_tile_clb_mode_default__fle_2 logical_tile_clb_mode_default__fle_2 ( 
    .prog_clk ( prog_clk ) , .Test_en ( Test_en ) , .clk ( clk ) , 
    .fle_in ( clb_I2 ) , 
    .fle_regin ( logical_tile_clb_mode_default__fle_1_fle_regout ) , 
    .fle_scin ( logical_tile_clb_mode_default__fle_1_fle_scout ) , 
    .fle_clk ( clb_clk ) , 
    .ccff_head ( logical_tile_clb_mode_default__fle_1_ccff_tail ) ,
    .fle_out ( { clb_O[5] , clb_O[4] } ) ,
    .fle_regout ( logical_tile_clb_mode_default__fle_2_fle_regout ) , 
    .fle_scout ( logical_tile_clb_mode_default__fle_2_fle_scout ) , 
    .ccff_tail ( logical_tile_clb_mode_default__fle_2_ccff_tail ) , 
    .p0 ( p0 ) ) ;
logical_tile_clb_mode_default__fle_3 logical_tile_clb_mode_default__fle_3 ( 
    .prog_clk ( prog_clk ) , .Test_en ( Test_en ) , .clk ( clk ) , 
    .fle_in ( clb_I3 ) , 
    .fle_regin ( logical_tile_clb_mode_default__fle_2_fle_regout ) , 
    .fle_scin ( logical_tile_clb_mode_default__fle_2_fle_scout ) , 
    .fle_clk ( clb_clk ) , 
    .ccff_head ( logical_tile_clb_mode_default__fle_2_ccff_tail ) , 
    .fle_out ( logical_tile_clb_mode_default__fle_3_fle_out ) , 
    .fle_regout ( logical_tile_clb_mode_default__fle_3_fle_regout ) , 
    .fle_scout ( logical_tile_clb_mode_default__fle_3_fle_scout ) , 
    .ccff_tail ( logical_tile_clb_mode_default__fle_3_ccff_tail ) , 
    .p0 ( p0 ) , .p3 ( p4 ) ) ;
logical_tile_clb_mode_default__fle_4 logical_tile_clb_mode_default__fle_4 ( 
    .prog_clk ( prog_clk ) , .Test_en ( Test_en ) , .clk ( clk ) , 
    .fle_in ( clb_I4 ) , 
    .fle_regin ( logical_tile_clb_mode_default__fle_3_fle_regout ) , 
    .fle_scin ( logical_tile_clb_mode_default__fle_3_fle_scout ) , 
    .fle_clk ( clb_clk ) , 
    .ccff_head ( logical_tile_clb_mode_default__fle_3_ccff_tail ) ,
    .fle_out ( { clb_O[9] , logical_tile_clb_mode_default__fle_4_fle_out[1] } ) ,
    .fle_regout ( logical_tile_clb_mode_default__fle_4_fle_regout ) , 
    .fle_scout ( logical_tile_clb_mode_default__fle_4_fle_scout ) , 
    .ccff_tail ( logical_tile_clb_mode_default__fle_4_ccff_tail ) , 
    .p1 ( p2 ) , .p3 ( p4 ) ) ;
logical_tile_clb_mode_default__fle_5 logical_tile_clb_mode_default__fle_5 ( 
    .prog_clk ( prog_clk ) , .Test_en ( Test_en ) , .clk ( clk ) , 
    .fle_in ( clb_I5 ) , 
    .fle_regin ( logical_tile_clb_mode_default__fle_4_fle_regout ) , 
    .fle_scin ( logical_tile_clb_mode_default__fle_4_fle_scout ) , 
    .fle_clk ( clb_clk ) , 
    .ccff_head ( logical_tile_clb_mode_default__fle_4_ccff_tail ) ,
    .fle_out ( { logical_tile_clb_mode_default__fle_5_fle_out[0] , clb_O[10] } ) ,
    .fle_regout ( logical_tile_clb_mode_default__fle_5_fle_regout ) , 
    .fle_scout ( logical_tile_clb_mode_default__fle_5_fle_scout ) , 
    .ccff_tail ( logical_tile_clb_mode_default__fle_5_ccff_tail ) , 
    .p1 ( p2 ) ) ;
logical_tile_clb_mode_default__fle_6 logical_tile_clb_mode_default__fle_6 ( 
    .prog_clk ( prog_clk ) , .Test_en ( Test_en ) , .clk ( clk ) , 
    .fle_in ( clb_I6 ) , 
    .fle_regin ( logical_tile_clb_mode_default__fle_5_fle_regout ) , 
    .fle_scin ( logical_tile_clb_mode_default__fle_5_fle_scout ) , 
    .fle_clk ( clb_clk ) , 
    .ccff_head ( logical_tile_clb_mode_default__fle_5_ccff_tail ) ,
    .fle_out ( { logical_tile_clb_mode_default__fle_6_fle_out[0] , clb_O[12] } ) ,
    .fle_regout ( logical_tile_clb_mode_default__fle_6_fle_regout ) , 
    .fle_scout ( logical_tile_clb_mode_default__fle_6_fle_scout ) , 
    .ccff_tail ( logical_tile_clb_mode_default__fle_6_ccff_tail ) , 
    .p1 ( p2 ) ) ;
logical_tile_clb_mode_default__fle logical_tile_clb_mode_default__fle_7 ( 
    .prog_clk ( prog_clk ) , .Test_en ( Test_en ) , .clk ( clk ) , 
    .fle_in ( clb_I7 ) , 
    .fle_regin ( logical_tile_clb_mode_default__fle_6_fle_regout ) , 
    .fle_scin ( logical_tile_clb_mode_default__fle_6_fle_scout ) , 
    .fle_clk ( clb_clk ) , 
    .ccff_head ( logical_tile_clb_mode_default__fle_6_ccff_tail ) ,
    .fle_out ( { p_abuf14 , clb_O[14] } ) ,
    .fle_regout ( clb_regout ) , .fle_scout ( clb_scout ) , 
    .ccff_tail ( ccff_tail ) , .p_abuf0 ( p_abuf16 ) , .p_abuf1 ( p_abuf17 ) , 
    .p2 ( p3 ) ) ;
direct_interc direct_interc_0_ (
    .in ( { SYNOPSYS_UNCONNECTED_1 } ) ,
    .out ( logical_tile_clb_mode_default__fle_0_fle_out ) ) ;
direct_interc direct_interc_1_ (
    .in ( { SYNOPSYS_UNCONNECTED_2 } ) ,
    .out ( clb_O[1] ) ) ;
direct_interc direct_interc_2_ (
    .in ( { SYNOPSYS_UNCONNECTED_3 } ) ,
    .out ( logical_tile_clb_mode_default__fle_1_fle_out ) ) ;
direct_interc direct_interc_3_ (
    .in ( { SYNOPSYS_UNCONNECTED_4 } ) ,
    .out ( clb_O[3] ) ) ;
direct_interc direct_interc_4_ (
    .in ( { SYNOPSYS_UNCONNECTED_5 } ) ,
    .out ( clb_O[4] ) ) ;
direct_interc direct_interc_5_ (
    .in ( { SYNOPSYS_UNCONNECTED_6 } ) ,
    .out ( clb_O[5] ) ) ;
direct_interc direct_interc_6_ (
    .in ( { SYNOPSYS_UNCONNECTED_7 } ) ,
    .out ( logical_tile_clb_mode_default__fle_3_fle_out[1] ) ) ;
direct_interc direct_interc_7_ (
    .in ( { SYNOPSYS_UNCONNECTED_8 } ) ,
    .out ( logical_tile_clb_mode_default__fle_3_fle_out[0] ) ) ;
direct_interc direct_interc_8_ (
    .in ( { SYNOPSYS_UNCONNECTED_9 } ) ,
    .out ( logical_tile_clb_mode_default__fle_4_fle_out ) ) ;
direct_interc direct_interc_9_ (
    .in ( { SYNOPSYS_UNCONNECTED_10 } ) ,
    .out ( clb_O[9] ) ) ;
direct_interc direct_interc_10_ (
    .in ( { SYNOPSYS_UNCONNECTED_11 } ) ,
    .out ( clb_O[10] ) ) ;
direct_interc direct_interc_11_ (
    .in ( { SYNOPSYS_UNCONNECTED_12 } ) ,
    .out ( logical_tile_clb_mode_default__fle_5_fle_out ) ) ;
direct_interc direct_interc_12_ (
    .in ( { SYNOPSYS_UNCONNECTED_13 } ) ,
    .out ( clb_O[12] ) ) ;
direct_interc direct_interc_13_ (
    .in ( { SYNOPSYS_UNCONNECTED_14 } ) ,
    .out ( logical_tile_clb_mode_default__fle_6_fle_out ) ) ;
direct_interc direct_interc_14_ (
    .in ( { SYNOPSYS_UNCONNECTED_15 } ) ,
    .out ( clb_O[14] ) ) ;
direct_interc direct_interc_15_ (
    .in ( { SYNOPSYS_UNCONNECTED_16 } ) ,
    .out ( { p_abuf14 } ) ) ;
direct_interc direct_interc_16_ (
    .in ( { SYNOPSYS_UNCONNECTED_17 } ) ,
    .out ( { p_abuf16 } ) ) ;
direct_interc direct_interc_17_ (
    .in ( { SYNOPSYS_UNCONNECTED_18 } ) ,
    .out ( { p_abuf17 } ) ) ;
direct_interc direct_interc_18_ (
    .in ( { SYNOPSYS_UNCONNECTED_19 } ) ,
    .out ( clb_I0[0] ) ) ;
direct_interc direct_interc_19_ (
    .in ( { SYNOPSYS_UNCONNECTED_20 } ) ,
    .out ( clb_I0[1] ) ) ;
direct_interc direct_interc_20_ (
    .in ( { SYNOPSYS_UNCONNECTED_21 } ) ,
    .out ( clb_I0[2] ) ) ;
direct_interc direct_interc_21_ (
    .in ( { SYNOPSYS_UNCONNECTED_22 } ) ,
    .out ( clb_I0[3] ) ) ;
direct_interc direct_interc_22_ (
    .in ( { SYNOPSYS_UNCONNECTED_23 } ) ,
    .out ( clb_regin ) ) ;
direct_interc direct_interc_23_ (
    .in ( { SYNOPSYS_UNCONNECTED_24 } ) ,
    .out ( clb_scin ) ) ;
direct_interc direct_interc_24_ (
    .in ( { SYNOPSYS_UNCONNECTED_25 } ) ,
    .out ( clb_clk ) ) ;
direct_interc direct_interc_25_ (
    .in ( { SYNOPSYS_UNCONNECTED_26 } ) ,
    .out ( clb_I1[0] ) ) ;
direct_interc direct_interc_26_ (
    .in ( { SYNOPSYS_UNCONNECTED_27 } ) ,
    .out ( clb_I1[1] ) ) ;
direct_interc direct_interc_27_ (
    .in ( { SYNOPSYS_UNCONNECTED_28 } ) ,
    .out ( clb_I1[2] ) ) ;
direct_interc direct_interc_28_ (
    .in ( { SYNOPSYS_UNCONNECTED_29 } ) ,
    .out ( clb_I1[3] ) ) ;
direct_interc direct_interc_29_ (
    .in ( { SYNOPSYS_UNCONNECTED_30 } ) ,
    .out ( logical_tile_clb_mode_default__fle_0_fle_regout ) ) ;
direct_interc direct_interc_30_ (
    .in ( { SYNOPSYS_UNCONNECTED_31 } ) ,
    .out ( logical_tile_clb_mode_default__fle_0_fle_scout ) ) ;
direct_interc direct_interc_31_ (
    .in ( { SYNOPSYS_UNCONNECTED_32 } ) ,
    .out ( clb_clk ) ) ;
direct_interc direct_interc_32_ (
    .in ( { SYNOPSYS_UNCONNECTED_33 } ) ,
    .out ( clb_I2[0] ) ) ;
direct_interc direct_interc_33_ (
    .in ( { SYNOPSYS_UNCONNECTED_34 } ) ,
    .out ( clb_I2[1] ) ) ;
direct_interc direct_interc_34_ (
    .in ( { SYNOPSYS_UNCONNECTED_35 } ) ,
    .out ( clb_I2[2] ) ) ;
direct_interc direct_interc_35_ (
    .in ( { SYNOPSYS_UNCONNECTED_36 } ) ,
    .out ( clb_I2[3] ) ) ;
direct_interc direct_interc_36_ (
    .in ( { SYNOPSYS_UNCONNECTED_37 } ) ,
    .out ( logical_tile_clb_mode_default__fle_1_fle_regout ) ) ;
direct_interc direct_interc_37_ (
    .in ( { SYNOPSYS_UNCONNECTED_38 } ) ,
    .out ( logical_tile_clb_mode_default__fle_1_fle_scout ) ) ;
direct_interc direct_interc_38_ (
    .in ( { SYNOPSYS_UNCONNECTED_39 } ) ,
    .out ( clb_clk ) ) ;
direct_interc direct_interc_39_ (
    .in ( { SYNOPSYS_UNCONNECTED_40 } ) ,
    .out ( clb_I3[0] ) ) ;
direct_interc direct_interc_40_ (
    .in ( { SYNOPSYS_UNCONNECTED_41 } ) ,
    .out ( clb_I3[1] ) ) ;
direct_interc direct_interc_41_ (
    .in ( { SYNOPSYS_UNCONNECTED_42 } ) ,
    .out ( clb_I3[2] ) ) ;
direct_interc direct_interc_42_ (
    .in ( { SYNOPSYS_UNCONNECTED_43 } ) ,
    .out ( clb_I3[3] ) ) ;
direct_interc direct_interc_43_ (
    .in ( { SYNOPSYS_UNCONNECTED_44 } ) ,
    .out ( logical_tile_clb_mode_default__fle_2_fle_regout ) ) ;
direct_interc direct_interc_44_ (
    .in ( { SYNOPSYS_UNCONNECTED_45 } ) ,
    .out ( logical_tile_clb_mode_default__fle_2_fle_scout ) ) ;
direct_interc direct_interc_45_ (
    .in ( { SYNOPSYS_UNCONNECTED_46 } ) ,
    .out ( clb_clk ) ) ;
direct_interc direct_interc_46_ (
    .in ( { SYNOPSYS_UNCONNECTED_47 } ) ,
    .out ( clb_I4[0] ) ) ;
direct_interc direct_interc_47_ (
    .in ( { SYNOPSYS_UNCONNECTED_48 } ) ,
    .out ( clb_I4[1] ) ) ;
direct_interc direct_interc_48_ (
    .in ( { SYNOPSYS_UNCONNECTED_49 } ) ,
    .out ( clb_I4[2] ) ) ;
direct_interc direct_interc_49_ (
    .in ( { SYNOPSYS_UNCONNECTED_50 } ) ,
    .out ( clb_I4[3] ) ) ;
direct_interc direct_interc_50_ (
    .in ( { SYNOPSYS_UNCONNECTED_51 } ) ,
    .out ( logical_tile_clb_mode_default__fle_3_fle_regout ) ) ;
direct_interc direct_interc_51_ (
    .in ( { SYNOPSYS_UNCONNECTED_52 } ) ,
    .out ( logical_tile_clb_mode_default__fle_3_fle_scout ) ) ;
direct_interc direct_interc_52_ (
    .in ( { SYNOPSYS_UNCONNECTED_53 } ) ,
    .out ( clb_clk ) ) ;
direct_interc direct_interc_53_ (
    .in ( { SYNOPSYS_UNCONNECTED_54 } ) ,
    .out ( clb_I5[0] ) ) ;
direct_interc direct_interc_54_ (
    .in ( { SYNOPSYS_UNCONNECTED_55 } ) ,
    .out ( clb_I5[1] ) ) ;
direct_interc direct_interc_55_ (
    .in ( { SYNOPSYS_UNCONNECTED_56 } ) ,
    .out ( clb_I5[2] ) ) ;
direct_interc direct_interc_56_ (
    .in ( { SYNOPSYS_UNCONNECTED_57 } ) ,
    .out ( clb_I5[3] ) ) ;
direct_interc direct_interc_57_ (
    .in ( { SYNOPSYS_UNCONNECTED_58 } ) ,
    .out ( logical_tile_clb_mode_default__fle_4_fle_regout ) ) ;
direct_interc direct_interc_58_ (
    .in ( { SYNOPSYS_UNCONNECTED_59 } ) ,
    .out ( logical_tile_clb_mode_default__fle_4_fle_scout ) ) ;
direct_interc direct_interc_59_ (
    .in ( { SYNOPSYS_UNCONNECTED_60 } ) ,
    .out ( clb_clk ) ) ;
direct_interc direct_interc_60_ (
    .in ( { SYNOPSYS_UNCONNECTED_61 } ) ,
    .out ( clb_I6[0] ) ) ;
direct_interc direct_interc_61_ (
    .in ( { SYNOPSYS_UNCONNECTED_62 } ) ,
    .out ( clb_I6[1] ) ) ;
direct_interc direct_interc_62_ (
    .in ( { SYNOPSYS_UNCONNECTED_63 } ) ,
    .out ( clb_I6[2] ) ) ;
direct_interc direct_interc_63_ (
    .in ( { SYNOPSYS_UNCONNECTED_64 } ) ,
    .out ( clb_I6[3] ) ) ;
direct_interc direct_interc_64_ (
    .in ( { SYNOPSYS_UNCONNECTED_65 } ) ,
    .out ( logical_tile_clb_mode_default__fle_5_fle_regout ) ) ;
direct_interc direct_interc_65_ (
    .in ( { SYNOPSYS_UNCONNECTED_66 } ) ,
    .out ( logical_tile_clb_mode_default__fle_5_fle_scout ) ) ;
direct_interc direct_interc_66_ (
    .in ( { SYNOPSYS_UNCONNECTED_67 } ) ,
    .out ( clb_clk ) ) ;
direct_interc direct_interc_67_ (
    .in ( { SYNOPSYS_UNCONNECTED_68 } ) ,
    .out ( clb_I7[0] ) ) ;
direct_interc direct_interc_68_ (
    .in ( { SYNOPSYS_UNCONNECTED_69 } ) ,
    .out ( clb_I7[1] ) ) ;
direct_interc direct_interc_69_ (
    .in ( { SYNOPSYS_UNCONNECTED_70 } ) ,
    .out ( clb_I7[2] ) ) ;
direct_interc direct_interc_70_ (
    .in ( { SYNOPSYS_UNCONNECTED_71 } ) ,
    .out ( clb_I7[3] ) ) ;
direct_interc direct_interc_71_ (
    .in ( { SYNOPSYS_UNCONNECTED_72 } ) ,
    .out ( logical_tile_clb_mode_default__fle_6_fle_regout ) ) ;
direct_interc direct_interc_72_ (
    .in ( { SYNOPSYS_UNCONNECTED_73 } ) ,
    .out ( logical_tile_clb_mode_default__fle_6_fle_scout ) ) ;
direct_interc direct_interc_73_ (
    .in ( { SYNOPSYS_UNCONNECTED_74 } ) ,
    .out ( clb_clk ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_59 ( 
    .A ( logical_tile_clb_mode_default__fle_0_fle_out[1] ) , .X ( clb_O[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_58 ( .A ( clb_O[1] ) , .X ( p_abuf0 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_60 ( 
    .A ( logical_tile_clb_mode_default__fle_0_fle_out[1] ) , .X ( p_abuf1 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_63 ( 
    .A ( logical_tile_clb_mode_default__fle_1_fle_out[1] ) , .X ( clb_O[2] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_62 ( .A ( clb_O[3] ) , .X ( p_abuf2 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_64 ( 
    .A ( logical_tile_clb_mode_default__fle_1_fle_out[1] ) , .X ( p_abuf3 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_69 ( 
    .A ( logical_tile_clb_mode_default__fle_3_fle_out[0] ) , .X ( clb_O[7] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_66 ( .A ( clb_O[5] ) , .X ( p_abuf4 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_68 ( .A ( clb_O[4] ) , .X ( p_abuf5 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_70 ( 
    .A ( logical_tile_clb_mode_default__fle_3_fle_out[0] ) , .X ( p_abuf6 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_71 ( 
    .A ( logical_tile_clb_mode_default__fle_3_fle_out[1] ) , .X ( clb_O[6] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_72 ( 
    .A ( logical_tile_clb_mode_default__fle_3_fle_out[1] ) , .X ( p_abuf7 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_75 ( 
    .A ( logical_tile_clb_mode_default__fle_4_fle_out[1] ) , .X ( clb_O[8] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_74 ( .A ( clb_O[9] ) , 
    .X ( BUF_net_74 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_76 ( 
    .A ( logical_tile_clb_mode_default__fle_4_fle_out[1] ) , 
    .X ( BUF_net_76 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_77 ( 
    .A ( logical_tile_clb_mode_default__fle_5_fle_out[0] ) , 
    .X ( clb_O[11] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_78 ( 
    .A ( logical_tile_clb_mode_default__fle_5_fle_out[0] ) , 
    .X ( BUF_net_78 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_81 ( 
    .A ( logical_tile_clb_mode_default__fle_6_fle_out[0] ) , 
    .X ( clb_O[13] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_80 ( .A ( clb_O[10] ) , 
    .X ( BUF_net_80 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_82 ( 
    .A ( logical_tile_clb_mode_default__fle_6_fle_out[0] ) , 
    .X ( BUF_net_82 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_85 ( .A ( p_abuf14 ) , 
    .X ( BUF_net_85 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_84 ( .A ( clb_O[12] ) , 
    .X ( BUF_net_84 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_101 ( .A ( BUF_net_74 ) , 
    .X ( p_abuf8 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_87 ( .A ( clb_O[14] ) , 
    .X ( BUF_net_87 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_102 ( .A ( BUF_net_78 ) , 
    .X ( p_abuf10 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_103 ( .A ( BUF_net_85 ) , 
    .X ( clb_O[15] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_104 ( .A ( BUF_net_84 ) , 
    .X ( p_abuf13 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_105 ( .A ( BUF_net_87 ) , 
    .X ( p_abuf15 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_P_106 ( .A ( BUF_net_76 ) , 
    .X ( p_abuf9 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_P_107 ( .A ( BUF_net_80 ) , 
    .X ( p_abuf11 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_P_108 ( .A ( BUF_net_82 ) , 
    .X ( p_abuf12 ) ) ;
endmodule


module grid_clb ( prog_clk , Test_en , clk , top_width_0_height_0__pin_32_ , 
    top_width_0_height_0__pin_33_ , right_width_0_height_0__pin_0_ , 
    right_width_0_height_0__pin_1_ , right_width_0_height_0__pin_2_ , 
    right_width_0_height_0__pin_3_ , right_width_0_height_0__pin_4_ , 
    right_width_0_height_0__pin_5_ , right_width_0_height_0__pin_6_ , 
    right_width_0_height_0__pin_7_ , right_width_0_height_0__pin_8_ , 
    right_width_0_height_0__pin_9_ , right_width_0_height_0__pin_10_ , 
    right_width_0_height_0__pin_11_ , right_width_0_height_0__pin_12_ , 
    right_width_0_height_0__pin_13_ , right_width_0_height_0__pin_14_ , 
    right_width_0_height_0__pin_15_ , bottom_width_0_height_0__pin_16_ , 
    bottom_width_0_height_0__pin_17_ , bottom_width_0_height_0__pin_18_ , 
    bottom_width_0_height_0__pin_19_ , bottom_width_0_height_0__pin_20_ , 
    bottom_width_0_height_0__pin_21_ , bottom_width_0_height_0__pin_22_ , 
    bottom_width_0_height_0__pin_23_ , bottom_width_0_height_0__pin_24_ , 
    bottom_width_0_height_0__pin_25_ , bottom_width_0_height_0__pin_26_ , 
    bottom_width_0_height_0__pin_27_ , bottom_width_0_height_0__pin_28_ , 
    bottom_width_0_height_0__pin_29_ , bottom_width_0_height_0__pin_30_ , 
    bottom_width_0_height_0__pin_31_ , left_width_0_height_0__pin_52_ , 
    ccff_head , right_width_0_height_0__pin_34_upper , 
    right_width_0_height_0__pin_34_lower , 
    right_width_0_height_0__pin_35_upper , 
    right_width_0_height_0__pin_35_lower , 
    right_width_0_height_0__pin_36_upper , 
    right_width_0_height_0__pin_36_lower , 
    right_width_0_height_0__pin_37_upper , 
    right_width_0_height_0__pin_37_lower , 
    right_width_0_height_0__pin_38_upper , 
    right_width_0_height_0__pin_38_lower , 
    right_width_0_height_0__pin_39_upper , 
    right_width_0_height_0__pin_39_lower , 
    right_width_0_height_0__pin_40_upper , 
    right_width_0_height_0__pin_40_lower , 
    right_width_0_height_0__pin_41_upper , 
    right_width_0_height_0__pin_41_lower , 
    bottom_width_0_height_0__pin_42_upper , 
    bottom_width_0_height_0__pin_42_lower , 
    bottom_width_0_height_0__pin_43_upper , 
    bottom_width_0_height_0__pin_43_lower , 
    bottom_width_0_height_0__pin_44_upper , 
    bottom_width_0_height_0__pin_44_lower , 
    bottom_width_0_height_0__pin_45_upper , 
    bottom_width_0_height_0__pin_45_lower , 
    bottom_width_0_height_0__pin_46_upper , 
    bottom_width_0_height_0__pin_46_lower , 
    bottom_width_0_height_0__pin_47_upper , 
    bottom_width_0_height_0__pin_47_lower , 
    bottom_width_0_height_0__pin_48_upper , 
    bottom_width_0_height_0__pin_48_lower , 
    bottom_width_0_height_0__pin_49_upper , 
    bottom_width_0_height_0__pin_49_lower , bottom_width_0_height_0__pin_50_ , 
    bottom_width_0_height_0__pin_51_ , ccff_tail ) ;
input  [0:0] prog_clk ;
input  [0:0] Test_en ;
input  [0:0] clk ;
input  [0:0] top_width_0_height_0__pin_32_ ;
input  [0:0] top_width_0_height_0__pin_33_ ;
input  [0:0] right_width_0_height_0__pin_0_ ;
input  [0:0] right_width_0_height_0__pin_1_ ;
input  [0:0] right_width_0_height_0__pin_2_ ;
input  [0:0] right_width_0_height_0__pin_3_ ;
input  [0:0] right_width_0_height_0__pin_4_ ;
input  [0:0] right_width_0_height_0__pin_5_ ;
input  [0:0] right_width_0_height_0__pin_6_ ;
input  [0:0] right_width_0_height_0__pin_7_ ;
input  [0:0] right_width_0_height_0__pin_8_ ;
input  [0:0] right_width_0_height_0__pin_9_ ;
input  [0:0] right_width_0_height_0__pin_10_ ;
input  [0:0] right_width_0_height_0__pin_11_ ;
input  [0:0] right_width_0_height_0__pin_12_ ;
input  [0:0] right_width_0_height_0__pin_13_ ;
input  [0:0] right_width_0_height_0__pin_14_ ;
input  [0:0] right_width_0_height_0__pin_15_ ;
input  [0:0] bottom_width_0_height_0__pin_16_ ;
input  [0:0] bottom_width_0_height_0__pin_17_ ;
input  [0:0] bottom_width_0_height_0__pin_18_ ;
input  [0:0] bottom_width_0_height_0__pin_19_ ;
input  [0:0] bottom_width_0_height_0__pin_20_ ;
input  [0:0] bottom_width_0_height_0__pin_21_ ;
input  [0:0] bottom_width_0_height_0__pin_22_ ;
input  [0:0] bottom_width_0_height_0__pin_23_ ;
input  [0:0] bottom_width_0_height_0__pin_24_ ;
input  [0:0] bottom_width_0_height_0__pin_25_ ;
input  [0:0] bottom_width_0_height_0__pin_26_ ;
input  [0:0] bottom_width_0_height_0__pin_27_ ;
input  [0:0] bottom_width_0_height_0__pin_28_ ;
input  [0:0] bottom_width_0_height_0__pin_29_ ;
input  [0:0] bottom_width_0_height_0__pin_30_ ;
input  [0:0] bottom_width_0_height_0__pin_31_ ;
input  [0:0] left_width_0_height_0__pin_52_ ;
input  [0:0] ccff_head ;
output [0:0] right_width_0_height_0__pin_34_upper ;
output [0:0] right_width_0_height_0__pin_34_lower ;
output [0:0] right_width_0_height_0__pin_35_upper ;
output [0:0] right_width_0_height_0__pin_35_lower ;
output [0:0] right_width_0_height_0__pin_36_upper ;
output [0:0] right_width_0_height_0__pin_36_lower ;
output [0:0] right_width_0_height_0__pin_37_upper ;
output [0:0] right_width_0_height_0__pin_37_lower ;
output [0:0] right_width_0_height_0__pin_38_upper ;
output [0:0] right_width_0_height_0__pin_38_lower ;
output [0:0] right_width_0_height_0__pin_39_upper ;
output [0:0] right_width_0_height_0__pin_39_lower ;
output [0:0] right_width_0_height_0__pin_40_upper ;
output [0:0] right_width_0_height_0__pin_40_lower ;
output [0:0] right_width_0_height_0__pin_41_upper ;
output [0:0] right_width_0_height_0__pin_41_lower ;
output [0:0] bottom_width_0_height_0__pin_42_upper ;
output [0:0] bottom_width_0_height_0__pin_42_lower ;
output [0:0] bottom_width_0_height_0__pin_43_upper ;
output [0:0] bottom_width_0_height_0__pin_43_lower ;
output [0:0] bottom_width_0_height_0__pin_44_upper ;
output [0:0] bottom_width_0_height_0__pin_44_lower ;
output [0:0] bottom_width_0_height_0__pin_45_upper ;
output [0:0] bottom_width_0_height_0__pin_45_lower ;
output [0:0] bottom_width_0_height_0__pin_46_upper ;
output [0:0] bottom_width_0_height_0__pin_46_lower ;
output [0:0] bottom_width_0_height_0__pin_47_upper ;
output [0:0] bottom_width_0_height_0__pin_47_lower ;
output [0:0] bottom_width_0_height_0__pin_48_upper ;
output [0:0] bottom_width_0_height_0__pin_48_lower ;
output [0:0] bottom_width_0_height_0__pin_49_upper ;
output [0:0] bottom_width_0_height_0__pin_49_lower ;
output [0:0] bottom_width_0_height_0__pin_50_ ;
output [0:0] bottom_width_0_height_0__pin_51_ ;
output [0:0] ccff_tail ;

wire ropt_net_128 ;
wire ropt_net_134 ;
wire ropt_net_136 ;
wire ropt_net_147 ;
wire ropt_net_133 ;
wire ropt_net_144 ;
wire ropt_net_126 ;
wire ropt_net_130 ;
wire ropt_net_135 ;
wire p_abuf14 ;

logical_tile_clb_mode_clb_ logical_tile_clb_mode_clb__0 ( 
    .prog_clk ( prog_clk ) , .Test_en ( Test_en ) , .clk ( clk ) ,
    .clb_I0 ( { right_width_0_height_0__pin_0_[0] , 
        right_width_0_height_0__pin_1_[0] , 
        right_width_0_height_0__pin_2_[0] , 
        right_width_0_height_0__pin_3_[0] } ) ,
    .clb_I1 ( { right_width_0_height_0__pin_4_[0] , 
        right_width_0_height_0__pin_5_[0] , 
        right_width_0_height_0__pin_6_[0] , 
        right_width_0_height_0__pin_7_[0] } ) ,
    .clb_I2 ( { right_width_0_height_0__pin_8_[0] , 
        right_width_0_height_0__pin_9_[0] , 
        right_width_0_height_0__pin_10_[0] , 
        right_width_0_height_0__pin_11_[0] } ) ,
    .clb_I3 ( { right_width_0_height_0__pin_12_[0] , 
        right_width_0_height_0__pin_13_[0] , 
        right_width_0_height_0__pin_14_[0] , 
        right_width_0_height_0__pin_15_[0] } ) ,
    .clb_I4 ( { bottom_width_0_height_0__pin_16_[0] , 
        bottom_width_0_height_0__pin_17_[0] , 
        bottom_width_0_height_0__pin_18_[0] , 
        bottom_width_0_height_0__pin_19_[0] } ) ,
    .clb_I5 ( { bottom_width_0_height_0__pin_20_[0] , 
        bottom_width_0_height_0__pin_21_[0] , 
        bottom_width_0_height_0__pin_22_[0] , 
        bottom_width_0_height_0__pin_23_[0] } ) ,
    .clb_I6 ( { bottom_width_0_height_0__pin_24_[0] , 
        bottom_width_0_height_0__pin_25_[0] , 
        bottom_width_0_height_0__pin_26_[0] , 
        bottom_width_0_height_0__pin_27_[0] } ) ,
    .clb_I7 ( { bottom_width_0_height_0__pin_28_[0] , 
        bottom_width_0_height_0__pin_29_[0] , 
        bottom_width_0_height_0__pin_30_[0] , 
        bottom_width_0_height_0__pin_31_[0] } ) ,
    .clb_regin ( top_width_0_height_0__pin_32_ ) , 
    .clb_scin ( top_width_0_height_0__pin_33_ ) , 
    .clb_clk ( left_width_0_height_0__pin_52_ ) , .ccff_head ( ccff_head ) ,
    .clb_O ( { aps_rename_129_ , aps_rename_130_ , aps_rename_132_ , 
        aps_rename_134_ , aps_rename_136_ , aps_rename_138_ , 
        aps_rename_140_ , aps_rename_141_ , aps_rename_143_ , 
        aps_rename_145_ , aps_rename_147_ , aps_rename_149_ , 
        aps_rename_151_ , aps_rename_153_ , aps_rename_155_ , 
        bottom_width_0_height_0__pin_49_upper[0] } ) ,
    .clb_regout ( bottom_width_0_height_0__pin_50_ ) , 
    .clb_scout ( bottom_width_0_height_0__pin_51_ ) ,
    .ccff_tail ( { ropt_net_124 } ) ,
    .p_abuf0 ( right_width_0_height_0__pin_35_upper[0] ) , 
    .p_abuf1 ( right_width_0_height_0__pin_34_upper[0] ) , 
    .p_abuf2 ( ropt_net_134 ) , .p_abuf3 ( ropt_net_128 ) , 
    .p_abuf4 ( right_width_0_height_0__pin_39_upper[0] ) , 
    .p_abuf5 ( ropt_net_136 ) , .p_abuf6 ( ropt_net_133 ) , 
    .p_abuf7 ( ropt_net_147 ) , .p_abuf8 ( ropt_net_144 ) , 
    .p_abuf9 ( bottom_width_0_height_0__pin_42_upper[0] ) , 
    .p_abuf10 ( ropt_net_126 ) , 
    .p_abuf11 ( bottom_width_0_height_0__pin_44_upper[0] ) , 
    .p_abuf12 ( bottom_width_0_height_0__pin_47_upper[0] ) , 
    .p_abuf13 ( ropt_net_130 ) , .p_abuf14 ( p_abuf14 ) , 
    .p_abuf15 ( ropt_net_135 ) , .p0 ( optlc_net_118 ) , 
    .p1 ( optlc_net_119 ) , .p2 ( optlc_net_120 ) , .p3 ( optlc_net_121 ) , 
    .p4 ( optlc_net_122 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_1__0 ( .A ( aps_rename_129_ ) , 
    .X ( ropt_net_129 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_2__1 ( .A ( aps_rename_130_ ) , 
    .X ( aps_rename_131_ ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_3__2 ( .A ( aps_rename_132_ ) , 
    .X ( aps_rename_133_ ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_4__3 ( .A ( aps_rename_134_ ) , 
    .X ( aps_rename_135_ ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_5__4 ( .A ( aps_rename_136_ ) , 
    .X ( aps_rename_137_ ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_6__5 ( .A ( aps_rename_138_ ) , 
    .X ( aps_rename_139_ ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_7__6 ( .A ( aps_rename_140_ ) , 
    .X ( ropt_net_131 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_8__7 ( .A ( aps_rename_141_ ) , 
    .X ( aps_rename_142_ ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_9__8 ( .A ( aps_rename_143_ ) , 
    .X ( aps_rename_144_ ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_10__9 ( .A ( aps_rename_145_ ) , 
    .X ( aps_rename_146_ ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_11__10 ( .A ( aps_rename_147_ ) , 
    .X ( aps_rename_148_ ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_12__11 ( .A ( aps_rename_149_ ) , 
    .X ( aps_rename_150_ ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_13__12 ( .A ( aps_rename_151_ ) , 
    .X ( aps_rename_152_ ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 FTB_14__13 ( .A ( aps_rename_153_ ) , 
    .X ( aps_rename_154_ ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_15__14 ( .A ( aps_rename_155_ ) , 
    .X ( bottom_width_0_height_0__pin_48_lower[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 FTB_16__15 ( .A ( p_abuf14 ) , 
    .X ( bottom_width_0_height_0__pin_49_lower[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_89 ( .A ( aps_rename_131_ ) , 
    .X ( BUF_net_89 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_90 ( .A ( aps_rename_133_ ) , 
    .X ( ropt_net_132 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_91 ( .A ( aps_rename_135_ ) , 
    .X ( ropt_net_125 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_92 ( .A ( aps_rename_137_ ) , 
    .X ( right_width_0_height_0__pin_38_lower[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_93 ( .A ( aps_rename_139_ ) , 
    .X ( ropt_net_137 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_94 ( .A ( aps_rename_142_ ) , 
    .X ( right_width_0_height_0__pin_41_lower[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_RR_95 ( .A ( aps_rename_144_ ) , 
    .X ( bottom_width_0_height_0__pin_42_lower[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_96 ( .A ( aps_rename_146_ ) , 
    .X ( BUF_net_96 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_97 ( .A ( aps_rename_148_ ) , 
    .X ( BUF_net_97 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_98 ( .A ( aps_rename_150_ ) , 
    .X ( ropt_net_138 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_99 ( .A ( aps_rename_152_ ) , 
    .X ( BUF_net_99 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_RR_100 ( .A ( aps_rename_154_ ) , 
    .X ( ropt_net_127 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 BUFT_P_110 ( .A ( BUF_net_89 ) , 
    .X ( ropt_net_146 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_P_111 ( .A ( BUF_net_96 ) , 
    .X ( bottom_width_0_height_0__pin_43_lower[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_P_112 ( .A ( BUF_net_97 ) , 
    .X ( bottom_width_0_height_0__pin_44_lower[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 BUFT_P_113 ( .A ( BUF_net_99 ) , 
    .X ( bottom_width_0_height_0__pin_46_lower[0] ) ) ;
sky130_fd_sc_hd__conb_1 optlc_119 ( .LO ( SYNOPSYS_UNCONNECTED_1 ) , 
    .HI ( optlc_net_118 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_122 ( .LO ( SYNOPSYS_UNCONNECTED_2 ) , 
    .HI ( optlc_net_119 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_125 ( .LO ( SYNOPSYS_UNCONNECTED_3 ) , 
    .HI ( optlc_net_120 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_127 ( .LO ( SYNOPSYS_UNCONNECTED_4 ) , 
    .HI ( optlc_net_121 ) ) ;
sky130_fd_sc_hd__conb_1 optlc_129 ( .LO ( SYNOPSYS_UNCONNECTED_5 ) , 
    .HI ( optlc_net_122 ) ) ;
sky130_fd_sc_hd__dlymetal6s2s_1 ropt_mt_inst_878 ( .A ( ropt_net_124 ) , 
    .X ( ropt_net_139 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 ropt_mt_inst_879 ( .A ( ropt_net_125 ) , 
    .X ( right_width_0_height_0__pin_37_lower[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 ropt_mt_inst_880 ( .A ( ropt_net_126 ) , 
    .X ( ropt_net_140 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 ropt_mt_inst_881 ( .A ( ropt_net_127 ) , 
    .X ( bottom_width_0_height_0__pin_47_lower[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 ropt_mt_inst_882 ( .A ( ropt_net_128 ) , 
    .X ( right_width_0_height_0__pin_36_upper[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 ropt_mt_inst_884 ( .A ( ropt_net_129 ) , 
    .X ( ropt_net_143 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 ropt_mt_inst_885 ( .A ( ropt_net_130 ) , 
    .X ( bottom_width_0_height_0__pin_46_upper[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 ropt_mt_inst_886 ( .A ( ropt_net_131 ) , 
    .X ( right_width_0_height_0__pin_40_lower[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 ropt_mt_inst_887 ( .A ( ropt_net_132 ) , 
    .X ( ropt_net_142 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 ropt_mt_inst_888 ( .A ( ropt_net_133 ) , 
    .X ( right_width_0_height_0__pin_41_upper[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 ropt_mt_inst_890 ( .A ( ropt_net_134 ) , 
    .X ( right_width_0_height_0__pin_37_upper[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 ropt_mt_inst_892 ( .A ( ropt_net_135 ) , 
    .X ( bottom_width_0_height_0__pin_48_upper[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 ropt_mt_inst_895 ( .A ( ropt_net_136 ) , 
    .X ( ropt_net_145 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 ropt_mt_inst_898 ( .A ( ropt_net_137 ) , 
    .X ( ropt_net_141 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 ropt_mt_inst_909 ( .A ( ropt_net_138 ) , 
    .X ( bottom_width_0_height_0__pin_45_lower[0] ) ) ;
sky130_fd_sc_hd__dlymetal6s6s_1 ropt_mt_inst_913 ( .A ( ropt_net_139 ) , 
    .X ( ccff_tail[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 ropt_mt_inst_914 ( .A ( ropt_net_140 ) , 
    .X ( bottom_width_0_height_0__pin_45_upper[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 ropt_mt_inst_915 ( .A ( ropt_net_141 ) , 
    .X ( right_width_0_height_0__pin_39_lower[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 ropt_mt_inst_916 ( .A ( ropt_net_142 ) , 
    .X ( right_width_0_height_0__pin_36_lower[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 ropt_mt_inst_917 ( .A ( ropt_net_143 ) , 
    .X ( right_width_0_height_0__pin_34_lower[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 ropt_mt_inst_918 ( .A ( ropt_net_144 ) , 
    .X ( bottom_width_0_height_0__pin_43_upper[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 ropt_mt_inst_919 ( .A ( ropt_net_145 ) , 
    .X ( right_width_0_height_0__pin_38_upper[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 ropt_mt_inst_920 ( .A ( ropt_net_146 ) , 
    .X ( right_width_0_height_0__pin_35_lower[0] ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 ropt_mt_inst_921 ( .A ( ropt_net_147 ) , 
    .X ( right_width_0_height_0__pin_40_upper[0] ) ) ;
endmodule


module fpga_core ( prog_clk , Test_en , clk , gfpga_pad_GPIO_A , 
    gfpga_pad_GPIO_IE , gfpga_pad_GPIO_OE , gfpga_pad_GPIO_Y , ccff_head , 
    ccff_tail ) ;
input  [0:0] prog_clk ;
input  [0:0] Test_en ;
input  [0:0] clk ;
output [0:7] gfpga_pad_GPIO_A ;
output [0:7] gfpga_pad_GPIO_IE ;
output [0:7] gfpga_pad_GPIO_OE ;
inout  [0:7] gfpga_pad_GPIO_Y ;
input  [0:0] ccff_head ;
output [0:0] ccff_tail ;

wire [0:0] cbx_1__0__0_bottom_grid_pin_0_ ;
wire [0:0] cbx_1__0__0_ccff_tail ;
wire [0:19] cbx_1__0__0_chanx_left_out ;
wire [0:19] cbx_1__0__0_chanx_right_out ;
wire [0:0] cbx_1__0__0_top_grid_pin_16_ ;
wire [0:0] cbx_1__0__0_top_grid_pin_17_ ;
wire [0:0] cbx_1__0__0_top_grid_pin_18_ ;
wire [0:0] cbx_1__0__0_top_grid_pin_19_ ;
wire [0:0] cbx_1__0__0_top_grid_pin_20_ ;
wire [0:0] cbx_1__0__0_top_grid_pin_21_ ;
wire [0:0] cbx_1__0__0_top_grid_pin_22_ ;
wire [0:0] cbx_1__0__0_top_grid_pin_23_ ;
wire [0:0] cbx_1__0__0_top_grid_pin_24_ ;
wire [0:0] cbx_1__0__0_top_grid_pin_25_ ;
wire [0:0] cbx_1__0__0_top_grid_pin_26_ ;
wire [0:0] cbx_1__0__0_top_grid_pin_27_ ;
wire [0:0] cbx_1__0__0_top_grid_pin_28_ ;
wire [0:0] cbx_1__0__0_top_grid_pin_29_ ;
wire [0:0] cbx_1__0__0_top_grid_pin_30_ ;
wire [0:0] cbx_1__0__0_top_grid_pin_31_ ;
wire [0:0] cbx_1__0__1_bottom_grid_pin_0_ ;
wire [0:0] cbx_1__0__1_ccff_tail ;
wire [0:19] cbx_1__0__1_chanx_left_out ;
wire [0:19] cbx_1__0__1_chanx_right_out ;
wire [0:0] cbx_1__0__1_top_grid_pin_16_ ;
wire [0:0] cbx_1__0__1_top_grid_pin_17_ ;
wire [0:0] cbx_1__0__1_top_grid_pin_18_ ;
wire [0:0] cbx_1__0__1_top_grid_pin_19_ ;
wire [0:0] cbx_1__0__1_top_grid_pin_20_ ;
wire [0:0] cbx_1__0__1_top_grid_pin_21_ ;
wire [0:0] cbx_1__0__1_top_grid_pin_22_ ;
wire [0:0] cbx_1__0__1_top_grid_pin_23_ ;
wire [0:0] cbx_1__0__1_top_grid_pin_24_ ;
wire [0:0] cbx_1__0__1_top_grid_pin_25_ ;
wire [0:0] cbx_1__0__1_top_grid_pin_26_ ;
wire [0:0] cbx_1__0__1_top_grid_pin_27_ ;
wire [0:0] cbx_1__0__1_top_grid_pin_28_ ;
wire [0:0] cbx_1__0__1_top_grid_pin_29_ ;
wire [0:0] cbx_1__0__1_top_grid_pin_30_ ;
wire [0:0] cbx_1__0__1_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__0_ccff_tail ;
wire [0:19] cbx_1__1__0_chanx_left_out ;
wire [0:19] cbx_1__1__0_chanx_right_out ;
wire [0:0] cbx_1__1__0_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__0_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__0_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__0_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__0_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__0_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__0_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__0_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__0_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__0_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__0_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__0_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__0_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__0_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__0_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__0_top_grid_pin_31_ ;
wire [0:0] cbx_1__1__1_ccff_tail ;
wire [0:19] cbx_1__1__1_chanx_left_out ;
wire [0:19] cbx_1__1__1_chanx_right_out ;
wire [0:0] cbx_1__1__1_top_grid_pin_16_ ;
wire [0:0] cbx_1__1__1_top_grid_pin_17_ ;
wire [0:0] cbx_1__1__1_top_grid_pin_18_ ;
wire [0:0] cbx_1__1__1_top_grid_pin_19_ ;
wire [0:0] cbx_1__1__1_top_grid_pin_20_ ;
wire [0:0] cbx_1__1__1_top_grid_pin_21_ ;
wire [0:0] cbx_1__1__1_top_grid_pin_22_ ;
wire [0:0] cbx_1__1__1_top_grid_pin_23_ ;
wire [0:0] cbx_1__1__1_top_grid_pin_24_ ;
wire [0:0] cbx_1__1__1_top_grid_pin_25_ ;
wire [0:0] cbx_1__1__1_top_grid_pin_26_ ;
wire [0:0] cbx_1__1__1_top_grid_pin_27_ ;
wire [0:0] cbx_1__1__1_top_grid_pin_28_ ;
wire [0:0] cbx_1__1__1_top_grid_pin_29_ ;
wire [0:0] cbx_1__1__1_top_grid_pin_30_ ;
wire [0:0] cbx_1__1__1_top_grid_pin_31_ ;
wire [0:0] cbx_1__2__0_ccff_tail ;
wire [0:19] cbx_1__2__0_chanx_left_out ;
wire [0:19] cbx_1__2__0_chanx_right_out ;
wire [0:0] cbx_1__2__0_top_grid_pin_0_ ;
wire [0:0] cbx_1__2__1_ccff_tail ;
wire [0:19] cbx_1__2__1_chanx_left_out ;
wire [0:19] cbx_1__2__1_chanx_right_out ;
wire [0:0] cbx_1__2__1_top_grid_pin_0_ ;
wire [0:0] cby_0__1__0_ccff_tail ;
wire [0:19] cby_0__1__0_chany_bottom_out ;
wire [0:19] cby_0__1__0_chany_top_out ;
wire [0:0] cby_0__1__0_left_grid_pin_0_ ;
wire [0:0] cby_0__1__0_right_grid_pin_52_ ;
wire [0:0] cby_0__1__1_ccff_tail ;
wire [0:19] cby_0__1__1_chany_bottom_out ;
wire [0:19] cby_0__1__1_chany_top_out ;
wire [0:0] cby_0__1__1_left_grid_pin_0_ ;
wire [0:0] cby_0__1__1_right_grid_pin_52_ ;
wire [0:0] cby_1__1__0_ccff_tail ;
wire [0:19] cby_1__1__0_chany_bottom_out ;
wire [0:19] cby_1__1__0_chany_top_out ;
wire [0:0] cby_1__1__0_left_grid_pin_0_ ;
wire [0:0] cby_1__1__0_left_grid_pin_10_ ;
wire [0:0] cby_1__1__0_left_grid_pin_11_ ;
wire [0:0] cby_1__1__0_left_grid_pin_12_ ;
wire [0:0] cby_1__1__0_left_grid_pin_13_ ;
wire [0:0] cby_1__1__0_left_grid_pin_14_ ;
wire [0:0] cby_1__1__0_left_grid_pin_15_ ;
wire [0:0] cby_1__1__0_left_grid_pin_1_ ;
wire [0:0] cby_1__1__0_left_grid_pin_2_ ;
wire [0:0] cby_1__1__0_left_grid_pin_3_ ;
wire [0:0] cby_1__1__0_left_grid_pin_4_ ;
wire [0:0] cby_1__1__0_left_grid_pin_5_ ;
wire [0:0] cby_1__1__0_left_grid_pin_6_ ;
wire [0:0] cby_1__1__0_left_grid_pin_7_ ;
wire [0:0] cby_1__1__0_left_grid_pin_8_ ;
wire [0:0] cby_1__1__0_left_grid_pin_9_ ;
wire [0:0] cby_1__1__0_right_grid_pin_52_ ;
wire [0:0] cby_1__1__1_ccff_tail ;
wire [0:19] cby_1__1__1_chany_bottom_out ;
wire [0:19] cby_1__1__1_chany_top_out ;
wire [0:0] cby_1__1__1_left_grid_pin_0_ ;
wire [0:0] cby_1__1__1_left_grid_pin_10_ ;
wire [0:0] cby_1__1__1_left_grid_pin_11_ ;
wire [0:0] cby_1__1__1_left_grid_pin_12_ ;
wire [0:0] cby_1__1__1_left_grid_pin_13_ ;
wire [0:0] cby_1__1__1_left_grid_pin_14_ ;
wire [0:0] cby_1__1__1_left_grid_pin_15_ ;
wire [0:0] cby_1__1__1_left_grid_pin_1_ ;
wire [0:0] cby_1__1__1_left_grid_pin_2_ ;
wire [0:0] cby_1__1__1_left_grid_pin_3_ ;
wire [0:0] cby_1__1__1_left_grid_pin_4_ ;
wire [0:0] cby_1__1__1_left_grid_pin_5_ ;
wire [0:0] cby_1__1__1_left_grid_pin_6_ ;
wire [0:0] cby_1__1__1_left_grid_pin_7_ ;
wire [0:0] cby_1__1__1_left_grid_pin_8_ ;
wire [0:0] cby_1__1__1_left_grid_pin_9_ ;
wire [0:0] cby_1__1__1_right_grid_pin_52_ ;
wire [0:0] cby_1__1__2_ccff_tail ;
wire [0:19] cby_1__1__2_chany_bottom_out ;
wire [0:19] cby_1__1__2_chany_top_out ;
wire [0:0] cby_1__1__2_left_grid_pin_0_ ;
wire [0:0] cby_1__1__2_left_grid_pin_10_ ;
wire [0:0] cby_1__1__2_left_grid_pin_11_ ;
wire [0:0] cby_1__1__2_left_grid_pin_12_ ;
wire [0:0] cby_1__1__2_left_grid_pin_13_ ;
wire [0:0] cby_1__1__2_left_grid_pin_14_ ;
wire [0:0] cby_1__1__2_left_grid_pin_15_ ;
wire [0:0] cby_1__1__2_left_grid_pin_1_ ;
wire [0:0] cby_1__1__2_left_grid_pin_2_ ;
wire [0:0] cby_1__1__2_left_grid_pin_3_ ;
wire [0:0] cby_1__1__2_left_grid_pin_4_ ;
wire [0:0] cby_1__1__2_left_grid_pin_5_ ;
wire [0:0] cby_1__1__2_left_grid_pin_6_ ;
wire [0:0] cby_1__1__2_left_grid_pin_7_ ;
wire [0:0] cby_1__1__2_left_grid_pin_8_ ;
wire [0:0] cby_1__1__2_left_grid_pin_9_ ;
wire [0:0] cby_1__1__2_right_grid_pin_52_ ;
wire [0:0] cby_1__1__3_ccff_tail ;
wire [0:19] cby_1__1__3_chany_bottom_out ;
wire [0:19] cby_1__1__3_chany_top_out ;
wire [0:0] cby_1__1__3_left_grid_pin_0_ ;
wire [0:0] cby_1__1__3_left_grid_pin_10_ ;
wire [0:0] cby_1__1__3_left_grid_pin_11_ ;
wire [0:0] cby_1__1__3_left_grid_pin_12_ ;
wire [0:0] cby_1__1__3_left_grid_pin_13_ ;
wire [0:0] cby_1__1__3_left_grid_pin_14_ ;
wire [0:0] cby_1__1__3_left_grid_pin_15_ ;
wire [0:0] cby_1__1__3_left_grid_pin_1_ ;
wire [0:0] cby_1__1__3_left_grid_pin_2_ ;
wire [0:0] cby_1__1__3_left_grid_pin_3_ ;
wire [0:0] cby_1__1__3_left_grid_pin_4_ ;
wire [0:0] cby_1__1__3_left_grid_pin_5_ ;
wire [0:0] cby_1__1__3_left_grid_pin_6_ ;
wire [0:0] cby_1__1__3_left_grid_pin_7_ ;
wire [0:0] cby_1__1__3_left_grid_pin_8_ ;
wire [0:0] cby_1__1__3_left_grid_pin_9_ ;
wire [0:0] cby_1__1__3_right_grid_pin_52_ ;
wire [0:0] direct_interc_0_out ;
wire [0:0] direct_interc_1_out ;
wire [0:0] direct_interc_2_out ;
wire [0:0] direct_interc_3_out ;
wire [0:0] direct_interc_4_out ;
wire [0:0] direct_interc_5_out ;
wire [0:0] grid_clb_0_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_0_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_0_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_0_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_0_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_0_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_0_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_0_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_0_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_0_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_0_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_0_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_0_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_0_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_0_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_0_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_0_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_0_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_0_ccff_tail ;
wire [0:0] grid_clb_0_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_0_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_0_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_0_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_0_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_0_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_0_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_0_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_0_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_0_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_0_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_0_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_0_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_0_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_0_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_0_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_1__2__undriven_top_width_0_height_0__pin_32_ ;
wire [0:0] grid_clb_1__2__undriven_top_width_0_height_0__pin_33_ ;
wire [0:0] grid_clb_1_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_1_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_1_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_1_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_1_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_1_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_1_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_1_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_1_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_1_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_1_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_1_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_1_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_1_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_1_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_1_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_1_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_1_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_1_ccff_tail ;
wire [0:0] grid_clb_1_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_1_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_1_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_1_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_1_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_1_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_1_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_1_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_1_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_1_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_1_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_1_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_1_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_1_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_1_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_1_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_2__1__undriven_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_2__1__undriven_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_2_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_2_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_2_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_2_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_2_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_2_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_2_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_2_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_2_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_2_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_2_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_2_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_2_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_2_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_2_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_2_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_2_ccff_tail ;
wire [0:0] grid_clb_2_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_2_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_2_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_2_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_2_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_2_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_2_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_2_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_2_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_2_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_2_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_2_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_2_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_2_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_2_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_2_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_clb_3_bottom_width_0_height_0__pin_42_lower ;
wire [0:0] grid_clb_3_bottom_width_0_height_0__pin_42_upper ;
wire [0:0] grid_clb_3_bottom_width_0_height_0__pin_43_lower ;
wire [0:0] grid_clb_3_bottom_width_0_height_0__pin_43_upper ;
wire [0:0] grid_clb_3_bottom_width_0_height_0__pin_44_lower ;
wire [0:0] grid_clb_3_bottom_width_0_height_0__pin_44_upper ;
wire [0:0] grid_clb_3_bottom_width_0_height_0__pin_45_lower ;
wire [0:0] grid_clb_3_bottom_width_0_height_0__pin_45_upper ;
wire [0:0] grid_clb_3_bottom_width_0_height_0__pin_46_lower ;
wire [0:0] grid_clb_3_bottom_width_0_height_0__pin_46_upper ;
wire [0:0] grid_clb_3_bottom_width_0_height_0__pin_47_lower ;
wire [0:0] grid_clb_3_bottom_width_0_height_0__pin_47_upper ;
wire [0:0] grid_clb_3_bottom_width_0_height_0__pin_48_lower ;
wire [0:0] grid_clb_3_bottom_width_0_height_0__pin_48_upper ;
wire [0:0] grid_clb_3_bottom_width_0_height_0__pin_49_lower ;
wire [0:0] grid_clb_3_bottom_width_0_height_0__pin_49_upper ;
wire [0:0] grid_clb_3_bottom_width_0_height_0__pin_50_ ;
wire [0:0] grid_clb_3_bottom_width_0_height_0__pin_51_ ;
wire [0:0] grid_clb_3_ccff_tail ;
wire [0:0] grid_clb_3_right_width_0_height_0__pin_34_lower ;
wire [0:0] grid_clb_3_right_width_0_height_0__pin_34_upper ;
wire [0:0] grid_clb_3_right_width_0_height_0__pin_35_lower ;
wire [0:0] grid_clb_3_right_width_0_height_0__pin_35_upper ;
wire [0:0] grid_clb_3_right_width_0_height_0__pin_36_lower ;
wire [0:0] grid_clb_3_right_width_0_height_0__pin_36_upper ;
wire [0:0] grid_clb_3_right_width_0_height_0__pin_37_lower ;
wire [0:0] grid_clb_3_right_width_0_height_0__pin_37_upper ;
wire [0:0] grid_clb_3_right_width_0_height_0__pin_38_lower ;
wire [0:0] grid_clb_3_right_width_0_height_0__pin_38_upper ;
wire [0:0] grid_clb_3_right_width_0_height_0__pin_39_lower ;
wire [0:0] grid_clb_3_right_width_0_height_0__pin_39_upper ;
wire [0:0] grid_clb_3_right_width_0_height_0__pin_40_lower ;
wire [0:0] grid_clb_3_right_width_0_height_0__pin_40_upper ;
wire [0:0] grid_clb_3_right_width_0_height_0__pin_41_lower ;
wire [0:0] grid_clb_3_right_width_0_height_0__pin_41_upper ;
wire [0:0] grid_io_bottom_0_ccff_tail ;
wire [0:0] grid_io_bottom_0_top_width_0_height_0__pin_1_lower ;
wire [0:0] grid_io_bottom_0_top_width_0_height_0__pin_1_upper ;
wire [0:0] grid_io_bottom_1_ccff_tail ;
wire [0:0] grid_io_bottom_1_top_width_0_height_0__pin_1_lower ;
wire [0:0] grid_io_bottom_1_top_width_0_height_0__pin_1_upper ;
wire [0:0] grid_io_left_0_ccff_tail ;
wire [0:0] grid_io_left_0_right_width_0_height_0__pin_1_lower ;
wire [0:0] grid_io_left_0_right_width_0_height_0__pin_1_upper ;
wire [0:0] grid_io_left_1_ccff_tail ;
wire [0:0] grid_io_left_1_right_width_0_height_0__pin_1_lower ;
wire [0:0] grid_io_left_1_right_width_0_height_0__pin_1_upper ;
wire [0:0] grid_io_right_0_ccff_tail ;
wire [0:0] grid_io_right_0_left_width_0_height_0__pin_1_lower ;
wire [0:0] grid_io_right_0_left_width_0_height_0__pin_1_upper ;
wire [0:0] grid_io_right_1_ccff_tail ;
wire [0:0] grid_io_right_1_left_width_0_height_0__pin_1_lower ;
wire [0:0] grid_io_right_1_left_width_0_height_0__pin_1_upper ;
wire [0:0] grid_io_top_0_bottom_width_0_height_0__pin_1_lower ;
wire [0:0] grid_io_top_0_bottom_width_0_height_0__pin_1_upper ;
wire [0:0] grid_io_top_0_ccff_tail ;
wire [0:0] grid_io_top_1_bottom_width_0_height_0__pin_1_lower ;
wire [0:0] grid_io_top_1_bottom_width_0_height_0__pin_1_upper ;
wire [0:0] grid_io_top_1_ccff_tail ;
wire [0:19] sb_0__0__0_chanx_right_out ;
wire [0:19] sb_0__0__0_chany_top_out ;
wire [0:0] sb_0__1__0_ccff_tail ;
wire [0:19] sb_0__1__0_chanx_right_out ;
wire [0:19] sb_0__1__0_chany_bottom_out ;
wire [0:19] sb_0__1__0_chany_top_out ;
wire [0:0] sb_0__2__0_ccff_tail ;
wire [0:19] sb_0__2__0_chanx_right_out ;
wire [0:19] sb_0__2__0_chany_bottom_out ;
wire [0:0] sb_1__0__0_ccff_tail ;
wire [0:19] sb_1__0__0_chanx_left_out ;
wire [0:19] sb_1__0__0_chanx_right_out ;
wire [0:19] sb_1__0__0_chany_top_out ;
wire [0:0] sb_1__1__0_ccff_tail ;
wire [0:19] sb_1__1__0_chanx_left_out ;
wire [0:19] sb_1__1__0_chanx_right_out ;
wire [0:19] sb_1__1__0_chany_bottom_out ;
wire [0:19] sb_1__1__0_chany_top_out ;
wire [0:0] sb_1__2__0_ccff_tail ;
wire [0:19] sb_1__2__0_chanx_left_out ;
wire [0:19] sb_1__2__0_chanx_right_out ;
wire [0:19] sb_1__2__0_chany_bottom_out ;
wire [0:0] sb_2__0__0_ccff_tail ;
wire [0:19] sb_2__0__0_chanx_left_out ;
wire [0:19] sb_2__0__0_chany_top_out ;
wire [0:0] sb_2__1__0_ccff_tail ;
wire [0:19] sb_2__1__0_chanx_left_out ;
wire [0:19] sb_2__1__0_chany_bottom_out ;
wire [0:19] sb_2__1__0_chany_top_out ;
wire [0:0] sb_2__2__0_ccff_tail ;
wire [0:19] sb_2__2__0_chanx_left_out ;
wire [0:19] sb_2__2__0_chany_bottom_out ;
//

grid_clb grid_clb_1__1_ (
    .prog_clk ( { ctsbuf_net_1722 } ) ,
    .Test_en ( Test_en ) , .clk ( clk ) , 
    .top_width_0_height_0__pin_32_ ( direct_interc_0_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_3_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__0_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__0_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__0_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__0_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__0_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__0_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__0_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__0_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__0_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__0_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__0_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__0_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__0_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__0_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__0_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__0_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__0__0_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__0__0_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__0__0_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__0__0_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__0__0_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__0__0_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__0__0_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__0__0_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__0__0_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__0__0_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__0__0_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__0__0_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__0__0_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__0__0_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__0__0_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__0__0_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_0__1__0_right_grid_pin_52_ ) ,
    .ccff_head ( { ropt_net_31 } ) ,
    
    .right_width_0_height_0__pin_34_upper ( grid_clb_0_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_0_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_0_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_0_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_0_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_0_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_0_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_0_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_0_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_0_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_0_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_0_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_0_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_0_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_0_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_0_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_0_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_0_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_0_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_0_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_0_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_0_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_0_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_0_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_0_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_0_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_0_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_0_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_0_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_0_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_0_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_0_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_0_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_0_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_0_ccff_tail ) ) ;
grid_clb grid_clb_1__2_ (
    .prog_clk ( { ctsbuf_net_1318 } ) ,
    .Test_en ( Test_en ) , .clk ( clk ) , 
    .top_width_0_height_0__pin_32_ ( grid_clb_1__2__undriven_top_width_0_height_0__pin_32_ ) , 
    .top_width_0_height_0__pin_33_ ( grid_clb_1__2__undriven_top_width_0_height_0__pin_33_ ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__1_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__1_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__1_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__1_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__1_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__1_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__1_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__1_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__1_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__1_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__1_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__1_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__1_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__1_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__1_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__1_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__0_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__0_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__0_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__0_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__0_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__0_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__0_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__0_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__0_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__0_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__0_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__0_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__0_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__0_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__0_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__0_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_0__1__1_right_grid_pin_52_ ) ,
    .ccff_head ( { ropt_net_27 } ) ,
    
    .right_width_0_height_0__pin_34_upper ( grid_clb_1_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_1_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_1_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_1_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_1_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_1_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_1_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_1_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_1_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_1_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_1_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_1_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_1_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_1_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_1_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_1_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_1_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_1_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_1_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_1_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_1_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_1_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_1_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_1_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_1_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_1_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_1_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_1_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_1_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_1_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_1_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_1_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_1_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_1_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_1_ccff_tail ) ) ;
grid_clb grid_clb_2__1_ (
    .prog_clk ( { ctsbuf_net_1116 } ) ,
    .Test_en ( Test_en ) , .clk ( clk ) , 
    .top_width_0_height_0__pin_32_ ( direct_interc_1_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_4_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__2_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__2_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__2_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__2_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__2_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__2_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__2_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__2_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__2_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__2_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__2_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__2_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__2_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__2_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__2_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__2_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__0__1_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__0__1_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__0__1_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__0__1_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__0__1_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__0__1_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__0__1_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__0__1_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__0__1_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__0__1_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__0__1_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__0__1_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__0__1_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__0__1_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__0__1_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__0__1_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__0_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__0_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_2_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_2_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_2_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_2_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_2_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_2_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_2_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_2_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_2_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_2_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_2_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_2_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_2_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_2_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_2_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_2_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_2_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_2_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_2_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_2_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_2_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_2_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_2_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_2_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_2_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_2_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_2_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_2_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_2_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_2_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_2_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_2_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_2__1__undriven_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_2__1__undriven_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_2_ccff_tail ) ) ;
grid_clb grid_clb_2__2_ (
    .prog_clk ( { ctsbuf_net_510 } ) ,
    .Test_en ( Test_en ) , .clk ( clk ) , 
    .top_width_0_height_0__pin_32_ ( direct_interc_2_out ) , 
    .top_width_0_height_0__pin_33_ ( direct_interc_5_out ) , 
    .right_width_0_height_0__pin_0_ ( cby_1__1__3_left_grid_pin_0_ ) , 
    .right_width_0_height_0__pin_1_ ( cby_1__1__3_left_grid_pin_1_ ) , 
    .right_width_0_height_0__pin_2_ ( cby_1__1__3_left_grid_pin_2_ ) , 
    .right_width_0_height_0__pin_3_ ( cby_1__1__3_left_grid_pin_3_ ) , 
    .right_width_0_height_0__pin_4_ ( cby_1__1__3_left_grid_pin_4_ ) , 
    .right_width_0_height_0__pin_5_ ( cby_1__1__3_left_grid_pin_5_ ) , 
    .right_width_0_height_0__pin_6_ ( cby_1__1__3_left_grid_pin_6_ ) , 
    .right_width_0_height_0__pin_7_ ( cby_1__1__3_left_grid_pin_7_ ) , 
    .right_width_0_height_0__pin_8_ ( cby_1__1__3_left_grid_pin_8_ ) , 
    .right_width_0_height_0__pin_9_ ( cby_1__1__3_left_grid_pin_9_ ) , 
    .right_width_0_height_0__pin_10_ ( cby_1__1__3_left_grid_pin_10_ ) , 
    .right_width_0_height_0__pin_11_ ( cby_1__1__3_left_grid_pin_11_ ) , 
    .right_width_0_height_0__pin_12_ ( cby_1__1__3_left_grid_pin_12_ ) , 
    .right_width_0_height_0__pin_13_ ( cby_1__1__3_left_grid_pin_13_ ) , 
    .right_width_0_height_0__pin_14_ ( cby_1__1__3_left_grid_pin_14_ ) , 
    .right_width_0_height_0__pin_15_ ( cby_1__1__3_left_grid_pin_15_ ) , 
    .bottom_width_0_height_0__pin_16_ ( cbx_1__1__1_top_grid_pin_16_ ) , 
    .bottom_width_0_height_0__pin_17_ ( cbx_1__1__1_top_grid_pin_17_ ) , 
    .bottom_width_0_height_0__pin_18_ ( cbx_1__1__1_top_grid_pin_18_ ) , 
    .bottom_width_0_height_0__pin_19_ ( cbx_1__1__1_top_grid_pin_19_ ) , 
    .bottom_width_0_height_0__pin_20_ ( cbx_1__1__1_top_grid_pin_20_ ) , 
    .bottom_width_0_height_0__pin_21_ ( cbx_1__1__1_top_grid_pin_21_ ) , 
    .bottom_width_0_height_0__pin_22_ ( cbx_1__1__1_top_grid_pin_22_ ) , 
    .bottom_width_0_height_0__pin_23_ ( cbx_1__1__1_top_grid_pin_23_ ) , 
    .bottom_width_0_height_0__pin_24_ ( cbx_1__1__1_top_grid_pin_24_ ) , 
    .bottom_width_0_height_0__pin_25_ ( cbx_1__1__1_top_grid_pin_25_ ) , 
    .bottom_width_0_height_0__pin_26_ ( cbx_1__1__1_top_grid_pin_26_ ) , 
    .bottom_width_0_height_0__pin_27_ ( cbx_1__1__1_top_grid_pin_27_ ) , 
    .bottom_width_0_height_0__pin_28_ ( cbx_1__1__1_top_grid_pin_28_ ) , 
    .bottom_width_0_height_0__pin_29_ ( cbx_1__1__1_top_grid_pin_29_ ) , 
    .bottom_width_0_height_0__pin_30_ ( cbx_1__1__1_top_grid_pin_30_ ) , 
    .bottom_width_0_height_0__pin_31_ ( cbx_1__1__1_top_grid_pin_31_ ) , 
    .left_width_0_height_0__pin_52_ ( cby_1__1__1_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__1_ccff_tail ) , 
    .right_width_0_height_0__pin_34_upper ( grid_clb_3_right_width_0_height_0__pin_34_upper ) , 
    .right_width_0_height_0__pin_34_lower ( grid_clb_3_right_width_0_height_0__pin_34_lower ) , 
    .right_width_0_height_0__pin_35_upper ( grid_clb_3_right_width_0_height_0__pin_35_upper ) , 
    .right_width_0_height_0__pin_35_lower ( grid_clb_3_right_width_0_height_0__pin_35_lower ) , 
    .right_width_0_height_0__pin_36_upper ( grid_clb_3_right_width_0_height_0__pin_36_upper ) , 
    .right_width_0_height_0__pin_36_lower ( grid_clb_3_right_width_0_height_0__pin_36_lower ) , 
    .right_width_0_height_0__pin_37_upper ( grid_clb_3_right_width_0_height_0__pin_37_upper ) , 
    .right_width_0_height_0__pin_37_lower ( grid_clb_3_right_width_0_height_0__pin_37_lower ) , 
    .right_width_0_height_0__pin_38_upper ( grid_clb_3_right_width_0_height_0__pin_38_upper ) , 
    .right_width_0_height_0__pin_38_lower ( grid_clb_3_right_width_0_height_0__pin_38_lower ) , 
    .right_width_0_height_0__pin_39_upper ( grid_clb_3_right_width_0_height_0__pin_39_upper ) , 
    .right_width_0_height_0__pin_39_lower ( grid_clb_3_right_width_0_height_0__pin_39_lower ) , 
    .right_width_0_height_0__pin_40_upper ( grid_clb_3_right_width_0_height_0__pin_40_upper ) , 
    .right_width_0_height_0__pin_40_lower ( grid_clb_3_right_width_0_height_0__pin_40_lower ) , 
    .right_width_0_height_0__pin_41_upper ( grid_clb_3_right_width_0_height_0__pin_41_upper ) , 
    .right_width_0_height_0__pin_41_lower ( grid_clb_3_right_width_0_height_0__pin_41_lower ) , 
    .bottom_width_0_height_0__pin_42_upper ( grid_clb_3_bottom_width_0_height_0__pin_42_upper ) , 
    .bottom_width_0_height_0__pin_42_lower ( grid_clb_3_bottom_width_0_height_0__pin_42_lower ) , 
    .bottom_width_0_height_0__pin_43_upper ( grid_clb_3_bottom_width_0_height_0__pin_43_upper ) , 
    .bottom_width_0_height_0__pin_43_lower ( grid_clb_3_bottom_width_0_height_0__pin_43_lower ) , 
    .bottom_width_0_height_0__pin_44_upper ( grid_clb_3_bottom_width_0_height_0__pin_44_upper ) , 
    .bottom_width_0_height_0__pin_44_lower ( grid_clb_3_bottom_width_0_height_0__pin_44_lower ) , 
    .bottom_width_0_height_0__pin_45_upper ( grid_clb_3_bottom_width_0_height_0__pin_45_upper ) , 
    .bottom_width_0_height_0__pin_45_lower ( grid_clb_3_bottom_width_0_height_0__pin_45_lower ) , 
    .bottom_width_0_height_0__pin_46_upper ( grid_clb_3_bottom_width_0_height_0__pin_46_upper ) , 
    .bottom_width_0_height_0__pin_46_lower ( grid_clb_3_bottom_width_0_height_0__pin_46_lower ) , 
    .bottom_width_0_height_0__pin_47_upper ( grid_clb_3_bottom_width_0_height_0__pin_47_upper ) , 
    .bottom_width_0_height_0__pin_47_lower ( grid_clb_3_bottom_width_0_height_0__pin_47_lower ) , 
    .bottom_width_0_height_0__pin_48_upper ( grid_clb_3_bottom_width_0_height_0__pin_48_upper ) , 
    .bottom_width_0_height_0__pin_48_lower ( grid_clb_3_bottom_width_0_height_0__pin_48_lower ) , 
    .bottom_width_0_height_0__pin_49_upper ( grid_clb_3_bottom_width_0_height_0__pin_49_upper ) , 
    .bottom_width_0_height_0__pin_49_lower ( grid_clb_3_bottom_width_0_height_0__pin_49_lower ) , 
    .bottom_width_0_height_0__pin_50_ ( grid_clb_3_bottom_width_0_height_0__pin_50_ ) , 
    .bottom_width_0_height_0__pin_51_ ( grid_clb_3_bottom_width_0_height_0__pin_51_ ) , 
    .ccff_tail ( grid_clb_3_ccff_tail ) ) ;
grid_io_top grid_io_top_1__3_ (
    .prog_clk ( { ctsbuf_net_914 } ) ,
    .gfpga_pad_GPIO_A ( gfpga_pad_GPIO_A[0] ) , 
    .gfpga_pad_GPIO_IE ( gfpga_pad_GPIO_IE[0] ) , 
    .gfpga_pad_GPIO_OE ( gfpga_pad_GPIO_OE[0] ) , 
    .gfpga_pad_GPIO_Y ( gfpga_pad_GPIO_Y[0] ) , 
    .bottom_width_0_height_0__pin_0_ ( cbx_1__2__0_top_grid_pin_0_ ) , 
    .ccff_head ( cbx_1__2__0_ccff_tail ) , 
    .bottom_width_0_height_0__pin_1_upper ( grid_io_top_0_bottom_width_0_height_0__pin_1_upper ) , 
    .bottom_width_0_height_0__pin_1_lower ( grid_io_top_0_bottom_width_0_height_0__pin_1_lower ) , 
    .ccff_tail ( grid_io_top_0_ccff_tail ) ) ;
grid_io_top grid_io_top_2__3_ (
    .prog_clk ( { ctsbuf_net_38 } ) ,
    .gfpga_pad_GPIO_A ( gfpga_pad_GPIO_A[1] ) , 
    .gfpga_pad_GPIO_IE ( gfpga_pad_GPIO_IE[1] ) , 
    .gfpga_pad_GPIO_OE ( gfpga_pad_GPIO_OE[1] ) , 
    .gfpga_pad_GPIO_Y ( gfpga_pad_GPIO_Y[1] ) , 
    .bottom_width_0_height_0__pin_0_ ( cbx_1__2__1_top_grid_pin_0_ ) , 
    .ccff_head ( cbx_1__2__1_ccff_tail ) , 
    .bottom_width_0_height_0__pin_1_upper ( grid_io_top_1_bottom_width_0_height_0__pin_1_upper ) , 
    .bottom_width_0_height_0__pin_1_lower ( grid_io_top_1_bottom_width_0_height_0__pin_1_lower ) , 
    .ccff_tail ( grid_io_top_1_ccff_tail ) ) ;
grid_io_right grid_io_right_3__1_ (
    .prog_clk ( { ctsbuf_net_49 } ) ,
    .gfpga_pad_GPIO_A ( gfpga_pad_GPIO_A[2] ) , 
    .gfpga_pad_GPIO_IE ( gfpga_pad_GPIO_IE[2] ) , 
    .gfpga_pad_GPIO_OE ( gfpga_pad_GPIO_OE[2] ) , 
    .gfpga_pad_GPIO_Y ( gfpga_pad_GPIO_Y[2] ) , 
    .left_width_0_height_0__pin_0_ ( cby_1__1__2_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__2_ccff_tail ) , 
    .left_width_0_height_0__pin_1_upper ( grid_io_right_0_left_width_0_height_0__pin_1_upper ) , 
    .left_width_0_height_0__pin_1_lower ( grid_io_right_0_left_width_0_height_0__pin_1_lower ) , 
    .ccff_tail ( grid_io_right_0_ccff_tail ) ) ;
grid_io_right grid_io_right_3__2_ (
    .prog_clk ( { ctsbuf_net_16 } ) ,
    .gfpga_pad_GPIO_A ( gfpga_pad_GPIO_A[3] ) , 
    .gfpga_pad_GPIO_IE ( gfpga_pad_GPIO_IE[3] ) , 
    .gfpga_pad_GPIO_OE ( gfpga_pad_GPIO_OE[3] ) , 
    .gfpga_pad_GPIO_Y ( gfpga_pad_GPIO_Y[3] ) , 
    .left_width_0_height_0__pin_0_ ( cby_1__1__3_right_grid_pin_52_ ) , 
    .ccff_head ( cby_1__1__3_ccff_tail ) , 
    .left_width_0_height_0__pin_1_upper ( grid_io_right_1_left_width_0_height_0__pin_1_upper ) , 
    .left_width_0_height_0__pin_1_lower ( grid_io_right_1_left_width_0_height_0__pin_1_lower ) , 
    .ccff_tail ( grid_io_right_1_ccff_tail ) ) ;
grid_io_bottom grid_io_bottom_1__0_ (
    .prog_clk ( { ctsbuf_net_611 } ) ,
    .gfpga_pad_GPIO_A ( gfpga_pad_GPIO_A[4] ) , 
    .gfpga_pad_GPIO_IE ( gfpga_pad_GPIO_IE[4] ) , 
    .gfpga_pad_GPIO_OE ( gfpga_pad_GPIO_OE[4] ) , 
    .gfpga_pad_GPIO_Y ( gfpga_pad_GPIO_Y[4] ) , 
    .top_width_0_height_0__pin_0_ ( cbx_1__0__0_bottom_grid_pin_0_ ) , 
    .ccff_head ( cbx_1__0__0_ccff_tail ) , 
    .top_width_0_height_0__pin_1_upper ( grid_io_bottom_0_top_width_0_height_0__pin_1_upper ) , 
    .top_width_0_height_0__pin_1_lower ( grid_io_bottom_0_top_width_0_height_0__pin_1_lower ) , 
    .ccff_tail ( grid_io_bottom_0_ccff_tail ) ) ;
grid_io_bottom grid_io_bottom_2__0_ (
    .prog_clk ( { ctsbuf_net_27 } ) ,
    .gfpga_pad_GPIO_A ( gfpga_pad_GPIO_A[5] ) , 
    .gfpga_pad_GPIO_IE ( gfpga_pad_GPIO_IE[5] ) , 
    .gfpga_pad_GPIO_OE ( gfpga_pad_GPIO_OE[5] ) , 
    .gfpga_pad_GPIO_Y ( gfpga_pad_GPIO_Y[5] ) , 
    .top_width_0_height_0__pin_0_ ( cbx_1__0__1_bottom_grid_pin_0_ ) , 
    .ccff_head ( cbx_1__0__1_ccff_tail ) , 
    .top_width_0_height_0__pin_1_upper ( grid_io_bottom_1_top_width_0_height_0__pin_1_upper ) , 
    .top_width_0_height_0__pin_1_lower ( grid_io_bottom_1_top_width_0_height_0__pin_1_lower ) , 
    .ccff_tail ( grid_io_bottom_1_ccff_tail ) ) ;
grid_io_left grid_io_left_0__1_ (
    .prog_clk ( { ctsbuf_net_1520 } ) ,
    .gfpga_pad_GPIO_A ( gfpga_pad_GPIO_A[6] ) , 
    .gfpga_pad_GPIO_IE ( gfpga_pad_GPIO_IE[6] ) , 
    .gfpga_pad_GPIO_OE ( gfpga_pad_GPIO_OE[6] ) , 
    .gfpga_pad_GPIO_Y ( gfpga_pad_GPIO_Y[6] ) , 
    .right_width_0_height_0__pin_0_ ( cby_0__1__0_left_grid_pin_0_ ) , 
    .ccff_head ( cby_0__1__0_ccff_tail ) , 
    .right_width_0_height_0__pin_1_upper ( grid_io_left_0_right_width_0_height_0__pin_1_upper ) , 
    .right_width_0_height_0__pin_1_lower ( grid_io_left_0_right_width_0_height_0__pin_1_lower ) , 
    .ccff_tail ( grid_io_left_0_ccff_tail ) ) ;
grid_io_left grid_io_left_0__2_ (
    .prog_clk ( { ctsbuf_net_1419 } ) ,
    .gfpga_pad_GPIO_A ( gfpga_pad_GPIO_A[7] ) , 
    .gfpga_pad_GPIO_IE ( gfpga_pad_GPIO_IE[7] ) , 
    .gfpga_pad_GPIO_OE ( gfpga_pad_GPIO_OE[7] ) , 
    .gfpga_pad_GPIO_Y ( gfpga_pad_GPIO_Y[7] ) , 
    .right_width_0_height_0__pin_0_ ( cby_0__1__1_left_grid_pin_0_ ) , 
    .ccff_head ( cby_0__1__1_ccff_tail ) , 
    .right_width_0_height_0__pin_1_upper ( grid_io_left_1_right_width_0_height_0__pin_1_upper ) , 
    .right_width_0_height_0__pin_1_lower ( grid_io_left_1_right_width_0_height_0__pin_1_lower ) , 
    .ccff_tail ( grid_io_left_1_ccff_tail ) ) ;
sb_0__0_ sb_0__0_ (
    .prog_clk ( { ctsbuf_net_1520 } ) ,
    .chany_top_in ( cby_0__1__0_chany_bottom_out ) , 
    .top_left_grid_pin_1_ ( grid_io_left_0_right_width_0_height_0__pin_1_lower ) , 
    .chanx_right_in ( cbx_1__0__0_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_0_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_0_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_0_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_0_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_0_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_0_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_0_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_0_bottom_width_0_height_0__pin_49_upper ) , 
    .right_bottom_grid_pin_1_ ( grid_io_bottom_0_top_width_0_height_0__pin_1_upper ) , 
    .ccff_head ( grid_io_bottom_0_ccff_tail ) , 
    .chany_top_out ( sb_0__0__0_chany_top_out ) , 
    .chanx_right_out ( sb_0__0__0_chanx_right_out ) , 
    .ccff_tail ( ccff_tail ) ) ;
sb_0__1_ sb_0__1_ (
    .prog_clk ( { p_abuf0 } ) ,
    .chany_top_in ( cby_0__1__1_chany_bottom_out ) , 
    .top_left_grid_pin_1_ ( grid_io_left_1_right_width_0_height_0__pin_1_lower ) , 
    .chanx_right_in ( cbx_1__1__0_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_1_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_1_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_1_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_1_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_1_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_1_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_1_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_1_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_0__1__0_chany_top_out ) , 
    .bottom_left_grid_pin_1_ ( grid_io_left_0_right_width_0_height_0__pin_1_upper ) , 
    .ccff_head ( cbx_1__1__0_ccff_tail ) , 
    .chany_top_out ( sb_0__1__0_chany_top_out ) , 
    .chanx_right_out ( sb_0__1__0_chanx_right_out ) , 
    .chany_bottom_out ( sb_0__1__0_chany_bottom_out ) , 
    .ccff_tail ( sb_0__1__0_ccff_tail ) ) ;
sb_0__2_ sb_0__2_ (
    .prog_clk ( { ctsbuf_net_1419 } ) ,
    .chanx_right_in ( cbx_1__2__0_chanx_left_out ) , 
    .right_top_grid_pin_1_ ( grid_io_top_0_bottom_width_0_height_0__pin_1_upper ) , 
    .chany_bottom_in ( cby_0__1__1_chany_top_out ) , 
    .bottom_left_grid_pin_1_ ( grid_io_left_1_right_width_0_height_0__pin_1_upper ) , 
    .ccff_head ( grid_io_top_0_ccff_tail ) , 
    .chanx_right_out ( sb_0__2__0_chanx_right_out ) , 
    .chany_bottom_out ( sb_0__2__0_chany_bottom_out ) , 
    .ccff_tail ( sb_0__2__0_ccff_tail ) ) ;
sb_1__0_ sb_1__0_ (
    .prog_clk ( { ctsbuf_net_813 } ) ,
    .chany_top_in ( cby_1__1__0_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_0_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_0_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_0_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_0_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_0_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_0_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_0_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_0_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__0__1_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_2_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_2_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_2_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_2_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_2_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_2_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_2_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_2_bottom_width_0_height_0__pin_49_upper ) , 
    .right_bottom_grid_pin_1_ ( grid_io_bottom_1_top_width_0_height_0__pin_1_upper ) , 
    .chanx_left_in ( cbx_1__0__0_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_0_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_0_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_0_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_0_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_0_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_0_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_0_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_0_bottom_width_0_height_0__pin_49_lower ) , 
    .left_bottom_grid_pin_1_ ( grid_io_bottom_0_top_width_0_height_0__pin_1_lower ) , 
    .ccff_head ( grid_io_bottom_1_ccff_tail ) , 
    .chany_top_out ( sb_1__0__0_chany_top_out ) , 
    .chanx_right_out ( sb_1__0__0_chanx_right_out ) , 
    .chanx_left_out ( sb_1__0__0_chanx_left_out ) , 
    .ccff_tail ( sb_1__0__0_ccff_tail ) ) ;
sb_1__1_ sb_1__1_ (
    .prog_clk ( { ctsbuf_net_1217 } ) ,
    .chany_top_in ( cby_1__1__1_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_1_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_1_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_1_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_1_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_1_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_1_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_1_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_1_right_width_0_height_0__pin_41_lower ) , 
    .chanx_right_in ( cbx_1__1__1_chanx_left_out ) , 
    .right_top_grid_pin_42_ ( grid_clb_3_bottom_width_0_height_0__pin_42_upper ) , 
    .right_top_grid_pin_43_ ( grid_clb_3_bottom_width_0_height_0__pin_43_upper ) , 
    .right_top_grid_pin_44_ ( grid_clb_3_bottom_width_0_height_0__pin_44_upper ) , 
    .right_top_grid_pin_45_ ( grid_clb_3_bottom_width_0_height_0__pin_45_upper ) , 
    .right_top_grid_pin_46_ ( grid_clb_3_bottom_width_0_height_0__pin_46_upper ) , 
    .right_top_grid_pin_47_ ( grid_clb_3_bottom_width_0_height_0__pin_47_upper ) , 
    .right_top_grid_pin_48_ ( grid_clb_3_bottom_width_0_height_0__pin_48_upper ) , 
    .right_top_grid_pin_49_ ( grid_clb_3_bottom_width_0_height_0__pin_49_upper ) , 
    .chany_bottom_in ( cby_1__1__0_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_0_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_0_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_0_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_0_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_0_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_0_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_0_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_0_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__0_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_1_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_1_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_1_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_1_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_1_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_1_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_1_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_1_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( cbx_1__1__1_ccff_tail ) , 
    .chany_top_out ( sb_1__1__0_chany_top_out ) , 
    .chanx_right_out ( sb_1__1__0_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__1__0_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__1__0_chanx_left_out ) , 
    .ccff_tail ( sb_1__1__0_ccff_tail ) ) ;
sb_1__2_ sb_1__2_ (
    .prog_clk ( { ctsbuf_net_712 } ) ,
    .chanx_right_in ( cbx_1__2__1_chanx_left_out ) , 
    .right_top_grid_pin_1_ ( grid_io_top_1_bottom_width_0_height_0__pin_1_upper ) , 
    .chany_bottom_in ( cby_1__1__1_chany_top_out ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_1_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_1_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_1_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_1_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_1_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_1_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_1_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_1_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__2__0_chanx_right_out ) , 
    .left_top_grid_pin_1_ ( grid_io_top_0_bottom_width_0_height_0__pin_1_lower ) ,
    .ccff_head ( { ropt_net_29 } ) ,
    .chanx_right_out ( sb_1__2__0_chanx_right_out ) , 
    .chany_bottom_out ( sb_1__2__0_chany_bottom_out ) , 
    .chanx_left_out ( sb_1__2__0_chanx_left_out ) , 
    .ccff_tail ( sb_1__2__0_ccff_tail ) ) ;
sb_2__0_ sb_2__0_ (
    .prog_clk ( { ctsbuf_net_27 } ) ,
    .chany_top_in ( cby_1__1__2_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_2_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_2_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_2_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_2_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_2_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_2_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_2_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_2_right_width_0_height_0__pin_41_lower ) , 
    .top_right_grid_pin_1_ ( grid_io_right_0_left_width_0_height_0__pin_1_lower ) , 
    .chanx_left_in ( cbx_1__0__1_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_2_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_2_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_2_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_2_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_2_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_2_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_2_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_2_bottom_width_0_height_0__pin_49_lower ) , 
    .left_bottom_grid_pin_1_ ( grid_io_bottom_1_top_width_0_height_0__pin_1_lower ) , 
    .ccff_head ( grid_io_right_0_ccff_tail ) , 
    .chany_top_out ( sb_2__0__0_chany_top_out ) , 
    .chanx_left_out ( sb_2__0__0_chanx_left_out ) , 
    .ccff_tail ( sb_2__0__0_ccff_tail ) ) ;
sb_2__1_ sb_2__1_ (
    .prog_clk ( { ctsbuf_net_49 } ) ,
    .chany_top_in ( cby_1__1__3_chany_bottom_out ) , 
    .top_left_grid_pin_34_ ( grid_clb_3_right_width_0_height_0__pin_34_lower ) , 
    .top_left_grid_pin_35_ ( grid_clb_3_right_width_0_height_0__pin_35_lower ) , 
    .top_left_grid_pin_36_ ( grid_clb_3_right_width_0_height_0__pin_36_lower ) , 
    .top_left_grid_pin_37_ ( grid_clb_3_right_width_0_height_0__pin_37_lower ) , 
    .top_left_grid_pin_38_ ( grid_clb_3_right_width_0_height_0__pin_38_lower ) , 
    .top_left_grid_pin_39_ ( grid_clb_3_right_width_0_height_0__pin_39_lower ) , 
    .top_left_grid_pin_40_ ( grid_clb_3_right_width_0_height_0__pin_40_lower ) , 
    .top_left_grid_pin_41_ ( grid_clb_3_right_width_0_height_0__pin_41_lower ) , 
    .top_right_grid_pin_1_ ( grid_io_right_1_left_width_0_height_0__pin_1_lower ) , 
    .chany_bottom_in ( cby_1__1__2_chany_top_out ) , 
    .bottom_right_grid_pin_1_ ( grid_io_right_0_left_width_0_height_0__pin_1_upper ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_2_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_2_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_2_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_2_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_2_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_2_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_2_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_2_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__1__1_chanx_right_out ) , 
    .left_top_grid_pin_42_ ( grid_clb_3_bottom_width_0_height_0__pin_42_lower ) , 
    .left_top_grid_pin_43_ ( grid_clb_3_bottom_width_0_height_0__pin_43_lower ) , 
    .left_top_grid_pin_44_ ( grid_clb_3_bottom_width_0_height_0__pin_44_lower ) , 
    .left_top_grid_pin_45_ ( grid_clb_3_bottom_width_0_height_0__pin_45_lower ) , 
    .left_top_grid_pin_46_ ( grid_clb_3_bottom_width_0_height_0__pin_46_lower ) , 
    .left_top_grid_pin_47_ ( grid_clb_3_bottom_width_0_height_0__pin_47_lower ) , 
    .left_top_grid_pin_48_ ( grid_clb_3_bottom_width_0_height_0__pin_48_lower ) , 
    .left_top_grid_pin_49_ ( grid_clb_3_bottom_width_0_height_0__pin_49_lower ) , 
    .ccff_head ( grid_io_right_1_ccff_tail ) , 
    .chany_top_out ( sb_2__1__0_chany_top_out ) , 
    .chany_bottom_out ( sb_2__1__0_chany_bottom_out ) , 
    .chanx_left_out ( sb_2__1__0_chanx_left_out ) , 
    .ccff_tail ( sb_2__1__0_ccff_tail ) ) ;
sb_2__2_ sb_2__2_ (
    .prog_clk ( { ctsbuf_net_16 } ) ,
    .chany_bottom_in ( cby_1__1__3_chany_top_out ) , 
    .bottom_right_grid_pin_1_ ( grid_io_right_1_left_width_0_height_0__pin_1_upper ) , 
    .bottom_left_grid_pin_34_ ( grid_clb_3_right_width_0_height_0__pin_34_upper ) , 
    .bottom_left_grid_pin_35_ ( grid_clb_3_right_width_0_height_0__pin_35_upper ) , 
    .bottom_left_grid_pin_36_ ( grid_clb_3_right_width_0_height_0__pin_36_upper ) , 
    .bottom_left_grid_pin_37_ ( grid_clb_3_right_width_0_height_0__pin_37_upper ) , 
    .bottom_left_grid_pin_38_ ( grid_clb_3_right_width_0_height_0__pin_38_upper ) , 
    .bottom_left_grid_pin_39_ ( grid_clb_3_right_width_0_height_0__pin_39_upper ) , 
    .bottom_left_grid_pin_40_ ( grid_clb_3_right_width_0_height_0__pin_40_upper ) , 
    .bottom_left_grid_pin_41_ ( grid_clb_3_right_width_0_height_0__pin_41_upper ) , 
    .chanx_left_in ( cbx_1__2__1_chanx_right_out ) , 
    .left_top_grid_pin_1_ ( grid_io_top_1_bottom_width_0_height_0__pin_1_lower ) , 
    .ccff_head ( ccff_head ) , 
    .chany_bottom_out ( sb_2__2__0_chany_bottom_out ) , 
    .chanx_left_out ( sb_2__2__0_chanx_left_out ) , 
    .ccff_tail ( sb_2__2__0_ccff_tail ) ) ;
cbx_1__0_ cbx_1__0_ (
    .prog_clk ( { ctsbuf_net_611 } ) ,
    .chanx_left_in ( sb_0__0__0_chanx_right_out ) , 
    .chanx_right_in ( sb_1__0__0_chanx_left_out ) , 
    .ccff_head ( sb_1__0__0_ccff_tail ) , 
    .chanx_left_out ( cbx_1__0__0_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__0__0_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__0__0_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__0__0_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__0__0_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__0__0_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__0__0_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__0__0_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__0__0_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__0__0_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__0__0_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__0__0_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__0__0_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__0__0_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__0__0_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__0__0_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__0__0_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__0__0_top_grid_pin_31_ ) , 
    .bottom_grid_pin_0_ ( cbx_1__0__0_bottom_grid_pin_0_ ) , 
    .ccff_tail ( cbx_1__0__0_ccff_tail ) ) ;
cbx_1__0_ cbx_2__0_ (
    .prog_clk ( { ctsbuf_net_27 } ) ,
    .chanx_left_in ( sb_1__0__0_chanx_right_out ) , 
    .chanx_right_in ( sb_2__0__0_chanx_left_out ) , 
    .ccff_head ( sb_2__0__0_ccff_tail ) , 
    .chanx_left_out ( cbx_1__0__1_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__0__1_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__0__1_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__0__1_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__0__1_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__0__1_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__0__1_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__0__1_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__0__1_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__0__1_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__0__1_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__0__1_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__0__1_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__0__1_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__0__1_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__0__1_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__0__1_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__0__1_top_grid_pin_31_ ) , 
    .bottom_grid_pin_0_ ( cbx_1__0__1_bottom_grid_pin_0_ ) , 
    .ccff_tail ( cbx_1__0__1_ccff_tail ) ) ;
cbx_1__1_ cbx_1__1_ (
    .prog_clk ( { ctsbuf_net_1621 } ) ,
    .chanx_left_in ( sb_0__1__0_chanx_right_out ) , 
    .chanx_right_in ( sb_1__1__0_chanx_left_out ) , 
    .ccff_head ( sb_1__1__0_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__0_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__0_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__0_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__0_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__0_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__0_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__0_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__0_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__0_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__0_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__0_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__0_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__0_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__0_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__0_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__0_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__0_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__0_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__0_ccff_tail ) ) ;
cbx_1__1_ cbx_2__1_ (
    .prog_clk ( { ctsbuf_net_1015 } ) ,
    .chanx_left_in ( sb_1__1__0_chanx_right_out ) , 
    .chanx_right_in ( sb_2__1__0_chanx_left_out ) , 
    .ccff_head ( sb_2__1__0_ccff_tail ) , 
    .chanx_left_out ( cbx_1__1__1_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__1__1_chanx_right_out ) , 
    .top_grid_pin_16_ ( cbx_1__1__1_top_grid_pin_16_ ) , 
    .top_grid_pin_17_ ( cbx_1__1__1_top_grid_pin_17_ ) , 
    .top_grid_pin_18_ ( cbx_1__1__1_top_grid_pin_18_ ) , 
    .top_grid_pin_19_ ( cbx_1__1__1_top_grid_pin_19_ ) , 
    .top_grid_pin_20_ ( cbx_1__1__1_top_grid_pin_20_ ) , 
    .top_grid_pin_21_ ( cbx_1__1__1_top_grid_pin_21_ ) , 
    .top_grid_pin_22_ ( cbx_1__1__1_top_grid_pin_22_ ) , 
    .top_grid_pin_23_ ( cbx_1__1__1_top_grid_pin_23_ ) , 
    .top_grid_pin_24_ ( cbx_1__1__1_top_grid_pin_24_ ) , 
    .top_grid_pin_25_ ( cbx_1__1__1_top_grid_pin_25_ ) , 
    .top_grid_pin_26_ ( cbx_1__1__1_top_grid_pin_26_ ) , 
    .top_grid_pin_27_ ( cbx_1__1__1_top_grid_pin_27_ ) , 
    .top_grid_pin_28_ ( cbx_1__1__1_top_grid_pin_28_ ) , 
    .top_grid_pin_29_ ( cbx_1__1__1_top_grid_pin_29_ ) , 
    .top_grid_pin_30_ ( cbx_1__1__1_top_grid_pin_30_ ) , 
    .top_grid_pin_31_ ( cbx_1__1__1_top_grid_pin_31_ ) , 
    .ccff_tail ( cbx_1__1__1_ccff_tail ) ) ;
cbx_1__2_ cbx_1__2_ (
    .prog_clk ( { ctsbuf_net_914 } ) ,
    .chanx_left_in ( sb_0__2__0_chanx_right_out ) , 
    .chanx_right_in ( sb_1__2__0_chanx_left_out ) , 
    .ccff_head ( sb_1__2__0_ccff_tail ) , 
    .chanx_left_out ( cbx_1__2__0_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__2__0_chanx_right_out ) , 
    .top_grid_pin_0_ ( cbx_1__2__0_top_grid_pin_0_ ) , 
    .ccff_tail ( cbx_1__2__0_ccff_tail ) ) ;
cbx_1__2_ cbx_2__2_ (
    .prog_clk ( { ctsbuf_net_16 } ) ,
    .chanx_left_in ( sb_1__2__0_chanx_right_out ) , 
    .chanx_right_in ( sb_2__2__0_chanx_left_out ) , 
    .ccff_head ( sb_2__2__0_ccff_tail ) , 
    .chanx_left_out ( cbx_1__2__1_chanx_left_out ) , 
    .chanx_right_out ( cbx_1__2__1_chanx_right_out ) , 
    .top_grid_pin_0_ ( cbx_1__2__1_top_grid_pin_0_ ) , 
    .ccff_tail ( cbx_1__2__1_ccff_tail ) ) ;
cby_0__1_ cby_0__1_ (
    .prog_clk ( { ctsbuf_net_1520 } ) ,
    .chany_bottom_in ( sb_0__0__0_chany_top_out ) , 
    .chany_top_in ( sb_0__1__0_chany_bottom_out ) , 
    .ccff_head ( sb_0__1__0_ccff_tail ) , 
    .chany_bottom_out ( cby_0__1__0_chany_bottom_out ) , 
    .chany_top_out ( cby_0__1__0_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_0__1__0_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_0__1__0_left_grid_pin_0_ ) , 
    .ccff_tail ( cby_0__1__0_ccff_tail ) ) ;
cby_0__1_ cby_0__2_ (
    .prog_clk ( { ctsbuf_net_1419 } ) ,
    .chany_bottom_in ( sb_0__1__0_chany_top_out ) , 
    .chany_top_in ( sb_0__2__0_chany_bottom_out ) , 
    .ccff_head ( sb_0__2__0_ccff_tail ) , 
    .chany_bottom_out ( cby_0__1__1_chany_bottom_out ) , 
    .chany_top_out ( cby_0__1__1_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_0__1__1_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_0__1__1_left_grid_pin_0_ ) , 
    .ccff_tail ( cby_0__1__1_ccff_tail ) ) ;
cby_1__1_ cby_1__1_ (
    .prog_clk ( { ctsbuf_net_1217 } ) ,
    .chany_bottom_in ( sb_1__0__0_chany_top_out ) , 
    .chany_top_in ( sb_1__1__0_chany_bottom_out ) , 
    .ccff_head ( grid_clb_0_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__0_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__0_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__0_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__0_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__0_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__0_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__0_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__0_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__0_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__0_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__0_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__0_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__0_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__0_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__0_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__0_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__0_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__0_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__0_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__0_ccff_tail ) ) ;
cby_1__1_ cby_1__2_ (
    .prog_clk ( { ctsbuf_net_712 } ) ,
    .chany_bottom_in ( sb_1__1__0_chany_top_out ) , 
    .chany_top_in ( sb_1__2__0_chany_bottom_out ) , 
    .ccff_head ( grid_clb_1_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__1_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__1_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__1_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__1_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__1_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__1_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__1_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__1_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__1_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__1_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__1_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__1_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__1_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__1_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__1_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__1_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__1_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__1_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__1_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__1_ccff_tail ) ) ;
cby_1__1_ cby_2__1_ (
    .prog_clk ( { ctsbuf_net_49 } ) ,
    .chany_bottom_in ( sb_2__0__0_chany_top_out ) , 
    .chany_top_in ( sb_2__1__0_chany_bottom_out ) , 
    .ccff_head ( grid_clb_2_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__2_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__2_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__2_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__2_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__2_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__2_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__2_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__2_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__2_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__2_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__2_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__2_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__2_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__2_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__2_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__2_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__2_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__2_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__2_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__2_ccff_tail ) ) ;
cby_1__1_ cby_2__2_ (
    .prog_clk ( { ctsbuf_net_16 } ) ,
    .chany_bottom_in ( sb_2__1__0_chany_top_out ) , 
    .chany_top_in ( sb_2__2__0_chany_bottom_out ) , 
    .ccff_head ( grid_clb_3_ccff_tail ) , 
    .chany_bottom_out ( cby_1__1__3_chany_bottom_out ) , 
    .chany_top_out ( cby_1__1__3_chany_top_out ) , 
    .right_grid_pin_52_ ( cby_1__1__3_right_grid_pin_52_ ) , 
    .left_grid_pin_0_ ( cby_1__1__3_left_grid_pin_0_ ) , 
    .left_grid_pin_1_ ( cby_1__1__3_left_grid_pin_1_ ) , 
    .left_grid_pin_2_ ( cby_1__1__3_left_grid_pin_2_ ) , 
    .left_grid_pin_3_ ( cby_1__1__3_left_grid_pin_3_ ) , 
    .left_grid_pin_4_ ( cby_1__1__3_left_grid_pin_4_ ) , 
    .left_grid_pin_5_ ( cby_1__1__3_left_grid_pin_5_ ) , 
    .left_grid_pin_6_ ( cby_1__1__3_left_grid_pin_6_ ) , 
    .left_grid_pin_7_ ( cby_1__1__3_left_grid_pin_7_ ) , 
    .left_grid_pin_8_ ( cby_1__1__3_left_grid_pin_8_ ) , 
    .left_grid_pin_9_ ( cby_1__1__3_left_grid_pin_9_ ) , 
    .left_grid_pin_10_ ( cby_1__1__3_left_grid_pin_10_ ) , 
    .left_grid_pin_11_ ( cby_1__1__3_left_grid_pin_11_ ) , 
    .left_grid_pin_12_ ( cby_1__1__3_left_grid_pin_12_ ) , 
    .left_grid_pin_13_ ( cby_1__1__3_left_grid_pin_13_ ) , 
    .left_grid_pin_14_ ( cby_1__1__3_left_grid_pin_14_ ) , 
    .left_grid_pin_15_ ( cby_1__1__3_left_grid_pin_15_ ) , 
    .ccff_tail ( cby_1__1__3_ccff_tail ) ) ;
direct_interc_0 direct_interc_0_ ( 
    .in ( grid_clb_1_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_0_out ) ) ;
direct_interc_1 direct_interc_1_ ( 
    .in ( grid_clb_3_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_1_out ) ) ;
direct_interc_2 direct_interc_2_ ( 
    .in ( grid_clb_0_bottom_width_0_height_0__pin_50_ ) , 
    .out ( direct_interc_2_out ) ) ;
direct_interc_3 direct_interc_3_ ( 
    .in ( grid_clb_1_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_3_out ) ) ;
direct_interc_4 direct_interc_4_ ( 
    .in ( grid_clb_3_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_4_out ) ) ;
direct_interc_5 direct_interc_5_ ( 
    .in ( grid_clb_0_bottom_width_0_height_0__pin_51_ ) , 
    .out ( direct_interc_5_out ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 ropt_h_inst_7301 ( 
    .A ( grid_io_left_1_ccff_tail[0] ) , .X ( ropt_net_25 ) ) ;
sky130_fd_sc_hd__clkinvlp_2 cts_inv_69097180 ( .A ( ctsbuf_net_1924 ) , 
    .Y ( ctsbuf_net_16 ) ) ;
sky130_fd_sc_hd__clkinvlp_2 cts_inv_69107181 ( .A ( ctsbuf_net_1924 ) , 
    .Y ( ctsbuf_net_27 ) ) ;
sky130_fd_sc_hd__clkinvlp_2 cts_inv_69117182 ( .A ( ctsbuf_net_1823 ) , 
    .Y ( ctsbuf_net_38 ) ) ;
sky130_fd_sc_hd__clkinvlp_2 cts_inv_69127183 ( .A ( ctsbuf_net_1924 ) , 
    .Y ( ctsbuf_net_49 ) ) ;
sky130_fd_sc_hd__clkinvlp_2 cts_inv_69137184 ( .A ( ctsbuf_net_1924 ) , 
    .Y ( ctsbuf_net_510 ) ) ;
sky130_fd_sc_hd__clkinvlp_2 cts_inv_69147185 ( .A ( ctsbuf_net_1823 ) , 
    .Y ( ctsbuf_net_611 ) ) ;
sky130_fd_sc_hd__clkinvlp_2 cts_inv_69157186 ( .A ( ctsbuf_net_1823 ) , 
    .Y ( ctsbuf_net_712 ) ) ;
sky130_fd_sc_hd__clkinvlp_2 cts_inv_69167187 ( .A ( ctsbuf_net_1924 ) , 
    .Y ( ctsbuf_net_813 ) ) ;
sky130_fd_sc_hd__clkinvlp_2 cts_inv_69177188 ( .A ( ctsbuf_net_1823 ) , 
    .Y ( ctsbuf_net_914 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 ropt_h_inst_7302 ( .A ( ropt_net_25 ) , 
    .X ( ropt_net_26 ) ) ;
sky130_fd_sc_hd__clkinvlp_2 cts_inv_69197190 ( .A ( ctsbuf_net_1924 ) , 
    .Y ( ctsbuf_net_1116 ) ) ;
sky130_fd_sc_hd__clkinvlp_2 cts_inv_69207191 ( .A ( ctsbuf_net_1924 ) , 
    .Y ( ctsbuf_net_1217 ) ) ;
sky130_fd_sc_hd__clkinvlp_2 cts_inv_69217192 ( .A ( ctsbuf_net_1823 ) , 
    .Y ( ctsbuf_net_1318 ) ) ;
sky130_fd_sc_hd__clkinvlp_2 cts_inv_69227193 ( .A ( ctsbuf_net_1823 ) , 
    .Y ( ctsbuf_net_1419 ) ) ;
sky130_fd_sc_hd__clkinvlp_2 cts_inv_69237194 ( .A ( ctsbuf_net_1823 ) , 
    .Y ( ctsbuf_net_1520 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 ropt_h_inst_7303 ( .A ( ropt_net_26 ) , 
    .X ( ropt_net_27 ) ) ;
sky130_fd_sc_hd__clkinvlp_2 cts_inv_69257196 ( .A ( ctsbuf_net_1924 ) , 
    .Y ( ctsbuf_net_1722 ) ) ;
sky130_fd_sc_hd__bufinv_8 cts_inv_69247195_69267197 ( 
    .A ( SYNOPSYS_UNCONNECTED_1 ) , .Y ( SYNOPSYS_UNCONNECTED_2 ) ) ;
sky130_fd_sc_hd__clkinv_16 cts_inv_69187189_69277198 ( 
    .A ( SYNOPSYS_UNCONNECTED_3 ) , .Y ( p_abuf0 ) ) ;
sky130_fd_sc_hd__clkinvlp_2 cts_inv_69397210 ( .A ( prog_clk[0] ) , 
    .Y ( ctsbuf_net_1823 ) ) ;
sky130_fd_sc_hd__clkinvlp_2 cts_inv_69407211 ( .A ( prog_clk[0] ) , 
    .Y ( ctsbuf_net_1924 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 ropt_h_inst_7304 ( 
    .A ( grid_io_top_1_ccff_tail[0] ) , .X ( ropt_net_28 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 ropt_h_inst_7305 ( .A ( ropt_net_28 ) , 
    .X ( ropt_net_29 ) ) ;
sky130_fd_sc_hd__dlygate4sd3_1 ropt_h_inst_7306 ( 
    .A ( grid_io_left_0_ccff_tail[0] ) , .X ( ropt_net_30 ) ) ;
sky130_fd_sc_hd__dlygate4sd2_1 ropt_h_inst_7307 ( .A ( ropt_net_30 ) , 
    .X ( ropt_net_31 ) ) ;
endmodule


