//Generated from netlist by SpyDrNet
//netlist name: FPGA88_SOFA_A
module EMBEDDED_IO_HD
(
    FPGA_DIR,
    FPGA_OUT,
    IO_ISOL_N,
    SOC_IN,
    FPGA_IN,
    SOC_DIR,
    SOC_OUT
);

    input FPGA_DIR;
    input FPGA_OUT;
    input IO_ISOL_N;
    input SOC_IN;
    output FPGA_IN;
    output SOC_DIR;
    output SOC_OUT;

    wire FPGA_DIR;
    wire FPGA_IN;
    wire FPGA_OUT;
    wire IO_ISOL_N;
    wire SOC_DIR;
    wire SOC_IN;
    wire SOC_OUT;

endmodule

